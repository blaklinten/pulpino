module matrix_multiply #(
  parameter mat_size = 2,
  parameter dat_size = 8
) (
//  input  logic            start        ,
//  output logic            done         ,
  input  logic            clk          , 
  input  logic [1023:0][7:0] mat_A ,
  input  logic [1023:0][7:0] mat_B ,
  output logic [1023:0][15:0] mat_C
);

  always @(posedge clk)
  begin
    mat_C[0] <= 
               mat_A[0];// * mat_B[0] +
//             mat_A[1] * mat_B[32] +
//             mat_A[2] * mat_B[64] +
//             mat_A[3] * mat_B[96] +
//             mat_A[4] * mat_B[128] +
//             mat_A[5] * mat_B[160] +
//             mat_A[6] * mat_B[192] +
//             mat_A[7] * mat_B[224] +
//             mat_A[8] * mat_B[256] +
//             mat_A[9] * mat_B[288] +
//             mat_A[10] * mat_B[320] +
//             mat_A[11] * mat_B[352] +
//             mat_A[12] * mat_B[384] +
//             mat_A[13] * mat_B[416] +
//             mat_A[14] * mat_B[448] +
//             mat_A[15] * mat_B[480] +
//             mat_A[16] * mat_B[512] +
//             mat_A[17] * mat_B[544] +
//             mat_A[18] * mat_B[576] +
//             mat_A[19] * mat_B[608] +
//             mat_A[20] * mat_B[640] +
//             mat_A[21] * mat_B[672] +
//             mat_A[22] * mat_B[704] +
//             mat_A[23] * mat_B[736] +
//             mat_A[24] * mat_B[768] +
//             mat_A[25] * mat_B[800] +
//             mat_A[26] * mat_B[832] +
//             mat_A[27] * mat_B[864] +
//             mat_A[28] * mat_B[896] +
//             mat_A[29] * mat_B[928] +
//             mat_A[30] * mat_B[960] +
//             mat_A[31] * mat_B[992];
    mat_C[1] <= 
//             mat_A[0] * mat_B[1] +
               mat_A[1];// * mat_B[33] +
//             mat_A[2] * mat_B[65] +
//             mat_A[3] * mat_B[97] +
//             mat_A[4] * mat_B[129] +
//             mat_A[5] * mat_B[161] +
//             mat_A[6] * mat_B[193] +
//             mat_A[7] * mat_B[225] +
//             mat_A[8] * mat_B[257] +
//             mat_A[9] * mat_B[289] +
//             mat_A[10] * mat_B[321] +
//             mat_A[11] * mat_B[353] +
//             mat_A[12] * mat_B[385] +
//             mat_A[13] * mat_B[417] +
//             mat_A[14] * mat_B[449] +
//             mat_A[15] * mat_B[481] +
//             mat_A[16] * mat_B[513] +
//             mat_A[17] * mat_B[545] +
//             mat_A[18] * mat_B[577] +
//             mat_A[19] * mat_B[609] +
//             mat_A[20] * mat_B[641] +
//             mat_A[21] * mat_B[673] +
//             mat_A[22] * mat_B[705] +
//             mat_A[23] * mat_B[737] +
//             mat_A[24] * mat_B[769] +
//             mat_A[25] * mat_B[801] +
//             mat_A[26] * mat_B[833] +
//             mat_A[27] * mat_B[865] +
//             mat_A[28] * mat_B[897] +
//             mat_A[29] * mat_B[929] +
//             mat_A[30] * mat_B[961] +
//             mat_A[31] * mat_B[993];
    mat_C[2] <= 
//             mat_A[0] * mat_B[2] +
//             mat_A[1] * mat_B[34] +
               mat_A[2];// * mat_B[66] +
//             mat_A[3] * mat_B[98] +
//             mat_A[4] * mat_B[130] +
//             mat_A[5] * mat_B[162] +
//             mat_A[6] * mat_B[194] +
//             mat_A[7] * mat_B[226] +
//             mat_A[8] * mat_B[258] +
//             mat_A[9] * mat_B[290] +
//             mat_A[10] * mat_B[322] +
//             mat_A[11] * mat_B[354] +
//             mat_A[12] * mat_B[386] +
//             mat_A[13] * mat_B[418] +
//             mat_A[14] * mat_B[450] +
//             mat_A[15] * mat_B[482] +
//             mat_A[16] * mat_B[514] +
//             mat_A[17] * mat_B[546] +
//             mat_A[18] * mat_B[578] +
//             mat_A[19] * mat_B[610] +
//             mat_A[20] * mat_B[642] +
//             mat_A[21] * mat_B[674] +
//             mat_A[22] * mat_B[706] +
//             mat_A[23] * mat_B[738] +
//             mat_A[24] * mat_B[770] +
//             mat_A[25] * mat_B[802] +
//             mat_A[26] * mat_B[834] +
//             mat_A[27] * mat_B[866] +
//             mat_A[28] * mat_B[898] +
//             mat_A[29] * mat_B[930] +
//             mat_A[30] * mat_B[962] +
//             mat_A[31] * mat_B[994];
    mat_C[3] <= 
//             mat_A[0] * mat_B[3] +
//             mat_A[1] * mat_B[35] +
//             mat_A[2] * mat_B[67] +
               mat_A[3];// * mat_B[99] +
//             mat_A[4] * mat_B[131] +
//             mat_A[5] * mat_B[163] +
//             mat_A[6] * mat_B[195] +
//             mat_A[7] * mat_B[227] +
//             mat_A[8] * mat_B[259] +
//             mat_A[9] * mat_B[291] +
//             mat_A[10] * mat_B[323] +
//             mat_A[11] * mat_B[355] +
//             mat_A[12] * mat_B[387] +
//             mat_A[13] * mat_B[419] +
//             mat_A[14] * mat_B[451] +
//             mat_A[15] * mat_B[483] +
//             mat_A[16] * mat_B[515] +
//             mat_A[17] * mat_B[547] +
//             mat_A[18] * mat_B[579] +
//             mat_A[19] * mat_B[611] +
//             mat_A[20] * mat_B[643] +
//             mat_A[21] * mat_B[675] +
//             mat_A[22] * mat_B[707] +
//             mat_A[23] * mat_B[739] +
//             mat_A[24] * mat_B[771] +
//             mat_A[25] * mat_B[803] +
//             mat_A[26] * mat_B[835] +
//             mat_A[27] * mat_B[867] +
//             mat_A[28] * mat_B[899] +
//             mat_A[29] * mat_B[931] +
//             mat_A[30] * mat_B[963] +
//             mat_A[31] * mat_B[995];
    mat_C[4] <= 
//             mat_A[0] * mat_B[4] +
//             mat_A[1] * mat_B[36] +
//             mat_A[2] * mat_B[68] +
//             mat_A[3] * mat_B[100] +
               mat_A[4];// * mat_B[132] +
//             mat_A[5] * mat_B[164] +
//             mat_A[6] * mat_B[196] +
//             mat_A[7] * mat_B[228] +
//             mat_A[8] * mat_B[260] +
//             mat_A[9] * mat_B[292] +
//             mat_A[10] * mat_B[324] +
//             mat_A[11] * mat_B[356] +
//             mat_A[12] * mat_B[388] +
//             mat_A[13] * mat_B[420] +
//             mat_A[14] * mat_B[452] +
//             mat_A[15] * mat_B[484] +
//             mat_A[16] * mat_B[516] +
//             mat_A[17] * mat_B[548] +
//             mat_A[18] * mat_B[580] +
//             mat_A[19] * mat_B[612] +
//             mat_A[20] * mat_B[644] +
//             mat_A[21] * mat_B[676] +
//             mat_A[22] * mat_B[708] +
//             mat_A[23] * mat_B[740] +
//             mat_A[24] * mat_B[772] +
//             mat_A[25] * mat_B[804] +
//             mat_A[26] * mat_B[836] +
//             mat_A[27] * mat_B[868] +
//             mat_A[28] * mat_B[900] +
//             mat_A[29] * mat_B[932] +
//             mat_A[30] * mat_B[964] +
//             mat_A[31] * mat_B[996];
    mat_C[5] <= 
//             mat_A[0] * mat_B[5] +
//             mat_A[1] * mat_B[37] +
//             mat_A[2] * mat_B[69] +
//             mat_A[3] * mat_B[101] +
//             mat_A[4] * mat_B[133] +
               mat_A[5];// * mat_B[165] +
//             mat_A[6] * mat_B[197] +
//             mat_A[7] * mat_B[229] +
//             mat_A[8] * mat_B[261] +
//             mat_A[9] * mat_B[293] +
//             mat_A[10] * mat_B[325] +
//             mat_A[11] * mat_B[357] +
//             mat_A[12] * mat_B[389] +
//             mat_A[13] * mat_B[421] +
//             mat_A[14] * mat_B[453] +
//             mat_A[15] * mat_B[485] +
//             mat_A[16] * mat_B[517] +
//             mat_A[17] * mat_B[549] +
//             mat_A[18] * mat_B[581] +
//             mat_A[19] * mat_B[613] +
//             mat_A[20] * mat_B[645] +
//             mat_A[21] * mat_B[677] +
//             mat_A[22] * mat_B[709] +
//             mat_A[23] * mat_B[741] +
//             mat_A[24] * mat_B[773] +
//             mat_A[25] * mat_B[805] +
//             mat_A[26] * mat_B[837] +
//             mat_A[27] * mat_B[869] +
//             mat_A[28] * mat_B[901] +
//             mat_A[29] * mat_B[933] +
//             mat_A[30] * mat_B[965] +
//             mat_A[31] * mat_B[997];
    mat_C[6] <= 
//             mat_A[0] * mat_B[6] +
//             mat_A[1] * mat_B[38] +
//             mat_A[2] * mat_B[70] +
//             mat_A[3] * mat_B[102] +
//             mat_A[4] * mat_B[134] +
//             mat_A[5] * mat_B[166] +
               mat_A[6];// * mat_B[198] +
//             mat_A[7] * mat_B[230] +
//             mat_A[8] * mat_B[262] +
//             mat_A[9] * mat_B[294] +
//             mat_A[10] * mat_B[326] +
//             mat_A[11] * mat_B[358] +
//             mat_A[12] * mat_B[390] +
//             mat_A[13] * mat_B[422] +
//             mat_A[14] * mat_B[454] +
//             mat_A[15] * mat_B[486] +
//             mat_A[16] * mat_B[518] +
//             mat_A[17] * mat_B[550] +
//             mat_A[18] * mat_B[582] +
//             mat_A[19] * mat_B[614] +
//             mat_A[20] * mat_B[646] +
//             mat_A[21] * mat_B[678] +
//             mat_A[22] * mat_B[710] +
//             mat_A[23] * mat_B[742] +
//             mat_A[24] * mat_B[774] +
//             mat_A[25] * mat_B[806] +
//             mat_A[26] * mat_B[838] +
//             mat_A[27] * mat_B[870] +
//             mat_A[28] * mat_B[902] +
//             mat_A[29] * mat_B[934] +
//             mat_A[30] * mat_B[966] +
//             mat_A[31] * mat_B[998];
    mat_C[7] <= 
//             mat_A[0] * mat_B[7] +
//             mat_A[1] * mat_B[39] +
//             mat_A[2] * mat_B[71] +
//             mat_A[3] * mat_B[103] +
//             mat_A[4] * mat_B[135] +
//             mat_A[5] * mat_B[167] +
//             mat_A[6] * mat_B[199] +
               mat_A[7];// * mat_B[231] +
//             mat_A[8] * mat_B[263] +
//             mat_A[9] * mat_B[295] +
//             mat_A[10] * mat_B[327] +
//             mat_A[11] * mat_B[359] +
//             mat_A[12] * mat_B[391] +
//             mat_A[13] * mat_B[423] +
//             mat_A[14] * mat_B[455] +
//             mat_A[15] * mat_B[487] +
//             mat_A[16] * mat_B[519] +
//             mat_A[17] * mat_B[551] +
//             mat_A[18] * mat_B[583] +
//             mat_A[19] * mat_B[615] +
//             mat_A[20] * mat_B[647] +
//             mat_A[21] * mat_B[679] +
//             mat_A[22] * mat_B[711] +
//             mat_A[23] * mat_B[743] +
//             mat_A[24] * mat_B[775] +
//             mat_A[25] * mat_B[807] +
//             mat_A[26] * mat_B[839] +
//             mat_A[27] * mat_B[871] +
//             mat_A[28] * mat_B[903] +
//             mat_A[29] * mat_B[935] +
//             mat_A[30] * mat_B[967] +
//             mat_A[31] * mat_B[999];
//  mat_C[8] <= 
//             mat_A[0] * mat_B[8] +
//             mat_A[1] * mat_B[40] +
//             mat_A[2] * mat_B[72] +
//             mat_A[3] * mat_B[104] +
//             mat_A[4] * mat_B[136] +
//             mat_A[5] * mat_B[168] +
//             mat_A[6] * mat_B[200] +
//             mat_A[7] * mat_B[232] +
//             mat_A[8] * mat_B[264] +
//             mat_A[9] * mat_B[296] +
//             mat_A[10] * mat_B[328] +
//             mat_A[11] * mat_B[360] +
//             mat_A[12] * mat_B[392] +
//             mat_A[13] * mat_B[424] +
//             mat_A[14] * mat_B[456] +
//             mat_A[15] * mat_B[488] +
//             mat_A[16] * mat_B[520] +
//             mat_A[17] * mat_B[552] +
//             mat_A[18] * mat_B[584] +
//             mat_A[19] * mat_B[616] +
//             mat_A[20] * mat_B[648] +
//             mat_A[21] * mat_B[680] +
//             mat_A[22] * mat_B[712] +
//             mat_A[23] * mat_B[744] +
//             mat_A[24] * mat_B[776] +
//             mat_A[25] * mat_B[808] +
//             mat_A[26] * mat_B[840] +
//             mat_A[27] * mat_B[872] +
//             mat_A[28] * mat_B[904] +
//             mat_A[29] * mat_B[936] +
//             mat_A[30] * mat_B[968] +
//             mat_A[31] * mat_B[1000];
//  mat_C[9] <= 
//             mat_A[0] * mat_B[9] +
//             mat_A[1] * mat_B[41] +
//             mat_A[2] * mat_B[73] +
//             mat_A[3] * mat_B[105] +
//             mat_A[4] * mat_B[137] +
//             mat_A[5] * mat_B[169] +
//             mat_A[6] * mat_B[201] +
//             mat_A[7] * mat_B[233] +
//             mat_A[8] * mat_B[265] +
//             mat_A[9] * mat_B[297] +
//             mat_A[10] * mat_B[329] +
//             mat_A[11] * mat_B[361] +
//             mat_A[12] * mat_B[393] +
//             mat_A[13] * mat_B[425] +
//             mat_A[14] * mat_B[457] +
//             mat_A[15] * mat_B[489] +
//             mat_A[16] * mat_B[521] +
//             mat_A[17] * mat_B[553] +
//             mat_A[18] * mat_B[585] +
//             mat_A[19] * mat_B[617] +
//             mat_A[20] * mat_B[649] +
//             mat_A[21] * mat_B[681] +
//             mat_A[22] * mat_B[713] +
//             mat_A[23] * mat_B[745] +
//             mat_A[24] * mat_B[777] +
//             mat_A[25] * mat_B[809] +
//             mat_A[26] * mat_B[841] +
//             mat_A[27] * mat_B[873] +
//             mat_A[28] * mat_B[905] +
//             mat_A[29] * mat_B[937] +
//             mat_A[30] * mat_B[969] +
//             mat_A[31] * mat_B[1001];
//  mat_C[10] <= 
//             mat_A[0] * mat_B[10] +
//             mat_A[1] * mat_B[42] +
//             mat_A[2] * mat_B[74] +
//             mat_A[3] * mat_B[106] +
//             mat_A[4] * mat_B[138] +
//             mat_A[5] * mat_B[170] +
//             mat_A[6] * mat_B[202] +
//             mat_A[7] * mat_B[234] +
//             mat_A[8] * mat_B[266] +
//             mat_A[9] * mat_B[298] +
//             mat_A[10] * mat_B[330] +
//             mat_A[11] * mat_B[362] +
//             mat_A[12] * mat_B[394] +
//             mat_A[13] * mat_B[426] +
//             mat_A[14] * mat_B[458] +
//             mat_A[15] * mat_B[490] +
//             mat_A[16] * mat_B[522] +
//             mat_A[17] * mat_B[554] +
//             mat_A[18] * mat_B[586] +
//             mat_A[19] * mat_B[618] +
//             mat_A[20] * mat_B[650] +
//             mat_A[21] * mat_B[682] +
//             mat_A[22] * mat_B[714] +
//             mat_A[23] * mat_B[746] +
//             mat_A[24] * mat_B[778] +
//             mat_A[25] * mat_B[810] +
//             mat_A[26] * mat_B[842] +
//             mat_A[27] * mat_B[874] +
//             mat_A[28] * mat_B[906] +
//             mat_A[29] * mat_B[938] +
//             mat_A[30] * mat_B[970] +
//             mat_A[31] * mat_B[1002];
//  mat_C[11] <= 
//             mat_A[0] * mat_B[11] +
//             mat_A[1] * mat_B[43] +
//             mat_A[2] * mat_B[75] +
//             mat_A[3] * mat_B[107] +
//             mat_A[4] * mat_B[139] +
//             mat_A[5] * mat_B[171] +
//             mat_A[6] * mat_B[203] +
//             mat_A[7] * mat_B[235] +
//             mat_A[8] * mat_B[267] +
//             mat_A[9] * mat_B[299] +
//             mat_A[10] * mat_B[331] +
//             mat_A[11] * mat_B[363] +
//             mat_A[12] * mat_B[395] +
//             mat_A[13] * mat_B[427] +
//             mat_A[14] * mat_B[459] +
//             mat_A[15] * mat_B[491] +
//             mat_A[16] * mat_B[523] +
//             mat_A[17] * mat_B[555] +
//             mat_A[18] * mat_B[587] +
//             mat_A[19] * mat_B[619] +
//             mat_A[20] * mat_B[651] +
//             mat_A[21] * mat_B[683] +
//             mat_A[22] * mat_B[715] +
//             mat_A[23] * mat_B[747] +
//             mat_A[24] * mat_B[779] +
//             mat_A[25] * mat_B[811] +
//             mat_A[26] * mat_B[843] +
//             mat_A[27] * mat_B[875] +
//             mat_A[28] * mat_B[907] +
//             mat_A[29] * mat_B[939] +
//             mat_A[30] * mat_B[971] +
//             mat_A[31] * mat_B[1003];
//  mat_C[12] <= 
//             mat_A[0] * mat_B[12] +
//             mat_A[1] * mat_B[44] +
//             mat_A[2] * mat_B[76] +
//             mat_A[3] * mat_B[108] +
//             mat_A[4] * mat_B[140] +
//             mat_A[5] * mat_B[172] +
//             mat_A[6] * mat_B[204] +
//             mat_A[7] * mat_B[236] +
//             mat_A[8] * mat_B[268] +
//             mat_A[9] * mat_B[300] +
//             mat_A[10] * mat_B[332] +
//             mat_A[11] * mat_B[364] +
//             mat_A[12] * mat_B[396] +
//             mat_A[13] * mat_B[428] +
//             mat_A[14] * mat_B[460] +
//             mat_A[15] * mat_B[492] +
//             mat_A[16] * mat_B[524] +
//             mat_A[17] * mat_B[556] +
//             mat_A[18] * mat_B[588] +
//             mat_A[19] * mat_B[620] +
//             mat_A[20] * mat_B[652] +
//             mat_A[21] * mat_B[684] +
//             mat_A[22] * mat_B[716] +
//             mat_A[23] * mat_B[748] +
//             mat_A[24] * mat_B[780] +
//             mat_A[25] * mat_B[812] +
//             mat_A[26] * mat_B[844] +
//             mat_A[27] * mat_B[876] +
//             mat_A[28] * mat_B[908] +
//             mat_A[29] * mat_B[940] +
//             mat_A[30] * mat_B[972] +
//             mat_A[31] * mat_B[1004];
//  mat_C[13] <= 
//             mat_A[0] * mat_B[13] +
//             mat_A[1] * mat_B[45] +
//             mat_A[2] * mat_B[77] +
//             mat_A[3] * mat_B[109] +
//             mat_A[4] * mat_B[141] +
//             mat_A[5] * mat_B[173] +
//             mat_A[6] * mat_B[205] +
//             mat_A[7] * mat_B[237] +
//             mat_A[8] * mat_B[269] +
//             mat_A[9] * mat_B[301] +
//             mat_A[10] * mat_B[333] +
//             mat_A[11] * mat_B[365] +
//             mat_A[12] * mat_B[397] +
//             mat_A[13] * mat_B[429] +
//             mat_A[14] * mat_B[461] +
//             mat_A[15] * mat_B[493] +
//             mat_A[16] * mat_B[525] +
//             mat_A[17] * mat_B[557] +
//             mat_A[18] * mat_B[589] +
//             mat_A[19] * mat_B[621] +
//             mat_A[20] * mat_B[653] +
//             mat_A[21] * mat_B[685] +
//             mat_A[22] * mat_B[717] +
//             mat_A[23] * mat_B[749] +
//             mat_A[24] * mat_B[781] +
//             mat_A[25] * mat_B[813] +
//             mat_A[26] * mat_B[845] +
//             mat_A[27] * mat_B[877] +
//             mat_A[28] * mat_B[909] +
//             mat_A[29] * mat_B[941] +
//             mat_A[30] * mat_B[973] +
//             mat_A[31] * mat_B[1005];
//  mat_C[14] <= 
//             mat_A[0] * mat_B[14] +
//             mat_A[1] * mat_B[46] +
//             mat_A[2] * mat_B[78] +
//             mat_A[3] * mat_B[110] +
//             mat_A[4] * mat_B[142] +
//             mat_A[5] * mat_B[174] +
//             mat_A[6] * mat_B[206] +
//             mat_A[7] * mat_B[238] +
//             mat_A[8] * mat_B[270] +
//             mat_A[9] * mat_B[302] +
//             mat_A[10] * mat_B[334] +
//             mat_A[11] * mat_B[366] +
//             mat_A[12] * mat_B[398] +
//             mat_A[13] * mat_B[430] +
//             mat_A[14] * mat_B[462] +
//             mat_A[15] * mat_B[494] +
//             mat_A[16] * mat_B[526] +
//             mat_A[17] * mat_B[558] +
//             mat_A[18] * mat_B[590] +
//             mat_A[19] * mat_B[622] +
//             mat_A[20] * mat_B[654] +
//             mat_A[21] * mat_B[686] +
//             mat_A[22] * mat_B[718] +
//             mat_A[23] * mat_B[750] +
//             mat_A[24] * mat_B[782] +
//             mat_A[25] * mat_B[814] +
//             mat_A[26] * mat_B[846] +
//             mat_A[27] * mat_B[878] +
//             mat_A[28] * mat_B[910] +
//             mat_A[29] * mat_B[942] +
//             mat_A[30] * mat_B[974] +
//             mat_A[31] * mat_B[1006];
//  mat_C[15] <= 
//             mat_A[0] * mat_B[15] +
//             mat_A[1] * mat_B[47] +
//             mat_A[2] * mat_B[79] +
//             mat_A[3] * mat_B[111] +
//             mat_A[4] * mat_B[143] +
//             mat_A[5] * mat_B[175] +
//             mat_A[6] * mat_B[207] +
//             mat_A[7] * mat_B[239] +
//             mat_A[8] * mat_B[271] +
//             mat_A[9] * mat_B[303] +
//             mat_A[10] * mat_B[335] +
//             mat_A[11] * mat_B[367] +
//             mat_A[12] * mat_B[399] +
//             mat_A[13] * mat_B[431] +
//             mat_A[14] * mat_B[463] +
//             mat_A[15] * mat_B[495] +
//             mat_A[16] * mat_B[527] +
//             mat_A[17] * mat_B[559] +
//             mat_A[18] * mat_B[591] +
//             mat_A[19] * mat_B[623] +
//             mat_A[20] * mat_B[655] +
//             mat_A[21] * mat_B[687] +
//             mat_A[22] * mat_B[719] +
//             mat_A[23] * mat_B[751] +
//             mat_A[24] * mat_B[783] +
//             mat_A[25] * mat_B[815] +
//             mat_A[26] * mat_B[847] +
//             mat_A[27] * mat_B[879] +
//             mat_A[28] * mat_B[911] +
//             mat_A[29] * mat_B[943] +
//             mat_A[30] * mat_B[975] +
//             mat_A[31] * mat_B[1007];
//  mat_C[16] <= 
//             mat_A[0] * mat_B[16] +
//             mat_A[1] * mat_B[48] +
//             mat_A[2] * mat_B[80] +
//             mat_A[3] * mat_B[112] +
//             mat_A[4] * mat_B[144] +
//             mat_A[5] * mat_B[176] +
//             mat_A[6] * mat_B[208] +
//             mat_A[7] * mat_B[240] +
//             mat_A[8] * mat_B[272] +
//             mat_A[9] * mat_B[304] +
//             mat_A[10] * mat_B[336] +
//             mat_A[11] * mat_B[368] +
//             mat_A[12] * mat_B[400] +
//             mat_A[13] * mat_B[432] +
//             mat_A[14] * mat_B[464] +
//             mat_A[15] * mat_B[496] +
//             mat_A[16] * mat_B[528] +
//             mat_A[17] * mat_B[560] +
//             mat_A[18] * mat_B[592] +
//             mat_A[19] * mat_B[624] +
//             mat_A[20] * mat_B[656] +
//             mat_A[21] * mat_B[688] +
//             mat_A[22] * mat_B[720] +
//             mat_A[23] * mat_B[752] +
//             mat_A[24] * mat_B[784] +
//             mat_A[25] * mat_B[816] +
//             mat_A[26] * mat_B[848] +
//             mat_A[27] * mat_B[880] +
//             mat_A[28] * mat_B[912] +
//             mat_A[29] * mat_B[944] +
//             mat_A[30] * mat_B[976] +
//             mat_A[31] * mat_B[1008];
//  mat_C[17] <= 
//             mat_A[0] * mat_B[17] +
//             mat_A[1] * mat_B[49] +
//             mat_A[2] * mat_B[81] +
//             mat_A[3] * mat_B[113] +
//             mat_A[4] * mat_B[145] +
//             mat_A[5] * mat_B[177] +
//             mat_A[6] * mat_B[209] +
//             mat_A[7] * mat_B[241] +
//             mat_A[8] * mat_B[273] +
//             mat_A[9] * mat_B[305] +
//             mat_A[10] * mat_B[337] +
//             mat_A[11] * mat_B[369] +
//             mat_A[12] * mat_B[401] +
//             mat_A[13] * mat_B[433] +
//             mat_A[14] * mat_B[465] +
//             mat_A[15] * mat_B[497] +
//             mat_A[16] * mat_B[529] +
//             mat_A[17] * mat_B[561] +
//             mat_A[18] * mat_B[593] +
//             mat_A[19] * mat_B[625] +
//             mat_A[20] * mat_B[657] +
//             mat_A[21] * mat_B[689] +
//             mat_A[22] * mat_B[721] +
//             mat_A[23] * mat_B[753] +
//             mat_A[24] * mat_B[785] +
//             mat_A[25] * mat_B[817] +
//             mat_A[26] * mat_B[849] +
//             mat_A[27] * mat_B[881] +
//             mat_A[28] * mat_B[913] +
//             mat_A[29] * mat_B[945] +
//             mat_A[30] * mat_B[977] +
//             mat_A[31] * mat_B[1009];
//  mat_C[18] <= 
//             mat_A[0] * mat_B[18] +
//             mat_A[1] * mat_B[50] +
//             mat_A[2] * mat_B[82] +
//             mat_A[3] * mat_B[114] +
//             mat_A[4] * mat_B[146] +
//             mat_A[5] * mat_B[178] +
//             mat_A[6] * mat_B[210] +
//             mat_A[7] * mat_B[242] +
//             mat_A[8] * mat_B[274] +
//             mat_A[9] * mat_B[306] +
//             mat_A[10] * mat_B[338] +
//             mat_A[11] * mat_B[370] +
//             mat_A[12] * mat_B[402] +
//             mat_A[13] * mat_B[434] +
//             mat_A[14] * mat_B[466] +
//             mat_A[15] * mat_B[498] +
//             mat_A[16] * mat_B[530] +
//             mat_A[17] * mat_B[562] +
//             mat_A[18] * mat_B[594] +
//             mat_A[19] * mat_B[626] +
//             mat_A[20] * mat_B[658] +
//             mat_A[21] * mat_B[690] +
//             mat_A[22] * mat_B[722] +
//             mat_A[23] * mat_B[754] +
//             mat_A[24] * mat_B[786] +
//             mat_A[25] * mat_B[818] +
//             mat_A[26] * mat_B[850] +
//             mat_A[27] * mat_B[882] +
//             mat_A[28] * mat_B[914] +
//             mat_A[29] * mat_B[946] +
//             mat_A[30] * mat_B[978] +
//             mat_A[31] * mat_B[1010];
//  mat_C[19] <= 
//             mat_A[0] * mat_B[19] +
//             mat_A[1] * mat_B[51] +
//             mat_A[2] * mat_B[83] +
//             mat_A[3] * mat_B[115] +
//             mat_A[4] * mat_B[147] +
//             mat_A[5] * mat_B[179] +
//             mat_A[6] * mat_B[211] +
//             mat_A[7] * mat_B[243] +
//             mat_A[8] * mat_B[275] +
//             mat_A[9] * mat_B[307] +
//             mat_A[10] * mat_B[339] +
//             mat_A[11] * mat_B[371] +
//             mat_A[12] * mat_B[403] +
//             mat_A[13] * mat_B[435] +
//             mat_A[14] * mat_B[467] +
//             mat_A[15] * mat_B[499] +
//             mat_A[16] * mat_B[531] +
//             mat_A[17] * mat_B[563] +
//             mat_A[18] * mat_B[595] +
//             mat_A[19] * mat_B[627] +
//             mat_A[20] * mat_B[659] +
//             mat_A[21] * mat_B[691] +
//             mat_A[22] * mat_B[723] +
//             mat_A[23] * mat_B[755] +
//             mat_A[24] * mat_B[787] +
//             mat_A[25] * mat_B[819] +
//             mat_A[26] * mat_B[851] +
//             mat_A[27] * mat_B[883] +
//             mat_A[28] * mat_B[915] +
//             mat_A[29] * mat_B[947] +
//             mat_A[30] * mat_B[979] +
//             mat_A[31] * mat_B[1011];
//  mat_C[20] <= 
//             mat_A[0] * mat_B[20] +
//             mat_A[1] * mat_B[52] +
//             mat_A[2] * mat_B[84] +
//             mat_A[3] * mat_B[116] +
//             mat_A[4] * mat_B[148] +
//             mat_A[5] * mat_B[180] +
//             mat_A[6] * mat_B[212] +
//             mat_A[7] * mat_B[244] +
//             mat_A[8] * mat_B[276] +
//             mat_A[9] * mat_B[308] +
//             mat_A[10] * mat_B[340] +
//             mat_A[11] * mat_B[372] +
//             mat_A[12] * mat_B[404] +
//             mat_A[13] * mat_B[436] +
//             mat_A[14] * mat_B[468] +
//             mat_A[15] * mat_B[500] +
//             mat_A[16] * mat_B[532] +
//             mat_A[17] * mat_B[564] +
//             mat_A[18] * mat_B[596] +
//             mat_A[19] * mat_B[628] +
//             mat_A[20] * mat_B[660] +
//             mat_A[21] * mat_B[692] +
//             mat_A[22] * mat_B[724] +
//             mat_A[23] * mat_B[756] +
//             mat_A[24] * mat_B[788] +
//             mat_A[25] * mat_B[820] +
//             mat_A[26] * mat_B[852] +
//             mat_A[27] * mat_B[884] +
//             mat_A[28] * mat_B[916] +
//             mat_A[29] * mat_B[948] +
//             mat_A[30] * mat_B[980] +
//             mat_A[31] * mat_B[1012];
//  mat_C[21] <= 
//             mat_A[0] * mat_B[21] +
//             mat_A[1] * mat_B[53] +
//             mat_A[2] * mat_B[85] +
//             mat_A[3] * mat_B[117] +
//             mat_A[4] * mat_B[149] +
//             mat_A[5] * mat_B[181] +
//             mat_A[6] * mat_B[213] +
//             mat_A[7] * mat_B[245] +
//             mat_A[8] * mat_B[277] +
//             mat_A[9] * mat_B[309] +
//             mat_A[10] * mat_B[341] +
//             mat_A[11] * mat_B[373] +
//             mat_A[12] * mat_B[405] +
//             mat_A[13] * mat_B[437] +
//             mat_A[14] * mat_B[469] +
//             mat_A[15] * mat_B[501] +
//             mat_A[16] * mat_B[533] +
//             mat_A[17] * mat_B[565] +
//             mat_A[18] * mat_B[597] +
//             mat_A[19] * mat_B[629] +
//             mat_A[20] * mat_B[661] +
//             mat_A[21] * mat_B[693] +
//             mat_A[22] * mat_B[725] +
//             mat_A[23] * mat_B[757] +
//             mat_A[24] * mat_B[789] +
//             mat_A[25] * mat_B[821] +
//             mat_A[26] * mat_B[853] +
//             mat_A[27] * mat_B[885] +
//             mat_A[28] * mat_B[917] +
//             mat_A[29] * mat_B[949] +
//             mat_A[30] * mat_B[981] +
//             mat_A[31] * mat_B[1013];
//  mat_C[22] <= 
//             mat_A[0] * mat_B[22] +
//             mat_A[1] * mat_B[54] +
//             mat_A[2] * mat_B[86] +
//             mat_A[3] * mat_B[118] +
//             mat_A[4] * mat_B[150] +
//             mat_A[5] * mat_B[182] +
//             mat_A[6] * mat_B[214] +
//             mat_A[7] * mat_B[246] +
//             mat_A[8] * mat_B[278] +
//             mat_A[9] * mat_B[310] +
//             mat_A[10] * mat_B[342] +
//             mat_A[11] * mat_B[374] +
//             mat_A[12] * mat_B[406] +
//             mat_A[13] * mat_B[438] +
//             mat_A[14] * mat_B[470] +
//             mat_A[15] * mat_B[502] +
//             mat_A[16] * mat_B[534] +
//             mat_A[17] * mat_B[566] +
//             mat_A[18] * mat_B[598] +
//             mat_A[19] * mat_B[630] +
//             mat_A[20] * mat_B[662] +
//             mat_A[21] * mat_B[694] +
//             mat_A[22] * mat_B[726] +
//             mat_A[23] * mat_B[758] +
//             mat_A[24] * mat_B[790] +
//             mat_A[25] * mat_B[822] +
//             mat_A[26] * mat_B[854] +
//             mat_A[27] * mat_B[886] +
//             mat_A[28] * mat_B[918] +
//             mat_A[29] * mat_B[950] +
//             mat_A[30] * mat_B[982] +
//             mat_A[31] * mat_B[1014];
//  mat_C[23] <= 
//             mat_A[0] * mat_B[23] +
//             mat_A[1] * mat_B[55] +
//             mat_A[2] * mat_B[87] +
//             mat_A[3] * mat_B[119] +
//             mat_A[4] * mat_B[151] +
//             mat_A[5] * mat_B[183] +
//             mat_A[6] * mat_B[215] +
//             mat_A[7] * mat_B[247] +
//             mat_A[8] * mat_B[279] +
//             mat_A[9] * mat_B[311] +
//             mat_A[10] * mat_B[343] +
//             mat_A[11] * mat_B[375] +
//             mat_A[12] * mat_B[407] +
//             mat_A[13] * mat_B[439] +
//             mat_A[14] * mat_B[471] +
//             mat_A[15] * mat_B[503] +
//             mat_A[16] * mat_B[535] +
//             mat_A[17] * mat_B[567] +
//             mat_A[18] * mat_B[599] +
//             mat_A[19] * mat_B[631] +
//             mat_A[20] * mat_B[663] +
//             mat_A[21] * mat_B[695] +
//             mat_A[22] * mat_B[727] +
//             mat_A[23] * mat_B[759] +
//             mat_A[24] * mat_B[791] +
//             mat_A[25] * mat_B[823] +
//             mat_A[26] * mat_B[855] +
//             mat_A[27] * mat_B[887] +
//             mat_A[28] * mat_B[919] +
//             mat_A[29] * mat_B[951] +
//             mat_A[30] * mat_B[983] +
//             mat_A[31] * mat_B[1015];
//  mat_C[24] <= 
//             mat_A[0] * mat_B[24] +
//             mat_A[1] * mat_B[56] +
//             mat_A[2] * mat_B[88] +
//             mat_A[3] * mat_B[120] +
//             mat_A[4] * mat_B[152] +
//             mat_A[5] * mat_B[184] +
//             mat_A[6] * mat_B[216] +
//             mat_A[7] * mat_B[248] +
//             mat_A[8] * mat_B[280] +
//             mat_A[9] * mat_B[312] +
//             mat_A[10] * mat_B[344] +
//             mat_A[11] * mat_B[376] +
//             mat_A[12] * mat_B[408] +
//             mat_A[13] * mat_B[440] +
//             mat_A[14] * mat_B[472] +
//             mat_A[15] * mat_B[504] +
//             mat_A[16] * mat_B[536] +
//             mat_A[17] * mat_B[568] +
//             mat_A[18] * mat_B[600] +
//             mat_A[19] * mat_B[632] +
//             mat_A[20] * mat_B[664] +
//             mat_A[21] * mat_B[696] +
//             mat_A[22] * mat_B[728] +
//             mat_A[23] * mat_B[760] +
//             mat_A[24] * mat_B[792] +
//             mat_A[25] * mat_B[824] +
//             mat_A[26] * mat_B[856] +
//             mat_A[27] * mat_B[888] +
//             mat_A[28] * mat_B[920] +
//             mat_A[29] * mat_B[952] +
//             mat_A[30] * mat_B[984] +
//             mat_A[31] * mat_B[1016];
//  mat_C[25] <= 
//             mat_A[0] * mat_B[25] +
//             mat_A[1] * mat_B[57] +
//             mat_A[2] * mat_B[89] +
//             mat_A[3] * mat_B[121] +
//             mat_A[4] * mat_B[153] +
//             mat_A[5] * mat_B[185] +
//             mat_A[6] * mat_B[217] +
//             mat_A[7] * mat_B[249] +
//             mat_A[8] * mat_B[281] +
//             mat_A[9] * mat_B[313] +
//             mat_A[10] * mat_B[345] +
//             mat_A[11] * mat_B[377] +
//             mat_A[12] * mat_B[409] +
//             mat_A[13] * mat_B[441] +
//             mat_A[14] * mat_B[473] +
//             mat_A[15] * mat_B[505] +
//             mat_A[16] * mat_B[537] +
//             mat_A[17] * mat_B[569] +
//             mat_A[18] * mat_B[601] +
//             mat_A[19] * mat_B[633] +
//             mat_A[20] * mat_B[665] +
//             mat_A[21] * mat_B[697] +
//             mat_A[22] * mat_B[729] +
//             mat_A[23] * mat_B[761] +
//             mat_A[24] * mat_B[793] +
//             mat_A[25] * mat_B[825] +
//             mat_A[26] * mat_B[857] +
//             mat_A[27] * mat_B[889] +
//             mat_A[28] * mat_B[921] +
//             mat_A[29] * mat_B[953] +
//             mat_A[30] * mat_B[985] +
//             mat_A[31] * mat_B[1017];
//  mat_C[26] <= 
//             mat_A[0] * mat_B[26] +
//             mat_A[1] * mat_B[58] +
//             mat_A[2] * mat_B[90] +
//             mat_A[3] * mat_B[122] +
//             mat_A[4] * mat_B[154] +
//             mat_A[5] * mat_B[186] +
//             mat_A[6] * mat_B[218] +
//             mat_A[7] * mat_B[250] +
//             mat_A[8] * mat_B[282] +
//             mat_A[9] * mat_B[314] +
//             mat_A[10] * mat_B[346] +
//             mat_A[11] * mat_B[378] +
//             mat_A[12] * mat_B[410] +
//             mat_A[13] * mat_B[442] +
//             mat_A[14] * mat_B[474] +
//             mat_A[15] * mat_B[506] +
//             mat_A[16] * mat_B[538] +
//             mat_A[17] * mat_B[570] +
//             mat_A[18] * mat_B[602] +
//             mat_A[19] * mat_B[634] +
//             mat_A[20] * mat_B[666] +
//             mat_A[21] * mat_B[698] +
//             mat_A[22] * mat_B[730] +
//             mat_A[23] * mat_B[762] +
//             mat_A[24] * mat_B[794] +
//             mat_A[25] * mat_B[826] +
//             mat_A[26] * mat_B[858] +
//             mat_A[27] * mat_B[890] +
//             mat_A[28] * mat_B[922] +
//             mat_A[29] * mat_B[954] +
//             mat_A[30] * mat_B[986] +
//             mat_A[31] * mat_B[1018];
//  mat_C[27] <= 
//             mat_A[0] * mat_B[27] +
//             mat_A[1] * mat_B[59] +
//             mat_A[2] * mat_B[91] +
//             mat_A[3] * mat_B[123] +
//             mat_A[4] * mat_B[155] +
//             mat_A[5] * mat_B[187] +
//             mat_A[6] * mat_B[219] +
//             mat_A[7] * mat_B[251] +
//             mat_A[8] * mat_B[283] +
//             mat_A[9] * mat_B[315] +
//             mat_A[10] * mat_B[347] +
//             mat_A[11] * mat_B[379] +
//             mat_A[12] * mat_B[411] +
//             mat_A[13] * mat_B[443] +
//             mat_A[14] * mat_B[475] +
//             mat_A[15] * mat_B[507] +
//             mat_A[16] * mat_B[539] +
//             mat_A[17] * mat_B[571] +
//             mat_A[18] * mat_B[603] +
//             mat_A[19] * mat_B[635] +
//             mat_A[20] * mat_B[667] +
//             mat_A[21] * mat_B[699] +
//             mat_A[22] * mat_B[731] +
//             mat_A[23] * mat_B[763] +
//             mat_A[24] * mat_B[795] +
//             mat_A[25] * mat_B[827] +
//             mat_A[26] * mat_B[859] +
//             mat_A[27] * mat_B[891] +
//             mat_A[28] * mat_B[923] +
//             mat_A[29] * mat_B[955] +
//             mat_A[30] * mat_B[987] +
//             mat_A[31] * mat_B[1019];
//  mat_C[28] <= 
//             mat_A[0] * mat_B[28] +
//             mat_A[1] * mat_B[60] +
//             mat_A[2] * mat_B[92] +
//             mat_A[3] * mat_B[124] +
//             mat_A[4] * mat_B[156] +
//             mat_A[5] * mat_B[188] +
//             mat_A[6] * mat_B[220] +
//             mat_A[7] * mat_B[252] +
//             mat_A[8] * mat_B[284] +
//             mat_A[9] * mat_B[316] +
//             mat_A[10] * mat_B[348] +
//             mat_A[11] * mat_B[380] +
//             mat_A[12] * mat_B[412] +
//             mat_A[13] * mat_B[444] +
//             mat_A[14] * mat_B[476] +
//             mat_A[15] * mat_B[508] +
//             mat_A[16] * mat_B[540] +
//             mat_A[17] * mat_B[572] +
//             mat_A[18] * mat_B[604] +
//             mat_A[19] * mat_B[636] +
//             mat_A[20] * mat_B[668] +
//             mat_A[21] * mat_B[700] +
//             mat_A[22] * mat_B[732] +
//             mat_A[23] * mat_B[764] +
//             mat_A[24] * mat_B[796] +
//             mat_A[25] * mat_B[828] +
//             mat_A[26] * mat_B[860] +
//             mat_A[27] * mat_B[892] +
//             mat_A[28] * mat_B[924] +
//             mat_A[29] * mat_B[956] +
//             mat_A[30] * mat_B[988] +
//             mat_A[31] * mat_B[1020];
//  mat_C[29] <= 
//             mat_A[0] * mat_B[29] +
//             mat_A[1] * mat_B[61] +
//             mat_A[2] * mat_B[93] +
//             mat_A[3] * mat_B[125] +
//             mat_A[4] * mat_B[157] +
//             mat_A[5] * mat_B[189] +
//             mat_A[6] * mat_B[221] +
//             mat_A[7] * mat_B[253] +
//             mat_A[8] * mat_B[285] +
//             mat_A[9] * mat_B[317] +
//             mat_A[10] * mat_B[349] +
//             mat_A[11] * mat_B[381] +
//             mat_A[12] * mat_B[413] +
//             mat_A[13] * mat_B[445] +
//             mat_A[14] * mat_B[477] +
//             mat_A[15] * mat_B[509] +
//             mat_A[16] * mat_B[541] +
//             mat_A[17] * mat_B[573] +
//             mat_A[18] * mat_B[605] +
//             mat_A[19] * mat_B[637] +
//             mat_A[20] * mat_B[669] +
//             mat_A[21] * mat_B[701] +
//             mat_A[22] * mat_B[733] +
//             mat_A[23] * mat_B[765] +
//             mat_A[24] * mat_B[797] +
//             mat_A[25] * mat_B[829] +
//             mat_A[26] * mat_B[861] +
//             mat_A[27] * mat_B[893] +
//             mat_A[28] * mat_B[925] +
//             mat_A[29] * mat_B[957] +
//             mat_A[30] * mat_B[989] +
//             mat_A[31] * mat_B[1021];
//  mat_C[30] <= 
//             mat_A[0] * mat_B[30] +
//             mat_A[1] * mat_B[62] +
//             mat_A[2] * mat_B[94] +
//             mat_A[3] * mat_B[126] +
//             mat_A[4] * mat_B[158] +
//             mat_A[5] * mat_B[190] +
//             mat_A[6] * mat_B[222] +
//             mat_A[7] * mat_B[254] +
//             mat_A[8] * mat_B[286] +
//             mat_A[9] * mat_B[318] +
//             mat_A[10] * mat_B[350] +
//             mat_A[11] * mat_B[382] +
//             mat_A[12] * mat_B[414] +
//             mat_A[13] * mat_B[446] +
//             mat_A[14] * mat_B[478] +
//             mat_A[15] * mat_B[510] +
//             mat_A[16] * mat_B[542] +
//             mat_A[17] * mat_B[574] +
//             mat_A[18] * mat_B[606] +
//             mat_A[19] * mat_B[638] +
//             mat_A[20] * mat_B[670] +
//             mat_A[21] * mat_B[702] +
//             mat_A[22] * mat_B[734] +
//             mat_A[23] * mat_B[766] +
//             mat_A[24] * mat_B[798] +
//             mat_A[25] * mat_B[830] +
//             mat_A[26] * mat_B[862] +
//             mat_A[27] * mat_B[894] +
//             mat_A[28] * mat_B[926] +
//             mat_A[29] * mat_B[958] +
//             mat_A[30] * mat_B[990] +
//             mat_A[31] * mat_B[1022];
//  mat_C[31] <= 
//             mat_A[0] * mat_B[31] +
//             mat_A[1] * mat_B[63] +
//             mat_A[2] * mat_B[95] +
//             mat_A[3] * mat_B[127] +
//             mat_A[4] * mat_B[159] +
//             mat_A[5] * mat_B[191] +
//             mat_A[6] * mat_B[223] +
//             mat_A[7] * mat_B[255] +
//             mat_A[8] * mat_B[287] +
//             mat_A[9] * mat_B[319] +
//             mat_A[10] * mat_B[351] +
//             mat_A[11] * mat_B[383] +
//             mat_A[12] * mat_B[415] +
//             mat_A[13] * mat_B[447] +
//             mat_A[14] * mat_B[479] +
//             mat_A[15] * mat_B[511] +
//             mat_A[16] * mat_B[543] +
//             mat_A[17] * mat_B[575] +
//             mat_A[18] * mat_B[607] +
//             mat_A[19] * mat_B[639] +
//             mat_A[20] * mat_B[671] +
//             mat_A[21] * mat_B[703] +
//             mat_A[22] * mat_B[735] +
//             mat_A[23] * mat_B[767] +
//             mat_A[24] * mat_B[799] +
//             mat_A[25] * mat_B[831] +
//             mat_A[26] * mat_B[863] +
//             mat_A[27] * mat_B[895] +
//             mat_A[28] * mat_B[927] +
//             mat_A[29] * mat_B[959] +
//             mat_A[30] * mat_B[991] +
//             mat_A[31] * mat_B[1023];
//  mat_C[32] <= 
//             mat_A[32] * mat_B[0] +
//             mat_A[33] * mat_B[32] +
//             mat_A[34] * mat_B[64] +
//             mat_A[35] * mat_B[96] +
//             mat_A[36] * mat_B[128] +
//             mat_A[37] * mat_B[160] +
//             mat_A[38] * mat_B[192] +
//             mat_A[39] * mat_B[224] +
//             mat_A[40] * mat_B[256] +
//             mat_A[41] * mat_B[288] +
//             mat_A[42] * mat_B[320] +
//             mat_A[43] * mat_B[352] +
//             mat_A[44] * mat_B[384] +
//             mat_A[45] * mat_B[416] +
//             mat_A[46] * mat_B[448] +
//             mat_A[47] * mat_B[480] +
//             mat_A[48] * mat_B[512] +
//             mat_A[49] * mat_B[544] +
//             mat_A[50] * mat_B[576] +
//             mat_A[51] * mat_B[608] +
//             mat_A[52] * mat_B[640] +
//             mat_A[53] * mat_B[672] +
//             mat_A[54] * mat_B[704] +
//             mat_A[55] * mat_B[736] +
//             mat_A[56] * mat_B[768] +
//             mat_A[57] * mat_B[800] +
//             mat_A[58] * mat_B[832] +
//             mat_A[59] * mat_B[864] +
//             mat_A[60] * mat_B[896] +
//             mat_A[61] * mat_B[928] +
//             mat_A[62] * mat_B[960] +
//             mat_A[63] * mat_B[992];
//  mat_C[33] <= 
//             mat_A[32] * mat_B[1] +
//             mat_A[33] * mat_B[33] +
//             mat_A[34] * mat_B[65] +
//             mat_A[35] * mat_B[97] +
//             mat_A[36] * mat_B[129] +
//             mat_A[37] * mat_B[161] +
//             mat_A[38] * mat_B[193] +
//             mat_A[39] * mat_B[225] +
//             mat_A[40] * mat_B[257] +
//             mat_A[41] * mat_B[289] +
//             mat_A[42] * mat_B[321] +
//             mat_A[43] * mat_B[353] +
//             mat_A[44] * mat_B[385] +
//             mat_A[45] * mat_B[417] +
//             mat_A[46] * mat_B[449] +
//             mat_A[47] * mat_B[481] +
//             mat_A[48] * mat_B[513] +
//             mat_A[49] * mat_B[545] +
//             mat_A[50] * mat_B[577] +
//             mat_A[51] * mat_B[609] +
//             mat_A[52] * mat_B[641] +
//             mat_A[53] * mat_B[673] +
//             mat_A[54] * mat_B[705] +
//             mat_A[55] * mat_B[737] +
//             mat_A[56] * mat_B[769] +
//             mat_A[57] * mat_B[801] +
//             mat_A[58] * mat_B[833] +
//             mat_A[59] * mat_B[865] +
//             mat_A[60] * mat_B[897] +
//             mat_A[61] * mat_B[929] +
//             mat_A[62] * mat_B[961] +
//             mat_A[63] * mat_B[993];
//  mat_C[34] <= 
//             mat_A[32] * mat_B[2] +
//             mat_A[33] * mat_B[34] +
//             mat_A[34] * mat_B[66] +
//             mat_A[35] * mat_B[98] +
//             mat_A[36] * mat_B[130] +
//             mat_A[37] * mat_B[162] +
//             mat_A[38] * mat_B[194] +
//             mat_A[39] * mat_B[226] +
//             mat_A[40] * mat_B[258] +
//             mat_A[41] * mat_B[290] +
//             mat_A[42] * mat_B[322] +
//             mat_A[43] * mat_B[354] +
//             mat_A[44] * mat_B[386] +
//             mat_A[45] * mat_B[418] +
//             mat_A[46] * mat_B[450] +
//             mat_A[47] * mat_B[482] +
//             mat_A[48] * mat_B[514] +
//             mat_A[49] * mat_B[546] +
//             mat_A[50] * mat_B[578] +
//             mat_A[51] * mat_B[610] +
//             mat_A[52] * mat_B[642] +
//             mat_A[53] * mat_B[674] +
//             mat_A[54] * mat_B[706] +
//             mat_A[55] * mat_B[738] +
//             mat_A[56] * mat_B[770] +
//             mat_A[57] * mat_B[802] +
//             mat_A[58] * mat_B[834] +
//             mat_A[59] * mat_B[866] +
//             mat_A[60] * mat_B[898] +
//             mat_A[61] * mat_B[930] +
//             mat_A[62] * mat_B[962] +
//             mat_A[63] * mat_B[994];
//  mat_C[35] <= 
//             mat_A[32] * mat_B[3] +
//             mat_A[33] * mat_B[35] +
//             mat_A[34] * mat_B[67] +
//             mat_A[35] * mat_B[99] +
//             mat_A[36] * mat_B[131] +
//             mat_A[37] * mat_B[163] +
//             mat_A[38] * mat_B[195] +
//             mat_A[39] * mat_B[227] +
//             mat_A[40] * mat_B[259] +
//             mat_A[41] * mat_B[291] +
//             mat_A[42] * mat_B[323] +
//             mat_A[43] * mat_B[355] +
//             mat_A[44] * mat_B[387] +
//             mat_A[45] * mat_B[419] +
//             mat_A[46] * mat_B[451] +
//             mat_A[47] * mat_B[483] +
//             mat_A[48] * mat_B[515] +
//             mat_A[49] * mat_B[547] +
//             mat_A[50] * mat_B[579] +
//             mat_A[51] * mat_B[611] +
//             mat_A[52] * mat_B[643] +
//             mat_A[53] * mat_B[675] +
//             mat_A[54] * mat_B[707] +
//             mat_A[55] * mat_B[739] +
//             mat_A[56] * mat_B[771] +
//             mat_A[57] * mat_B[803] +
//             mat_A[58] * mat_B[835] +
//             mat_A[59] * mat_B[867] +
//             mat_A[60] * mat_B[899] +
//             mat_A[61] * mat_B[931] +
//             mat_A[62] * mat_B[963] +
//             mat_A[63] * mat_B[995];
//  mat_C[36] <= 
//             mat_A[32] * mat_B[4] +
//             mat_A[33] * mat_B[36] +
//             mat_A[34] * mat_B[68] +
//             mat_A[35] * mat_B[100] +
//             mat_A[36] * mat_B[132] +
//             mat_A[37] * mat_B[164] +
//             mat_A[38] * mat_B[196] +
//             mat_A[39] * mat_B[228] +
//             mat_A[40] * mat_B[260] +
//             mat_A[41] * mat_B[292] +
//             mat_A[42] * mat_B[324] +
//             mat_A[43] * mat_B[356] +
//             mat_A[44] * mat_B[388] +
//             mat_A[45] * mat_B[420] +
//             mat_A[46] * mat_B[452] +
//             mat_A[47] * mat_B[484] +
//             mat_A[48] * mat_B[516] +
//             mat_A[49] * mat_B[548] +
//             mat_A[50] * mat_B[580] +
//             mat_A[51] * mat_B[612] +
//             mat_A[52] * mat_B[644] +
//             mat_A[53] * mat_B[676] +
//             mat_A[54] * mat_B[708] +
//             mat_A[55] * mat_B[740] +
//             mat_A[56] * mat_B[772] +
//             mat_A[57] * mat_B[804] +
//             mat_A[58] * mat_B[836] +
//             mat_A[59] * mat_B[868] +
//             mat_A[60] * mat_B[900] +
//             mat_A[61] * mat_B[932] +
//             mat_A[62] * mat_B[964] +
//             mat_A[63] * mat_B[996];
//  mat_C[37] <= 
//             mat_A[32] * mat_B[5] +
//             mat_A[33] * mat_B[37] +
//             mat_A[34] * mat_B[69] +
//             mat_A[35] * mat_B[101] +
//             mat_A[36] * mat_B[133] +
//             mat_A[37] * mat_B[165] +
//             mat_A[38] * mat_B[197] +
//             mat_A[39] * mat_B[229] +
//             mat_A[40] * mat_B[261] +
//             mat_A[41] * mat_B[293] +
//             mat_A[42] * mat_B[325] +
//             mat_A[43] * mat_B[357] +
//             mat_A[44] * mat_B[389] +
//             mat_A[45] * mat_B[421] +
//             mat_A[46] * mat_B[453] +
//             mat_A[47] * mat_B[485] +
//             mat_A[48] * mat_B[517] +
//             mat_A[49] * mat_B[549] +
//             mat_A[50] * mat_B[581] +
//             mat_A[51] * mat_B[613] +
//             mat_A[52] * mat_B[645] +
//             mat_A[53] * mat_B[677] +
//             mat_A[54] * mat_B[709] +
//             mat_A[55] * mat_B[741] +
//             mat_A[56] * mat_B[773] +
//             mat_A[57] * mat_B[805] +
//             mat_A[58] * mat_B[837] +
//             mat_A[59] * mat_B[869] +
//             mat_A[60] * mat_B[901] +
//             mat_A[61] * mat_B[933] +
//             mat_A[62] * mat_B[965] +
//             mat_A[63] * mat_B[997];
//  mat_C[38] <= 
//             mat_A[32] * mat_B[6] +
//             mat_A[33] * mat_B[38] +
//             mat_A[34] * mat_B[70] +
//             mat_A[35] * mat_B[102] +
//             mat_A[36] * mat_B[134] +
//             mat_A[37] * mat_B[166] +
//             mat_A[38] * mat_B[198] +
//             mat_A[39] * mat_B[230] +
//             mat_A[40] * mat_B[262] +
//             mat_A[41] * mat_B[294] +
//             mat_A[42] * mat_B[326] +
//             mat_A[43] * mat_B[358] +
//             mat_A[44] * mat_B[390] +
//             mat_A[45] * mat_B[422] +
//             mat_A[46] * mat_B[454] +
//             mat_A[47] * mat_B[486] +
//             mat_A[48] * mat_B[518] +
//             mat_A[49] * mat_B[550] +
//             mat_A[50] * mat_B[582] +
//             mat_A[51] * mat_B[614] +
//             mat_A[52] * mat_B[646] +
//             mat_A[53] * mat_B[678] +
//             mat_A[54] * mat_B[710] +
//             mat_A[55] * mat_B[742] +
//             mat_A[56] * mat_B[774] +
//             mat_A[57] * mat_B[806] +
//             mat_A[58] * mat_B[838] +
//             mat_A[59] * mat_B[870] +
//             mat_A[60] * mat_B[902] +
//             mat_A[61] * mat_B[934] +
//             mat_A[62] * mat_B[966] +
//             mat_A[63] * mat_B[998];
//  mat_C[39] <= 
//             mat_A[32] * mat_B[7] +
//             mat_A[33] * mat_B[39] +
//             mat_A[34] * mat_B[71] +
//             mat_A[35] * mat_B[103] +
//             mat_A[36] * mat_B[135] +
//             mat_A[37] * mat_B[167] +
//             mat_A[38] * mat_B[199] +
//             mat_A[39] * mat_B[231] +
//             mat_A[40] * mat_B[263] +
//             mat_A[41] * mat_B[295] +
//             mat_A[42] * mat_B[327] +
//             mat_A[43] * mat_B[359] +
//             mat_A[44] * mat_B[391] +
//             mat_A[45] * mat_B[423] +
//             mat_A[46] * mat_B[455] +
//             mat_A[47] * mat_B[487] +
//             mat_A[48] * mat_B[519] +
//             mat_A[49] * mat_B[551] +
//             mat_A[50] * mat_B[583] +
//             mat_A[51] * mat_B[615] +
//             mat_A[52] * mat_B[647] +
//             mat_A[53] * mat_B[679] +
//             mat_A[54] * mat_B[711] +
//             mat_A[55] * mat_B[743] +
//             mat_A[56] * mat_B[775] +
//             mat_A[57] * mat_B[807] +
//             mat_A[58] * mat_B[839] +
//             mat_A[59] * mat_B[871] +
//             mat_A[60] * mat_B[903] +
//             mat_A[61] * mat_B[935] +
//             mat_A[62] * mat_B[967] +
//             mat_A[63] * mat_B[999];
//  mat_C[40] <= 
//             mat_A[32] * mat_B[8] +
//             mat_A[33] * mat_B[40] +
//             mat_A[34] * mat_B[72] +
//             mat_A[35] * mat_B[104] +
//             mat_A[36] * mat_B[136] +
//             mat_A[37] * mat_B[168] +
//             mat_A[38] * mat_B[200] +
//             mat_A[39] * mat_B[232] +
//             mat_A[40] * mat_B[264] +
//             mat_A[41] * mat_B[296] +
//             mat_A[42] * mat_B[328] +
//             mat_A[43] * mat_B[360] +
//             mat_A[44] * mat_B[392] +
//             mat_A[45] * mat_B[424] +
//             mat_A[46] * mat_B[456] +
//             mat_A[47] * mat_B[488] +
//             mat_A[48] * mat_B[520] +
//             mat_A[49] * mat_B[552] +
//             mat_A[50] * mat_B[584] +
//             mat_A[51] * mat_B[616] +
//             mat_A[52] * mat_B[648] +
//             mat_A[53] * mat_B[680] +
//             mat_A[54] * mat_B[712] +
//             mat_A[55] * mat_B[744] +
//             mat_A[56] * mat_B[776] +
//             mat_A[57] * mat_B[808] +
//             mat_A[58] * mat_B[840] +
//             mat_A[59] * mat_B[872] +
//             mat_A[60] * mat_B[904] +
//             mat_A[61] * mat_B[936] +
//             mat_A[62] * mat_B[968] +
//             mat_A[63] * mat_B[1000];
//  mat_C[41] <= 
//             mat_A[32] * mat_B[9] +
//             mat_A[33] * mat_B[41] +
//             mat_A[34] * mat_B[73] +
//             mat_A[35] * mat_B[105] +
//             mat_A[36] * mat_B[137] +
//             mat_A[37] * mat_B[169] +
//             mat_A[38] * mat_B[201] +
//             mat_A[39] * mat_B[233] +
//             mat_A[40] * mat_B[265] +
//             mat_A[41] * mat_B[297] +
//             mat_A[42] * mat_B[329] +
//             mat_A[43] * mat_B[361] +
//             mat_A[44] * mat_B[393] +
//             mat_A[45] * mat_B[425] +
//             mat_A[46] * mat_B[457] +
//             mat_A[47] * mat_B[489] +
//             mat_A[48] * mat_B[521] +
//             mat_A[49] * mat_B[553] +
//             mat_A[50] * mat_B[585] +
//             mat_A[51] * mat_B[617] +
//             mat_A[52] * mat_B[649] +
//             mat_A[53] * mat_B[681] +
//             mat_A[54] * mat_B[713] +
//             mat_A[55] * mat_B[745] +
//             mat_A[56] * mat_B[777] +
//             mat_A[57] * mat_B[809] +
//             mat_A[58] * mat_B[841] +
//             mat_A[59] * mat_B[873] +
//             mat_A[60] * mat_B[905] +
//             mat_A[61] * mat_B[937] +
//             mat_A[62] * mat_B[969] +
//             mat_A[63] * mat_B[1001];
//  mat_C[42] <= 
//             mat_A[32] * mat_B[10] +
//             mat_A[33] * mat_B[42] +
//             mat_A[34] * mat_B[74] +
//             mat_A[35] * mat_B[106] +
//             mat_A[36] * mat_B[138] +
//             mat_A[37] * mat_B[170] +
//             mat_A[38] * mat_B[202] +
//             mat_A[39] * mat_B[234] +
//             mat_A[40] * mat_B[266] +
//             mat_A[41] * mat_B[298] +
//             mat_A[42] * mat_B[330] +
//             mat_A[43] * mat_B[362] +
//             mat_A[44] * mat_B[394] +
//             mat_A[45] * mat_B[426] +
//             mat_A[46] * mat_B[458] +
//             mat_A[47] * mat_B[490] +
//             mat_A[48] * mat_B[522] +
//             mat_A[49] * mat_B[554] +
//             mat_A[50] * mat_B[586] +
//             mat_A[51] * mat_B[618] +
//             mat_A[52] * mat_B[650] +
//             mat_A[53] * mat_B[682] +
//             mat_A[54] * mat_B[714] +
//             mat_A[55] * mat_B[746] +
//             mat_A[56] * mat_B[778] +
//             mat_A[57] * mat_B[810] +
//             mat_A[58] * mat_B[842] +
//             mat_A[59] * mat_B[874] +
//             mat_A[60] * mat_B[906] +
//             mat_A[61] * mat_B[938] +
//             mat_A[62] * mat_B[970] +
//             mat_A[63] * mat_B[1002];
//  mat_C[43] <= 
//             mat_A[32] * mat_B[11] +
//             mat_A[33] * mat_B[43] +
//             mat_A[34] * mat_B[75] +
//             mat_A[35] * mat_B[107] +
//             mat_A[36] * mat_B[139] +
//             mat_A[37] * mat_B[171] +
//             mat_A[38] * mat_B[203] +
//             mat_A[39] * mat_B[235] +
//             mat_A[40] * mat_B[267] +
//             mat_A[41] * mat_B[299] +
//             mat_A[42] * mat_B[331] +
//             mat_A[43] * mat_B[363] +
//             mat_A[44] * mat_B[395] +
//             mat_A[45] * mat_B[427] +
//             mat_A[46] * mat_B[459] +
//             mat_A[47] * mat_B[491] +
//             mat_A[48] * mat_B[523] +
//             mat_A[49] * mat_B[555] +
//             mat_A[50] * mat_B[587] +
//             mat_A[51] * mat_B[619] +
//             mat_A[52] * mat_B[651] +
//             mat_A[53] * mat_B[683] +
//             mat_A[54] * mat_B[715] +
//             mat_A[55] * mat_B[747] +
//             mat_A[56] * mat_B[779] +
//             mat_A[57] * mat_B[811] +
//             mat_A[58] * mat_B[843] +
//             mat_A[59] * mat_B[875] +
//             mat_A[60] * mat_B[907] +
//             mat_A[61] * mat_B[939] +
//             mat_A[62] * mat_B[971] +
//             mat_A[63] * mat_B[1003];
//  mat_C[44] <= 
//             mat_A[32] * mat_B[12] +
//             mat_A[33] * mat_B[44] +
//             mat_A[34] * mat_B[76] +
//             mat_A[35] * mat_B[108] +
//             mat_A[36] * mat_B[140] +
//             mat_A[37] * mat_B[172] +
//             mat_A[38] * mat_B[204] +
//             mat_A[39] * mat_B[236] +
//             mat_A[40] * mat_B[268] +
//             mat_A[41] * mat_B[300] +
//             mat_A[42] * mat_B[332] +
//             mat_A[43] * mat_B[364] +
//             mat_A[44] * mat_B[396] +
//             mat_A[45] * mat_B[428] +
//             mat_A[46] * mat_B[460] +
//             mat_A[47] * mat_B[492] +
//             mat_A[48] * mat_B[524] +
//             mat_A[49] * mat_B[556] +
//             mat_A[50] * mat_B[588] +
//             mat_A[51] * mat_B[620] +
//             mat_A[52] * mat_B[652] +
//             mat_A[53] * mat_B[684] +
//             mat_A[54] * mat_B[716] +
//             mat_A[55] * mat_B[748] +
//             mat_A[56] * mat_B[780] +
//             mat_A[57] * mat_B[812] +
//             mat_A[58] * mat_B[844] +
//             mat_A[59] * mat_B[876] +
//             mat_A[60] * mat_B[908] +
//             mat_A[61] * mat_B[940] +
//             mat_A[62] * mat_B[972] +
//             mat_A[63] * mat_B[1004];
//  mat_C[45] <= 
//             mat_A[32] * mat_B[13] +
//             mat_A[33] * mat_B[45] +
//             mat_A[34] * mat_B[77] +
//             mat_A[35] * mat_B[109] +
//             mat_A[36] * mat_B[141] +
//             mat_A[37] * mat_B[173] +
//             mat_A[38] * mat_B[205] +
//             mat_A[39] * mat_B[237] +
//             mat_A[40] * mat_B[269] +
//             mat_A[41] * mat_B[301] +
//             mat_A[42] * mat_B[333] +
//             mat_A[43] * mat_B[365] +
//             mat_A[44] * mat_B[397] +
//             mat_A[45] * mat_B[429] +
//             mat_A[46] * mat_B[461] +
//             mat_A[47] * mat_B[493] +
//             mat_A[48] * mat_B[525] +
//             mat_A[49] * mat_B[557] +
//             mat_A[50] * mat_B[589] +
//             mat_A[51] * mat_B[621] +
//             mat_A[52] * mat_B[653] +
//             mat_A[53] * mat_B[685] +
//             mat_A[54] * mat_B[717] +
//             mat_A[55] * mat_B[749] +
//             mat_A[56] * mat_B[781] +
//             mat_A[57] * mat_B[813] +
//             mat_A[58] * mat_B[845] +
//             mat_A[59] * mat_B[877] +
//             mat_A[60] * mat_B[909] +
//             mat_A[61] * mat_B[941] +
//             mat_A[62] * mat_B[973] +
//             mat_A[63] * mat_B[1005];
//  mat_C[46] <= 
//             mat_A[32] * mat_B[14] +
//             mat_A[33] * mat_B[46] +
//             mat_A[34] * mat_B[78] +
//             mat_A[35] * mat_B[110] +
//             mat_A[36] * mat_B[142] +
//             mat_A[37] * mat_B[174] +
//             mat_A[38] * mat_B[206] +
//             mat_A[39] * mat_B[238] +
//             mat_A[40] * mat_B[270] +
//             mat_A[41] * mat_B[302] +
//             mat_A[42] * mat_B[334] +
//             mat_A[43] * mat_B[366] +
//             mat_A[44] * mat_B[398] +
//             mat_A[45] * mat_B[430] +
//             mat_A[46] * mat_B[462] +
//             mat_A[47] * mat_B[494] +
//             mat_A[48] * mat_B[526] +
//             mat_A[49] * mat_B[558] +
//             mat_A[50] * mat_B[590] +
//             mat_A[51] * mat_B[622] +
//             mat_A[52] * mat_B[654] +
//             mat_A[53] * mat_B[686] +
//             mat_A[54] * mat_B[718] +
//             mat_A[55] * mat_B[750] +
//             mat_A[56] * mat_B[782] +
//             mat_A[57] * mat_B[814] +
//             mat_A[58] * mat_B[846] +
//             mat_A[59] * mat_B[878] +
//             mat_A[60] * mat_B[910] +
//             mat_A[61] * mat_B[942] +
//             mat_A[62] * mat_B[974] +
//             mat_A[63] * mat_B[1006];
//  mat_C[47] <= 
//             mat_A[32] * mat_B[15] +
//             mat_A[33] * mat_B[47] +
//             mat_A[34] * mat_B[79] +
//             mat_A[35] * mat_B[111] +
//             mat_A[36] * mat_B[143] +
//             mat_A[37] * mat_B[175] +
//             mat_A[38] * mat_B[207] +
//             mat_A[39] * mat_B[239] +
//             mat_A[40] * mat_B[271] +
//             mat_A[41] * mat_B[303] +
//             mat_A[42] * mat_B[335] +
//             mat_A[43] * mat_B[367] +
//             mat_A[44] * mat_B[399] +
//             mat_A[45] * mat_B[431] +
//             mat_A[46] * mat_B[463] +
//             mat_A[47] * mat_B[495] +
//             mat_A[48] * mat_B[527] +
//             mat_A[49] * mat_B[559] +
//             mat_A[50] * mat_B[591] +
//             mat_A[51] * mat_B[623] +
//             mat_A[52] * mat_B[655] +
//             mat_A[53] * mat_B[687] +
//             mat_A[54] * mat_B[719] +
//             mat_A[55] * mat_B[751] +
//             mat_A[56] * mat_B[783] +
//             mat_A[57] * mat_B[815] +
//             mat_A[58] * mat_B[847] +
//             mat_A[59] * mat_B[879] +
//             mat_A[60] * mat_B[911] +
//             mat_A[61] * mat_B[943] +
//             mat_A[62] * mat_B[975] +
//             mat_A[63] * mat_B[1007];
//  mat_C[48] <= 
//             mat_A[32] * mat_B[16] +
//             mat_A[33] * mat_B[48] +
//             mat_A[34] * mat_B[80] +
//             mat_A[35] * mat_B[112] +
//             mat_A[36] * mat_B[144] +
//             mat_A[37] * mat_B[176] +
//             mat_A[38] * mat_B[208] +
//             mat_A[39] * mat_B[240] +
//             mat_A[40] * mat_B[272] +
//             mat_A[41] * mat_B[304] +
//             mat_A[42] * mat_B[336] +
//             mat_A[43] * mat_B[368] +
//             mat_A[44] * mat_B[400] +
//             mat_A[45] * mat_B[432] +
//             mat_A[46] * mat_B[464] +
//             mat_A[47] * mat_B[496] +
//             mat_A[48] * mat_B[528] +
//             mat_A[49] * mat_B[560] +
//             mat_A[50] * mat_B[592] +
//             mat_A[51] * mat_B[624] +
//             mat_A[52] * mat_B[656] +
//             mat_A[53] * mat_B[688] +
//             mat_A[54] * mat_B[720] +
//             mat_A[55] * mat_B[752] +
//             mat_A[56] * mat_B[784] +
//             mat_A[57] * mat_B[816] +
//             mat_A[58] * mat_B[848] +
//             mat_A[59] * mat_B[880] +
//             mat_A[60] * mat_B[912] +
//             mat_A[61] * mat_B[944] +
//             mat_A[62] * mat_B[976] +
//             mat_A[63] * mat_B[1008];
//  mat_C[49] <= 
//             mat_A[32] * mat_B[17] +
//             mat_A[33] * mat_B[49] +
//             mat_A[34] * mat_B[81] +
//             mat_A[35] * mat_B[113] +
//             mat_A[36] * mat_B[145] +
//             mat_A[37] * mat_B[177] +
//             mat_A[38] * mat_B[209] +
//             mat_A[39] * mat_B[241] +
//             mat_A[40] * mat_B[273] +
//             mat_A[41] * mat_B[305] +
//             mat_A[42] * mat_B[337] +
//             mat_A[43] * mat_B[369] +
//             mat_A[44] * mat_B[401] +
//             mat_A[45] * mat_B[433] +
//             mat_A[46] * mat_B[465] +
//             mat_A[47] * mat_B[497] +
//             mat_A[48] * mat_B[529] +
//             mat_A[49] * mat_B[561] +
//             mat_A[50] * mat_B[593] +
//             mat_A[51] * mat_B[625] +
//             mat_A[52] * mat_B[657] +
//             mat_A[53] * mat_B[689] +
//             mat_A[54] * mat_B[721] +
//             mat_A[55] * mat_B[753] +
//             mat_A[56] * mat_B[785] +
//             mat_A[57] * mat_B[817] +
//             mat_A[58] * mat_B[849] +
//             mat_A[59] * mat_B[881] +
//             mat_A[60] * mat_B[913] +
//             mat_A[61] * mat_B[945] +
//             mat_A[62] * mat_B[977] +
//             mat_A[63] * mat_B[1009];
//  mat_C[50] <= 
//             mat_A[32] * mat_B[18] +
//             mat_A[33] * mat_B[50] +
//             mat_A[34] * mat_B[82] +
//             mat_A[35] * mat_B[114] +
//             mat_A[36] * mat_B[146] +
//             mat_A[37] * mat_B[178] +
//             mat_A[38] * mat_B[210] +
//             mat_A[39] * mat_B[242] +
//             mat_A[40] * mat_B[274] +
//             mat_A[41] * mat_B[306] +
//             mat_A[42] * mat_B[338] +
//             mat_A[43] * mat_B[370] +
//             mat_A[44] * mat_B[402] +
//             mat_A[45] * mat_B[434] +
//             mat_A[46] * mat_B[466] +
//             mat_A[47] * mat_B[498] +
//             mat_A[48] * mat_B[530] +
//             mat_A[49] * mat_B[562] +
//             mat_A[50] * mat_B[594] +
//             mat_A[51] * mat_B[626] +
//             mat_A[52] * mat_B[658] +
//             mat_A[53] * mat_B[690] +
//             mat_A[54] * mat_B[722] +
//             mat_A[55] * mat_B[754] +
//             mat_A[56] * mat_B[786] +
//             mat_A[57] * mat_B[818] +
//             mat_A[58] * mat_B[850] +
//             mat_A[59] * mat_B[882] +
//             mat_A[60] * mat_B[914] +
//             mat_A[61] * mat_B[946] +
//             mat_A[62] * mat_B[978] +
//             mat_A[63] * mat_B[1010];
//  mat_C[51] <= 
//             mat_A[32] * mat_B[19] +
//             mat_A[33] * mat_B[51] +
//             mat_A[34] * mat_B[83] +
//             mat_A[35] * mat_B[115] +
//             mat_A[36] * mat_B[147] +
//             mat_A[37] * mat_B[179] +
//             mat_A[38] * mat_B[211] +
//             mat_A[39] * mat_B[243] +
//             mat_A[40] * mat_B[275] +
//             mat_A[41] * mat_B[307] +
//             mat_A[42] * mat_B[339] +
//             mat_A[43] * mat_B[371] +
//             mat_A[44] * mat_B[403] +
//             mat_A[45] * mat_B[435] +
//             mat_A[46] * mat_B[467] +
//             mat_A[47] * mat_B[499] +
//             mat_A[48] * mat_B[531] +
//             mat_A[49] * mat_B[563] +
//             mat_A[50] * mat_B[595] +
//             mat_A[51] * mat_B[627] +
//             mat_A[52] * mat_B[659] +
//             mat_A[53] * mat_B[691] +
//             mat_A[54] * mat_B[723] +
//             mat_A[55] * mat_B[755] +
//             mat_A[56] * mat_B[787] +
//             mat_A[57] * mat_B[819] +
//             mat_A[58] * mat_B[851] +
//             mat_A[59] * mat_B[883] +
//             mat_A[60] * mat_B[915] +
//             mat_A[61] * mat_B[947] +
//             mat_A[62] * mat_B[979] +
//             mat_A[63] * mat_B[1011];
//  mat_C[52] <= 
//             mat_A[32] * mat_B[20] +
//             mat_A[33] * mat_B[52] +
//             mat_A[34] * mat_B[84] +
//             mat_A[35] * mat_B[116] +
//             mat_A[36] * mat_B[148] +
//             mat_A[37] * mat_B[180] +
//             mat_A[38] * mat_B[212] +
//             mat_A[39] * mat_B[244] +
//             mat_A[40] * mat_B[276] +
//             mat_A[41] * mat_B[308] +
//             mat_A[42] * mat_B[340] +
//             mat_A[43] * mat_B[372] +
//             mat_A[44] * mat_B[404] +
//             mat_A[45] * mat_B[436] +
//             mat_A[46] * mat_B[468] +
//             mat_A[47] * mat_B[500] +
//             mat_A[48] * mat_B[532] +
//             mat_A[49] * mat_B[564] +
//             mat_A[50] * mat_B[596] +
//             mat_A[51] * mat_B[628] +
//             mat_A[52] * mat_B[660] +
//             mat_A[53] * mat_B[692] +
//             mat_A[54] * mat_B[724] +
//             mat_A[55] * mat_B[756] +
//             mat_A[56] * mat_B[788] +
//             mat_A[57] * mat_B[820] +
//             mat_A[58] * mat_B[852] +
//             mat_A[59] * mat_B[884] +
//             mat_A[60] * mat_B[916] +
//             mat_A[61] * mat_B[948] +
//             mat_A[62] * mat_B[980] +
//             mat_A[63] * mat_B[1012];
//  mat_C[53] <= 
//             mat_A[32] * mat_B[21] +
//             mat_A[33] * mat_B[53] +
//             mat_A[34] * mat_B[85] +
//             mat_A[35] * mat_B[117] +
//             mat_A[36] * mat_B[149] +
//             mat_A[37] * mat_B[181] +
//             mat_A[38] * mat_B[213] +
//             mat_A[39] * mat_B[245] +
//             mat_A[40] * mat_B[277] +
//             mat_A[41] * mat_B[309] +
//             mat_A[42] * mat_B[341] +
//             mat_A[43] * mat_B[373] +
//             mat_A[44] * mat_B[405] +
//             mat_A[45] * mat_B[437] +
//             mat_A[46] * mat_B[469] +
//             mat_A[47] * mat_B[501] +
//             mat_A[48] * mat_B[533] +
//             mat_A[49] * mat_B[565] +
//             mat_A[50] * mat_B[597] +
//             mat_A[51] * mat_B[629] +
//             mat_A[52] * mat_B[661] +
//             mat_A[53] * mat_B[693] +
//             mat_A[54] * mat_B[725] +
//             mat_A[55] * mat_B[757] +
//             mat_A[56] * mat_B[789] +
//             mat_A[57] * mat_B[821] +
//             mat_A[58] * mat_B[853] +
//             mat_A[59] * mat_B[885] +
//             mat_A[60] * mat_B[917] +
//             mat_A[61] * mat_B[949] +
//             mat_A[62] * mat_B[981] +
//             mat_A[63] * mat_B[1013];
//  mat_C[54] <= 
//             mat_A[32] * mat_B[22] +
//             mat_A[33] * mat_B[54] +
//             mat_A[34] * mat_B[86] +
//             mat_A[35] * mat_B[118] +
//             mat_A[36] * mat_B[150] +
//             mat_A[37] * mat_B[182] +
//             mat_A[38] * mat_B[214] +
//             mat_A[39] * mat_B[246] +
//             mat_A[40] * mat_B[278] +
//             mat_A[41] * mat_B[310] +
//             mat_A[42] * mat_B[342] +
//             mat_A[43] * mat_B[374] +
//             mat_A[44] * mat_B[406] +
//             mat_A[45] * mat_B[438] +
//             mat_A[46] * mat_B[470] +
//             mat_A[47] * mat_B[502] +
//             mat_A[48] * mat_B[534] +
//             mat_A[49] * mat_B[566] +
//             mat_A[50] * mat_B[598] +
//             mat_A[51] * mat_B[630] +
//             mat_A[52] * mat_B[662] +
//             mat_A[53] * mat_B[694] +
//             mat_A[54] * mat_B[726] +
//             mat_A[55] * mat_B[758] +
//             mat_A[56] * mat_B[790] +
//             mat_A[57] * mat_B[822] +
//             mat_A[58] * mat_B[854] +
//             mat_A[59] * mat_B[886] +
//             mat_A[60] * mat_B[918] +
//             mat_A[61] * mat_B[950] +
//             mat_A[62] * mat_B[982] +
//             mat_A[63] * mat_B[1014];
//  mat_C[55] <= 
//             mat_A[32] * mat_B[23] +
//             mat_A[33] * mat_B[55] +
//             mat_A[34] * mat_B[87] +
//             mat_A[35] * mat_B[119] +
//             mat_A[36] * mat_B[151] +
//             mat_A[37] * mat_B[183] +
//             mat_A[38] * mat_B[215] +
//             mat_A[39] * mat_B[247] +
//             mat_A[40] * mat_B[279] +
//             mat_A[41] * mat_B[311] +
//             mat_A[42] * mat_B[343] +
//             mat_A[43] * mat_B[375] +
//             mat_A[44] * mat_B[407] +
//             mat_A[45] * mat_B[439] +
//             mat_A[46] * mat_B[471] +
//             mat_A[47] * mat_B[503] +
//             mat_A[48] * mat_B[535] +
//             mat_A[49] * mat_B[567] +
//             mat_A[50] * mat_B[599] +
//             mat_A[51] * mat_B[631] +
//             mat_A[52] * mat_B[663] +
//             mat_A[53] * mat_B[695] +
//             mat_A[54] * mat_B[727] +
//             mat_A[55] * mat_B[759] +
//             mat_A[56] * mat_B[791] +
//             mat_A[57] * mat_B[823] +
//             mat_A[58] * mat_B[855] +
//             mat_A[59] * mat_B[887] +
//             mat_A[60] * mat_B[919] +
//             mat_A[61] * mat_B[951] +
//             mat_A[62] * mat_B[983] +
//             mat_A[63] * mat_B[1015];
//  mat_C[56] <= 
//             mat_A[32] * mat_B[24] +
//             mat_A[33] * mat_B[56] +
//             mat_A[34] * mat_B[88] +
//             mat_A[35] * mat_B[120] +
//             mat_A[36] * mat_B[152] +
//             mat_A[37] * mat_B[184] +
//             mat_A[38] * mat_B[216] +
//             mat_A[39] * mat_B[248] +
//             mat_A[40] * mat_B[280] +
//             mat_A[41] * mat_B[312] +
//             mat_A[42] * mat_B[344] +
//             mat_A[43] * mat_B[376] +
//             mat_A[44] * mat_B[408] +
//             mat_A[45] * mat_B[440] +
//             mat_A[46] * mat_B[472] +
//             mat_A[47] * mat_B[504] +
//             mat_A[48] * mat_B[536] +
//             mat_A[49] * mat_B[568] +
//             mat_A[50] * mat_B[600] +
//             mat_A[51] * mat_B[632] +
//             mat_A[52] * mat_B[664] +
//             mat_A[53] * mat_B[696] +
//             mat_A[54] * mat_B[728] +
//             mat_A[55] * mat_B[760] +
//             mat_A[56] * mat_B[792] +
//             mat_A[57] * mat_B[824] +
//             mat_A[58] * mat_B[856] +
//             mat_A[59] * mat_B[888] +
//             mat_A[60] * mat_B[920] +
//             mat_A[61] * mat_B[952] +
//             mat_A[62] * mat_B[984] +
//             mat_A[63] * mat_B[1016];
//  mat_C[57] <= 
//             mat_A[32] * mat_B[25] +
//             mat_A[33] * mat_B[57] +
//             mat_A[34] * mat_B[89] +
//             mat_A[35] * mat_B[121] +
//             mat_A[36] * mat_B[153] +
//             mat_A[37] * mat_B[185] +
//             mat_A[38] * mat_B[217] +
//             mat_A[39] * mat_B[249] +
//             mat_A[40] * mat_B[281] +
//             mat_A[41] * mat_B[313] +
//             mat_A[42] * mat_B[345] +
//             mat_A[43] * mat_B[377] +
//             mat_A[44] * mat_B[409] +
//             mat_A[45] * mat_B[441] +
//             mat_A[46] * mat_B[473] +
//             mat_A[47] * mat_B[505] +
//             mat_A[48] * mat_B[537] +
//             mat_A[49] * mat_B[569] +
//             mat_A[50] * mat_B[601] +
//             mat_A[51] * mat_B[633] +
//             mat_A[52] * mat_B[665] +
//             mat_A[53] * mat_B[697] +
//             mat_A[54] * mat_B[729] +
//             mat_A[55] * mat_B[761] +
//             mat_A[56] * mat_B[793] +
//             mat_A[57] * mat_B[825] +
//             mat_A[58] * mat_B[857] +
//             mat_A[59] * mat_B[889] +
//             mat_A[60] * mat_B[921] +
//             mat_A[61] * mat_B[953] +
//             mat_A[62] * mat_B[985] +
//             mat_A[63] * mat_B[1017];
//  mat_C[58] <= 
//             mat_A[32] * mat_B[26] +
//             mat_A[33] * mat_B[58] +
//             mat_A[34] * mat_B[90] +
//             mat_A[35] * mat_B[122] +
//             mat_A[36] * mat_B[154] +
//             mat_A[37] * mat_B[186] +
//             mat_A[38] * mat_B[218] +
//             mat_A[39] * mat_B[250] +
//             mat_A[40] * mat_B[282] +
//             mat_A[41] * mat_B[314] +
//             mat_A[42] * mat_B[346] +
//             mat_A[43] * mat_B[378] +
//             mat_A[44] * mat_B[410] +
//             mat_A[45] * mat_B[442] +
//             mat_A[46] * mat_B[474] +
//             mat_A[47] * mat_B[506] +
//             mat_A[48] * mat_B[538] +
//             mat_A[49] * mat_B[570] +
//             mat_A[50] * mat_B[602] +
//             mat_A[51] * mat_B[634] +
//             mat_A[52] * mat_B[666] +
//             mat_A[53] * mat_B[698] +
//             mat_A[54] * mat_B[730] +
//             mat_A[55] * mat_B[762] +
//             mat_A[56] * mat_B[794] +
//             mat_A[57] * mat_B[826] +
//             mat_A[58] * mat_B[858] +
//             mat_A[59] * mat_B[890] +
//             mat_A[60] * mat_B[922] +
//             mat_A[61] * mat_B[954] +
//             mat_A[62] * mat_B[986] +
//             mat_A[63] * mat_B[1018];
//  mat_C[59] <= 
//             mat_A[32] * mat_B[27] +
//             mat_A[33] * mat_B[59] +
//             mat_A[34] * mat_B[91] +
//             mat_A[35] * mat_B[123] +
//             mat_A[36] * mat_B[155] +
//             mat_A[37] * mat_B[187] +
//             mat_A[38] * mat_B[219] +
//             mat_A[39] * mat_B[251] +
//             mat_A[40] * mat_B[283] +
//             mat_A[41] * mat_B[315] +
//             mat_A[42] * mat_B[347] +
//             mat_A[43] * mat_B[379] +
//             mat_A[44] * mat_B[411] +
//             mat_A[45] * mat_B[443] +
//             mat_A[46] * mat_B[475] +
//             mat_A[47] * mat_B[507] +
//             mat_A[48] * mat_B[539] +
//             mat_A[49] * mat_B[571] +
//             mat_A[50] * mat_B[603] +
//             mat_A[51] * mat_B[635] +
//             mat_A[52] * mat_B[667] +
//             mat_A[53] * mat_B[699] +
//             mat_A[54] * mat_B[731] +
//             mat_A[55] * mat_B[763] +
//             mat_A[56] * mat_B[795] +
//             mat_A[57] * mat_B[827] +
//             mat_A[58] * mat_B[859] +
//             mat_A[59] * mat_B[891] +
//             mat_A[60] * mat_B[923] +
//             mat_A[61] * mat_B[955] +
//             mat_A[62] * mat_B[987] +
//             mat_A[63] * mat_B[1019];
//  mat_C[60] <= 
//             mat_A[32] * mat_B[28] +
//             mat_A[33] * mat_B[60] +
//             mat_A[34] * mat_B[92] +
//             mat_A[35] * mat_B[124] +
//             mat_A[36] * mat_B[156] +
//             mat_A[37] * mat_B[188] +
//             mat_A[38] * mat_B[220] +
//             mat_A[39] * mat_B[252] +
//             mat_A[40] * mat_B[284] +
//             mat_A[41] * mat_B[316] +
//             mat_A[42] * mat_B[348] +
//             mat_A[43] * mat_B[380] +
//             mat_A[44] * mat_B[412] +
//             mat_A[45] * mat_B[444] +
//             mat_A[46] * mat_B[476] +
//             mat_A[47] * mat_B[508] +
//             mat_A[48] * mat_B[540] +
//             mat_A[49] * mat_B[572] +
//             mat_A[50] * mat_B[604] +
//             mat_A[51] * mat_B[636] +
//             mat_A[52] * mat_B[668] +
//             mat_A[53] * mat_B[700] +
//             mat_A[54] * mat_B[732] +
//             mat_A[55] * mat_B[764] +
//             mat_A[56] * mat_B[796] +
//             mat_A[57] * mat_B[828] +
//             mat_A[58] * mat_B[860] +
//             mat_A[59] * mat_B[892] +
//             mat_A[60] * mat_B[924] +
//             mat_A[61] * mat_B[956] +
//             mat_A[62] * mat_B[988] +
//             mat_A[63] * mat_B[1020];
//  mat_C[61] <= 
//             mat_A[32] * mat_B[29] +
//             mat_A[33] * mat_B[61] +
//             mat_A[34] * mat_B[93] +
//             mat_A[35] * mat_B[125] +
//             mat_A[36] * mat_B[157] +
//             mat_A[37] * mat_B[189] +
//             mat_A[38] * mat_B[221] +
//             mat_A[39] * mat_B[253] +
//             mat_A[40] * mat_B[285] +
//             mat_A[41] * mat_B[317] +
//             mat_A[42] * mat_B[349] +
//             mat_A[43] * mat_B[381] +
//             mat_A[44] * mat_B[413] +
//             mat_A[45] * mat_B[445] +
//             mat_A[46] * mat_B[477] +
//             mat_A[47] * mat_B[509] +
//             mat_A[48] * mat_B[541] +
//             mat_A[49] * mat_B[573] +
//             mat_A[50] * mat_B[605] +
//             mat_A[51] * mat_B[637] +
//             mat_A[52] * mat_B[669] +
//             mat_A[53] * mat_B[701] +
//             mat_A[54] * mat_B[733] +
//             mat_A[55] * mat_B[765] +
//             mat_A[56] * mat_B[797] +
//             mat_A[57] * mat_B[829] +
//             mat_A[58] * mat_B[861] +
//             mat_A[59] * mat_B[893] +
//             mat_A[60] * mat_B[925] +
//             mat_A[61] * mat_B[957] +
//             mat_A[62] * mat_B[989] +
//             mat_A[63] * mat_B[1021];
//  mat_C[62] <= 
//             mat_A[32] * mat_B[30] +
//             mat_A[33] * mat_B[62] +
//             mat_A[34] * mat_B[94] +
//             mat_A[35] * mat_B[126] +
//             mat_A[36] * mat_B[158] +
//             mat_A[37] * mat_B[190] +
//             mat_A[38] * mat_B[222] +
//             mat_A[39] * mat_B[254] +
//             mat_A[40] * mat_B[286] +
//             mat_A[41] * mat_B[318] +
//             mat_A[42] * mat_B[350] +
//             mat_A[43] * mat_B[382] +
//             mat_A[44] * mat_B[414] +
//             mat_A[45] * mat_B[446] +
//             mat_A[46] * mat_B[478] +
//             mat_A[47] * mat_B[510] +
//             mat_A[48] * mat_B[542] +
//             mat_A[49] * mat_B[574] +
//             mat_A[50] * mat_B[606] +
//             mat_A[51] * mat_B[638] +
//             mat_A[52] * mat_B[670] +
//             mat_A[53] * mat_B[702] +
//             mat_A[54] * mat_B[734] +
//             mat_A[55] * mat_B[766] +
//             mat_A[56] * mat_B[798] +
//             mat_A[57] * mat_B[830] +
//             mat_A[58] * mat_B[862] +
//             mat_A[59] * mat_B[894] +
//             mat_A[60] * mat_B[926] +
//             mat_A[61] * mat_B[958] +
//             mat_A[62] * mat_B[990] +
//             mat_A[63] * mat_B[1022];
//  mat_C[63] <= 
//             mat_A[32] * mat_B[31] +
//             mat_A[33] * mat_B[63] +
//             mat_A[34] * mat_B[95] +
//             mat_A[35] * mat_B[127] +
//             mat_A[36] * mat_B[159] +
//             mat_A[37] * mat_B[191] +
//             mat_A[38] * mat_B[223] +
//             mat_A[39] * mat_B[255] +
//             mat_A[40] * mat_B[287] +
//             mat_A[41] * mat_B[319] +
//             mat_A[42] * mat_B[351] +
//             mat_A[43] * mat_B[383] +
//             mat_A[44] * mat_B[415] +
//             mat_A[45] * mat_B[447] +
//             mat_A[46] * mat_B[479] +
//             mat_A[47] * mat_B[511] +
//             mat_A[48] * mat_B[543] +
//             mat_A[49] * mat_B[575] +
//             mat_A[50] * mat_B[607] +
//             mat_A[51] * mat_B[639] +
//             mat_A[52] * mat_B[671] +
//             mat_A[53] * mat_B[703] +
//             mat_A[54] * mat_B[735] +
//             mat_A[55] * mat_B[767] +
//             mat_A[56] * mat_B[799] +
//             mat_A[57] * mat_B[831] +
//             mat_A[58] * mat_B[863] +
//             mat_A[59] * mat_B[895] +
//             mat_A[60] * mat_B[927] +
//             mat_A[61] * mat_B[959] +
//             mat_A[62] * mat_B[991] +
//             mat_A[63] * mat_B[1023];
//  mat_C[64] <= 
//             mat_A[64] * mat_B[0] +
//             mat_A[65] * mat_B[32] +
//             mat_A[66] * mat_B[64] +
//             mat_A[67] * mat_B[96] +
//             mat_A[68] * mat_B[128] +
//             mat_A[69] * mat_B[160] +
//             mat_A[70] * mat_B[192] +
//             mat_A[71] * mat_B[224] +
//             mat_A[72] * mat_B[256] +
//             mat_A[73] * mat_B[288] +
//             mat_A[74] * mat_B[320] +
//             mat_A[75] * mat_B[352] +
//             mat_A[76] * mat_B[384] +
//             mat_A[77] * mat_B[416] +
//             mat_A[78] * mat_B[448] +
//             mat_A[79] * mat_B[480] +
//             mat_A[80] * mat_B[512] +
//             mat_A[81] * mat_B[544] +
//             mat_A[82] * mat_B[576] +
//             mat_A[83] * mat_B[608] +
//             mat_A[84] * mat_B[640] +
//             mat_A[85] * mat_B[672] +
//             mat_A[86] * mat_B[704] +
//             mat_A[87] * mat_B[736] +
//             mat_A[88] * mat_B[768] +
//             mat_A[89] * mat_B[800] +
//             mat_A[90] * mat_B[832] +
//             mat_A[91] * mat_B[864] +
//             mat_A[92] * mat_B[896] +
//             mat_A[93] * mat_B[928] +
//             mat_A[94] * mat_B[960] +
//             mat_A[95] * mat_B[992];
//  mat_C[65] <= 
//             mat_A[64] * mat_B[1] +
//             mat_A[65] * mat_B[33] +
//             mat_A[66] * mat_B[65] +
//             mat_A[67] * mat_B[97] +
//             mat_A[68] * mat_B[129] +
//             mat_A[69] * mat_B[161] +
//             mat_A[70] * mat_B[193] +
//             mat_A[71] * mat_B[225] +
//             mat_A[72] * mat_B[257] +
//             mat_A[73] * mat_B[289] +
//             mat_A[74] * mat_B[321] +
//             mat_A[75] * mat_B[353] +
//             mat_A[76] * mat_B[385] +
//             mat_A[77] * mat_B[417] +
//             mat_A[78] * mat_B[449] +
//             mat_A[79] * mat_B[481] +
//             mat_A[80] * mat_B[513] +
//             mat_A[81] * mat_B[545] +
//             mat_A[82] * mat_B[577] +
//             mat_A[83] * mat_B[609] +
//             mat_A[84] * mat_B[641] +
//             mat_A[85] * mat_B[673] +
//             mat_A[86] * mat_B[705] +
//             mat_A[87] * mat_B[737] +
//             mat_A[88] * mat_B[769] +
//             mat_A[89] * mat_B[801] +
//             mat_A[90] * mat_B[833] +
//             mat_A[91] * mat_B[865] +
//             mat_A[92] * mat_B[897] +
//             mat_A[93] * mat_B[929] +
//             mat_A[94] * mat_B[961] +
//             mat_A[95] * mat_B[993];
//  mat_C[66] <= 
//             mat_A[64] * mat_B[2] +
//             mat_A[65] * mat_B[34] +
//             mat_A[66] * mat_B[66] +
//             mat_A[67] * mat_B[98] +
//             mat_A[68] * mat_B[130] +
//             mat_A[69] * mat_B[162] +
//             mat_A[70] * mat_B[194] +
//             mat_A[71] * mat_B[226] +
//             mat_A[72] * mat_B[258] +
//             mat_A[73] * mat_B[290] +
//             mat_A[74] * mat_B[322] +
//             mat_A[75] * mat_B[354] +
//             mat_A[76] * mat_B[386] +
//             mat_A[77] * mat_B[418] +
//             mat_A[78] * mat_B[450] +
//             mat_A[79] * mat_B[482] +
//             mat_A[80] * mat_B[514] +
//             mat_A[81] * mat_B[546] +
//             mat_A[82] * mat_B[578] +
//             mat_A[83] * mat_B[610] +
//             mat_A[84] * mat_B[642] +
//             mat_A[85] * mat_B[674] +
//             mat_A[86] * mat_B[706] +
//             mat_A[87] * mat_B[738] +
//             mat_A[88] * mat_B[770] +
//             mat_A[89] * mat_B[802] +
//             mat_A[90] * mat_B[834] +
//             mat_A[91] * mat_B[866] +
//             mat_A[92] * mat_B[898] +
//             mat_A[93] * mat_B[930] +
//             mat_A[94] * mat_B[962] +
//             mat_A[95] * mat_B[994];
//  mat_C[67] <= 
//             mat_A[64] * mat_B[3] +
//             mat_A[65] * mat_B[35] +
//             mat_A[66] * mat_B[67] +
//             mat_A[67] * mat_B[99] +
//             mat_A[68] * mat_B[131] +
//             mat_A[69] * mat_B[163] +
//             mat_A[70] * mat_B[195] +
//             mat_A[71] * mat_B[227] +
//             mat_A[72] * mat_B[259] +
//             mat_A[73] * mat_B[291] +
//             mat_A[74] * mat_B[323] +
//             mat_A[75] * mat_B[355] +
//             mat_A[76] * mat_B[387] +
//             mat_A[77] * mat_B[419] +
//             mat_A[78] * mat_B[451] +
//             mat_A[79] * mat_B[483] +
//             mat_A[80] * mat_B[515] +
//             mat_A[81] * mat_B[547] +
//             mat_A[82] * mat_B[579] +
//             mat_A[83] * mat_B[611] +
//             mat_A[84] * mat_B[643] +
//             mat_A[85] * mat_B[675] +
//             mat_A[86] * mat_B[707] +
//             mat_A[87] * mat_B[739] +
//             mat_A[88] * mat_B[771] +
//             mat_A[89] * mat_B[803] +
//             mat_A[90] * mat_B[835] +
//             mat_A[91] * mat_B[867] +
//             mat_A[92] * mat_B[899] +
//             mat_A[93] * mat_B[931] +
//             mat_A[94] * mat_B[963] +
//             mat_A[95] * mat_B[995];
//  mat_C[68] <= 
//             mat_A[64] * mat_B[4] +
//             mat_A[65] * mat_B[36] +
//             mat_A[66] * mat_B[68] +
//             mat_A[67] * mat_B[100] +
//             mat_A[68] * mat_B[132] +
//             mat_A[69] * mat_B[164] +
//             mat_A[70] * mat_B[196] +
//             mat_A[71] * mat_B[228] +
//             mat_A[72] * mat_B[260] +
//             mat_A[73] * mat_B[292] +
//             mat_A[74] * mat_B[324] +
//             mat_A[75] * mat_B[356] +
//             mat_A[76] * mat_B[388] +
//             mat_A[77] * mat_B[420] +
//             mat_A[78] * mat_B[452] +
//             mat_A[79] * mat_B[484] +
//             mat_A[80] * mat_B[516] +
//             mat_A[81] * mat_B[548] +
//             mat_A[82] * mat_B[580] +
//             mat_A[83] * mat_B[612] +
//             mat_A[84] * mat_B[644] +
//             mat_A[85] * mat_B[676] +
//             mat_A[86] * mat_B[708] +
//             mat_A[87] * mat_B[740] +
//             mat_A[88] * mat_B[772] +
//             mat_A[89] * mat_B[804] +
//             mat_A[90] * mat_B[836] +
//             mat_A[91] * mat_B[868] +
//             mat_A[92] * mat_B[900] +
//             mat_A[93] * mat_B[932] +
//             mat_A[94] * mat_B[964] +
//             mat_A[95] * mat_B[996];
//  mat_C[69] <= 
//             mat_A[64] * mat_B[5] +
//             mat_A[65] * mat_B[37] +
//             mat_A[66] * mat_B[69] +
//             mat_A[67] * mat_B[101] +
//             mat_A[68] * mat_B[133] +
//             mat_A[69] * mat_B[165] +
//             mat_A[70] * mat_B[197] +
//             mat_A[71] * mat_B[229] +
//             mat_A[72] * mat_B[261] +
//             mat_A[73] * mat_B[293] +
//             mat_A[74] * mat_B[325] +
//             mat_A[75] * mat_B[357] +
//             mat_A[76] * mat_B[389] +
//             mat_A[77] * mat_B[421] +
//             mat_A[78] * mat_B[453] +
//             mat_A[79] * mat_B[485] +
//             mat_A[80] * mat_B[517] +
//             mat_A[81] * mat_B[549] +
//             mat_A[82] * mat_B[581] +
//             mat_A[83] * mat_B[613] +
//             mat_A[84] * mat_B[645] +
//             mat_A[85] * mat_B[677] +
//             mat_A[86] * mat_B[709] +
//             mat_A[87] * mat_B[741] +
//             mat_A[88] * mat_B[773] +
//             mat_A[89] * mat_B[805] +
//             mat_A[90] * mat_B[837] +
//             mat_A[91] * mat_B[869] +
//             mat_A[92] * mat_B[901] +
//             mat_A[93] * mat_B[933] +
//             mat_A[94] * mat_B[965] +
//             mat_A[95] * mat_B[997];
//  mat_C[70] <= 
//             mat_A[64] * mat_B[6] +
//             mat_A[65] * mat_B[38] +
//             mat_A[66] * mat_B[70] +
//             mat_A[67] * mat_B[102] +
//             mat_A[68] * mat_B[134] +
//             mat_A[69] * mat_B[166] +
//             mat_A[70] * mat_B[198] +
//             mat_A[71] * mat_B[230] +
//             mat_A[72] * mat_B[262] +
//             mat_A[73] * mat_B[294] +
//             mat_A[74] * mat_B[326] +
//             mat_A[75] * mat_B[358] +
//             mat_A[76] * mat_B[390] +
//             mat_A[77] * mat_B[422] +
//             mat_A[78] * mat_B[454] +
//             mat_A[79] * mat_B[486] +
//             mat_A[80] * mat_B[518] +
//             mat_A[81] * mat_B[550] +
//             mat_A[82] * mat_B[582] +
//             mat_A[83] * mat_B[614] +
//             mat_A[84] * mat_B[646] +
//             mat_A[85] * mat_B[678] +
//             mat_A[86] * mat_B[710] +
//             mat_A[87] * mat_B[742] +
//             mat_A[88] * mat_B[774] +
//             mat_A[89] * mat_B[806] +
//             mat_A[90] * mat_B[838] +
//             mat_A[91] * mat_B[870] +
//             mat_A[92] * mat_B[902] +
//             mat_A[93] * mat_B[934] +
//             mat_A[94] * mat_B[966] +
//             mat_A[95] * mat_B[998];
//  mat_C[71] <= 
//             mat_A[64] * mat_B[7] +
//             mat_A[65] * mat_B[39] +
//             mat_A[66] * mat_B[71] +
//             mat_A[67] * mat_B[103] +
//             mat_A[68] * mat_B[135] +
//             mat_A[69] * mat_B[167] +
//             mat_A[70] * mat_B[199] +
//             mat_A[71] * mat_B[231] +
//             mat_A[72] * mat_B[263] +
//             mat_A[73] * mat_B[295] +
//             mat_A[74] * mat_B[327] +
//             mat_A[75] * mat_B[359] +
//             mat_A[76] * mat_B[391] +
//             mat_A[77] * mat_B[423] +
//             mat_A[78] * mat_B[455] +
//             mat_A[79] * mat_B[487] +
//             mat_A[80] * mat_B[519] +
//             mat_A[81] * mat_B[551] +
//             mat_A[82] * mat_B[583] +
//             mat_A[83] * mat_B[615] +
//             mat_A[84] * mat_B[647] +
//             mat_A[85] * mat_B[679] +
//             mat_A[86] * mat_B[711] +
//             mat_A[87] * mat_B[743] +
//             mat_A[88] * mat_B[775] +
//             mat_A[89] * mat_B[807] +
//             mat_A[90] * mat_B[839] +
//             mat_A[91] * mat_B[871] +
//             mat_A[92] * mat_B[903] +
//             mat_A[93] * mat_B[935] +
//             mat_A[94] * mat_B[967] +
//             mat_A[95] * mat_B[999];
//  mat_C[72] <= 
//             mat_A[64] * mat_B[8] +
//             mat_A[65] * mat_B[40] +
//             mat_A[66] * mat_B[72] +
//             mat_A[67] * mat_B[104] +
//             mat_A[68] * mat_B[136] +
//             mat_A[69] * mat_B[168] +
//             mat_A[70] * mat_B[200] +
//             mat_A[71] * mat_B[232] +
//             mat_A[72] * mat_B[264] +
//             mat_A[73] * mat_B[296] +
//             mat_A[74] * mat_B[328] +
//             mat_A[75] * mat_B[360] +
//             mat_A[76] * mat_B[392] +
//             mat_A[77] * mat_B[424] +
//             mat_A[78] * mat_B[456] +
//             mat_A[79] * mat_B[488] +
//             mat_A[80] * mat_B[520] +
//             mat_A[81] * mat_B[552] +
//             mat_A[82] * mat_B[584] +
//             mat_A[83] * mat_B[616] +
//             mat_A[84] * mat_B[648] +
//             mat_A[85] * mat_B[680] +
//             mat_A[86] * mat_B[712] +
//             mat_A[87] * mat_B[744] +
//             mat_A[88] * mat_B[776] +
//             mat_A[89] * mat_B[808] +
//             mat_A[90] * mat_B[840] +
//             mat_A[91] * mat_B[872] +
//             mat_A[92] * mat_B[904] +
//             mat_A[93] * mat_B[936] +
//             mat_A[94] * mat_B[968] +
//             mat_A[95] * mat_B[1000];
//  mat_C[73] <= 
//             mat_A[64] * mat_B[9] +
//             mat_A[65] * mat_B[41] +
//             mat_A[66] * mat_B[73] +
//             mat_A[67] * mat_B[105] +
//             mat_A[68] * mat_B[137] +
//             mat_A[69] * mat_B[169] +
//             mat_A[70] * mat_B[201] +
//             mat_A[71] * mat_B[233] +
//             mat_A[72] * mat_B[265] +
//             mat_A[73] * mat_B[297] +
//             mat_A[74] * mat_B[329] +
//             mat_A[75] * mat_B[361] +
//             mat_A[76] * mat_B[393] +
//             mat_A[77] * mat_B[425] +
//             mat_A[78] * mat_B[457] +
//             mat_A[79] * mat_B[489] +
//             mat_A[80] * mat_B[521] +
//             mat_A[81] * mat_B[553] +
//             mat_A[82] * mat_B[585] +
//             mat_A[83] * mat_B[617] +
//             mat_A[84] * mat_B[649] +
//             mat_A[85] * mat_B[681] +
//             mat_A[86] * mat_B[713] +
//             mat_A[87] * mat_B[745] +
//             mat_A[88] * mat_B[777] +
//             mat_A[89] * mat_B[809] +
//             mat_A[90] * mat_B[841] +
//             mat_A[91] * mat_B[873] +
//             mat_A[92] * mat_B[905] +
//             mat_A[93] * mat_B[937] +
//             mat_A[94] * mat_B[969] +
//             mat_A[95] * mat_B[1001];
//  mat_C[74] <= 
//             mat_A[64] * mat_B[10] +
//             mat_A[65] * mat_B[42] +
//             mat_A[66] * mat_B[74] +
//             mat_A[67] * mat_B[106] +
//             mat_A[68] * mat_B[138] +
//             mat_A[69] * mat_B[170] +
//             mat_A[70] * mat_B[202] +
//             mat_A[71] * mat_B[234] +
//             mat_A[72] * mat_B[266] +
//             mat_A[73] * mat_B[298] +
//             mat_A[74] * mat_B[330] +
//             mat_A[75] * mat_B[362] +
//             mat_A[76] * mat_B[394] +
//             mat_A[77] * mat_B[426] +
//             mat_A[78] * mat_B[458] +
//             mat_A[79] * mat_B[490] +
//             mat_A[80] * mat_B[522] +
//             mat_A[81] * mat_B[554] +
//             mat_A[82] * mat_B[586] +
//             mat_A[83] * mat_B[618] +
//             mat_A[84] * mat_B[650] +
//             mat_A[85] * mat_B[682] +
//             mat_A[86] * mat_B[714] +
//             mat_A[87] * mat_B[746] +
//             mat_A[88] * mat_B[778] +
//             mat_A[89] * mat_B[810] +
//             mat_A[90] * mat_B[842] +
//             mat_A[91] * mat_B[874] +
//             mat_A[92] * mat_B[906] +
//             mat_A[93] * mat_B[938] +
//             mat_A[94] * mat_B[970] +
//             mat_A[95] * mat_B[1002];
//  mat_C[75] <= 
//             mat_A[64] * mat_B[11] +
//             mat_A[65] * mat_B[43] +
//             mat_A[66] * mat_B[75] +
//             mat_A[67] * mat_B[107] +
//             mat_A[68] * mat_B[139] +
//             mat_A[69] * mat_B[171] +
//             mat_A[70] * mat_B[203] +
//             mat_A[71] * mat_B[235] +
//             mat_A[72] * mat_B[267] +
//             mat_A[73] * mat_B[299] +
//             mat_A[74] * mat_B[331] +
//             mat_A[75] * mat_B[363] +
//             mat_A[76] * mat_B[395] +
//             mat_A[77] * mat_B[427] +
//             mat_A[78] * mat_B[459] +
//             mat_A[79] * mat_B[491] +
//             mat_A[80] * mat_B[523] +
//             mat_A[81] * mat_B[555] +
//             mat_A[82] * mat_B[587] +
//             mat_A[83] * mat_B[619] +
//             mat_A[84] * mat_B[651] +
//             mat_A[85] * mat_B[683] +
//             mat_A[86] * mat_B[715] +
//             mat_A[87] * mat_B[747] +
//             mat_A[88] * mat_B[779] +
//             mat_A[89] * mat_B[811] +
//             mat_A[90] * mat_B[843] +
//             mat_A[91] * mat_B[875] +
//             mat_A[92] * mat_B[907] +
//             mat_A[93] * mat_B[939] +
//             mat_A[94] * mat_B[971] +
//             mat_A[95] * mat_B[1003];
//  mat_C[76] <= 
//             mat_A[64] * mat_B[12] +
//             mat_A[65] * mat_B[44] +
//             mat_A[66] * mat_B[76] +
//             mat_A[67] * mat_B[108] +
//             mat_A[68] * mat_B[140] +
//             mat_A[69] * mat_B[172] +
//             mat_A[70] * mat_B[204] +
//             mat_A[71] * mat_B[236] +
//             mat_A[72] * mat_B[268] +
//             mat_A[73] * mat_B[300] +
//             mat_A[74] * mat_B[332] +
//             mat_A[75] * mat_B[364] +
//             mat_A[76] * mat_B[396] +
//             mat_A[77] * mat_B[428] +
//             mat_A[78] * mat_B[460] +
//             mat_A[79] * mat_B[492] +
//             mat_A[80] * mat_B[524] +
//             mat_A[81] * mat_B[556] +
//             mat_A[82] * mat_B[588] +
//             mat_A[83] * mat_B[620] +
//             mat_A[84] * mat_B[652] +
//             mat_A[85] * mat_B[684] +
//             mat_A[86] * mat_B[716] +
//             mat_A[87] * mat_B[748] +
//             mat_A[88] * mat_B[780] +
//             mat_A[89] * mat_B[812] +
//             mat_A[90] * mat_B[844] +
//             mat_A[91] * mat_B[876] +
//             mat_A[92] * mat_B[908] +
//             mat_A[93] * mat_B[940] +
//             mat_A[94] * mat_B[972] +
//             mat_A[95] * mat_B[1004];
//  mat_C[77] <= 
//             mat_A[64] * mat_B[13] +
//             mat_A[65] * mat_B[45] +
//             mat_A[66] * mat_B[77] +
//             mat_A[67] * mat_B[109] +
//             mat_A[68] * mat_B[141] +
//             mat_A[69] * mat_B[173] +
//             mat_A[70] * mat_B[205] +
//             mat_A[71] * mat_B[237] +
//             mat_A[72] * mat_B[269] +
//             mat_A[73] * mat_B[301] +
//             mat_A[74] * mat_B[333] +
//             mat_A[75] * mat_B[365] +
//             mat_A[76] * mat_B[397] +
//             mat_A[77] * mat_B[429] +
//             mat_A[78] * mat_B[461] +
//             mat_A[79] * mat_B[493] +
//             mat_A[80] * mat_B[525] +
//             mat_A[81] * mat_B[557] +
//             mat_A[82] * mat_B[589] +
//             mat_A[83] * mat_B[621] +
//             mat_A[84] * mat_B[653] +
//             mat_A[85] * mat_B[685] +
//             mat_A[86] * mat_B[717] +
//             mat_A[87] * mat_B[749] +
//             mat_A[88] * mat_B[781] +
//             mat_A[89] * mat_B[813] +
//             mat_A[90] * mat_B[845] +
//             mat_A[91] * mat_B[877] +
//             mat_A[92] * mat_B[909] +
//             mat_A[93] * mat_B[941] +
//             mat_A[94] * mat_B[973] +
//             mat_A[95] * mat_B[1005];
//  mat_C[78] <= 
//             mat_A[64] * mat_B[14] +
//             mat_A[65] * mat_B[46] +
//             mat_A[66] * mat_B[78] +
//             mat_A[67] * mat_B[110] +
//             mat_A[68] * mat_B[142] +
//             mat_A[69] * mat_B[174] +
//             mat_A[70] * mat_B[206] +
//             mat_A[71] * mat_B[238] +
//             mat_A[72] * mat_B[270] +
//             mat_A[73] * mat_B[302] +
//             mat_A[74] * mat_B[334] +
//             mat_A[75] * mat_B[366] +
//             mat_A[76] * mat_B[398] +
//             mat_A[77] * mat_B[430] +
//             mat_A[78] * mat_B[462] +
//             mat_A[79] * mat_B[494] +
//             mat_A[80] * mat_B[526] +
//             mat_A[81] * mat_B[558] +
//             mat_A[82] * mat_B[590] +
//             mat_A[83] * mat_B[622] +
//             mat_A[84] * mat_B[654] +
//             mat_A[85] * mat_B[686] +
//             mat_A[86] * mat_B[718] +
//             mat_A[87] * mat_B[750] +
//             mat_A[88] * mat_B[782] +
//             mat_A[89] * mat_B[814] +
//             mat_A[90] * mat_B[846] +
//             mat_A[91] * mat_B[878] +
//             mat_A[92] * mat_B[910] +
//             mat_A[93] * mat_B[942] +
//             mat_A[94] * mat_B[974] +
//             mat_A[95] * mat_B[1006];
//  mat_C[79] <= 
//             mat_A[64] * mat_B[15] +
//             mat_A[65] * mat_B[47] +
//             mat_A[66] * mat_B[79] +
//             mat_A[67] * mat_B[111] +
//             mat_A[68] * mat_B[143] +
//             mat_A[69] * mat_B[175] +
//             mat_A[70] * mat_B[207] +
//             mat_A[71] * mat_B[239] +
//             mat_A[72] * mat_B[271] +
//             mat_A[73] * mat_B[303] +
//             mat_A[74] * mat_B[335] +
//             mat_A[75] * mat_B[367] +
//             mat_A[76] * mat_B[399] +
//             mat_A[77] * mat_B[431] +
//             mat_A[78] * mat_B[463] +
//             mat_A[79] * mat_B[495] +
//             mat_A[80] * mat_B[527] +
//             mat_A[81] * mat_B[559] +
//             mat_A[82] * mat_B[591] +
//             mat_A[83] * mat_B[623] +
//             mat_A[84] * mat_B[655] +
//             mat_A[85] * mat_B[687] +
//             mat_A[86] * mat_B[719] +
//             mat_A[87] * mat_B[751] +
//             mat_A[88] * mat_B[783] +
//             mat_A[89] * mat_B[815] +
//             mat_A[90] * mat_B[847] +
//             mat_A[91] * mat_B[879] +
//             mat_A[92] * mat_B[911] +
//             mat_A[93] * mat_B[943] +
//             mat_A[94] * mat_B[975] +
//             mat_A[95] * mat_B[1007];
//  mat_C[80] <= 
//             mat_A[64] * mat_B[16] +
//             mat_A[65] * mat_B[48] +
//             mat_A[66] * mat_B[80] +
//             mat_A[67] * mat_B[112] +
//             mat_A[68] * mat_B[144] +
//             mat_A[69] * mat_B[176] +
//             mat_A[70] * mat_B[208] +
//             mat_A[71] * mat_B[240] +
//             mat_A[72] * mat_B[272] +
//             mat_A[73] * mat_B[304] +
//             mat_A[74] * mat_B[336] +
//             mat_A[75] * mat_B[368] +
//             mat_A[76] * mat_B[400] +
//             mat_A[77] * mat_B[432] +
//             mat_A[78] * mat_B[464] +
//             mat_A[79] * mat_B[496] +
//             mat_A[80] * mat_B[528] +
//             mat_A[81] * mat_B[560] +
//             mat_A[82] * mat_B[592] +
//             mat_A[83] * mat_B[624] +
//             mat_A[84] * mat_B[656] +
//             mat_A[85] * mat_B[688] +
//             mat_A[86] * mat_B[720] +
//             mat_A[87] * mat_B[752] +
//             mat_A[88] * mat_B[784] +
//             mat_A[89] * mat_B[816] +
//             mat_A[90] * mat_B[848] +
//             mat_A[91] * mat_B[880] +
//             mat_A[92] * mat_B[912] +
//             mat_A[93] * mat_B[944] +
//             mat_A[94] * mat_B[976] +
//             mat_A[95] * mat_B[1008];
//  mat_C[81] <= 
//             mat_A[64] * mat_B[17] +
//             mat_A[65] * mat_B[49] +
//             mat_A[66] * mat_B[81] +
//             mat_A[67] * mat_B[113] +
//             mat_A[68] * mat_B[145] +
//             mat_A[69] * mat_B[177] +
//             mat_A[70] * mat_B[209] +
//             mat_A[71] * mat_B[241] +
//             mat_A[72] * mat_B[273] +
//             mat_A[73] * mat_B[305] +
//             mat_A[74] * mat_B[337] +
//             mat_A[75] * mat_B[369] +
//             mat_A[76] * mat_B[401] +
//             mat_A[77] * mat_B[433] +
//             mat_A[78] * mat_B[465] +
//             mat_A[79] * mat_B[497] +
//             mat_A[80] * mat_B[529] +
//             mat_A[81] * mat_B[561] +
//             mat_A[82] * mat_B[593] +
//             mat_A[83] * mat_B[625] +
//             mat_A[84] * mat_B[657] +
//             mat_A[85] * mat_B[689] +
//             mat_A[86] * mat_B[721] +
//             mat_A[87] * mat_B[753] +
//             mat_A[88] * mat_B[785] +
//             mat_A[89] * mat_B[817] +
//             mat_A[90] * mat_B[849] +
//             mat_A[91] * mat_B[881] +
//             mat_A[92] * mat_B[913] +
//             mat_A[93] * mat_B[945] +
//             mat_A[94] * mat_B[977] +
//             mat_A[95] * mat_B[1009];
//  mat_C[82] <= 
//             mat_A[64] * mat_B[18] +
//             mat_A[65] * mat_B[50] +
//             mat_A[66] * mat_B[82] +
//             mat_A[67] * mat_B[114] +
//             mat_A[68] * mat_B[146] +
//             mat_A[69] * mat_B[178] +
//             mat_A[70] * mat_B[210] +
//             mat_A[71] * mat_B[242] +
//             mat_A[72] * mat_B[274] +
//             mat_A[73] * mat_B[306] +
//             mat_A[74] * mat_B[338] +
//             mat_A[75] * mat_B[370] +
//             mat_A[76] * mat_B[402] +
//             mat_A[77] * mat_B[434] +
//             mat_A[78] * mat_B[466] +
//             mat_A[79] * mat_B[498] +
//             mat_A[80] * mat_B[530] +
//             mat_A[81] * mat_B[562] +
//             mat_A[82] * mat_B[594] +
//             mat_A[83] * mat_B[626] +
//             mat_A[84] * mat_B[658] +
//             mat_A[85] * mat_B[690] +
//             mat_A[86] * mat_B[722] +
//             mat_A[87] * mat_B[754] +
//             mat_A[88] * mat_B[786] +
//             mat_A[89] * mat_B[818] +
//             mat_A[90] * mat_B[850] +
//             mat_A[91] * mat_B[882] +
//             mat_A[92] * mat_B[914] +
//             mat_A[93] * mat_B[946] +
//             mat_A[94] * mat_B[978] +
//             mat_A[95] * mat_B[1010];
//  mat_C[83] <= 
//             mat_A[64] * mat_B[19] +
//             mat_A[65] * mat_B[51] +
//             mat_A[66] * mat_B[83] +
//             mat_A[67] * mat_B[115] +
//             mat_A[68] * mat_B[147] +
//             mat_A[69] * mat_B[179] +
//             mat_A[70] * mat_B[211] +
//             mat_A[71] * mat_B[243] +
//             mat_A[72] * mat_B[275] +
//             mat_A[73] * mat_B[307] +
//             mat_A[74] * mat_B[339] +
//             mat_A[75] * mat_B[371] +
//             mat_A[76] * mat_B[403] +
//             mat_A[77] * mat_B[435] +
//             mat_A[78] * mat_B[467] +
//             mat_A[79] * mat_B[499] +
//             mat_A[80] * mat_B[531] +
//             mat_A[81] * mat_B[563] +
//             mat_A[82] * mat_B[595] +
//             mat_A[83] * mat_B[627] +
//             mat_A[84] * mat_B[659] +
//             mat_A[85] * mat_B[691] +
//             mat_A[86] * mat_B[723] +
//             mat_A[87] * mat_B[755] +
//             mat_A[88] * mat_B[787] +
//             mat_A[89] * mat_B[819] +
//             mat_A[90] * mat_B[851] +
//             mat_A[91] * mat_B[883] +
//             mat_A[92] * mat_B[915] +
//             mat_A[93] * mat_B[947] +
//             mat_A[94] * mat_B[979] +
//             mat_A[95] * mat_B[1011];
//  mat_C[84] <= 
//             mat_A[64] * mat_B[20] +
//             mat_A[65] * mat_B[52] +
//             mat_A[66] * mat_B[84] +
//             mat_A[67] * mat_B[116] +
//             mat_A[68] * mat_B[148] +
//             mat_A[69] * mat_B[180] +
//             mat_A[70] * mat_B[212] +
//             mat_A[71] * mat_B[244] +
//             mat_A[72] * mat_B[276] +
//             mat_A[73] * mat_B[308] +
//             mat_A[74] * mat_B[340] +
//             mat_A[75] * mat_B[372] +
//             mat_A[76] * mat_B[404] +
//             mat_A[77] * mat_B[436] +
//             mat_A[78] * mat_B[468] +
//             mat_A[79] * mat_B[500] +
//             mat_A[80] * mat_B[532] +
//             mat_A[81] * mat_B[564] +
//             mat_A[82] * mat_B[596] +
//             mat_A[83] * mat_B[628] +
//             mat_A[84] * mat_B[660] +
//             mat_A[85] * mat_B[692] +
//             mat_A[86] * mat_B[724] +
//             mat_A[87] * mat_B[756] +
//             mat_A[88] * mat_B[788] +
//             mat_A[89] * mat_B[820] +
//             mat_A[90] * mat_B[852] +
//             mat_A[91] * mat_B[884] +
//             mat_A[92] * mat_B[916] +
//             mat_A[93] * mat_B[948] +
//             mat_A[94] * mat_B[980] +
//             mat_A[95] * mat_B[1012];
//  mat_C[85] <= 
//             mat_A[64] * mat_B[21] +
//             mat_A[65] * mat_B[53] +
//             mat_A[66] * mat_B[85] +
//             mat_A[67] * mat_B[117] +
//             mat_A[68] * mat_B[149] +
//             mat_A[69] * mat_B[181] +
//             mat_A[70] * mat_B[213] +
//             mat_A[71] * mat_B[245] +
//             mat_A[72] * mat_B[277] +
//             mat_A[73] * mat_B[309] +
//             mat_A[74] * mat_B[341] +
//             mat_A[75] * mat_B[373] +
//             mat_A[76] * mat_B[405] +
//             mat_A[77] * mat_B[437] +
//             mat_A[78] * mat_B[469] +
//             mat_A[79] * mat_B[501] +
//             mat_A[80] * mat_B[533] +
//             mat_A[81] * mat_B[565] +
//             mat_A[82] * mat_B[597] +
//             mat_A[83] * mat_B[629] +
//             mat_A[84] * mat_B[661] +
//             mat_A[85] * mat_B[693] +
//             mat_A[86] * mat_B[725] +
//             mat_A[87] * mat_B[757] +
//             mat_A[88] * mat_B[789] +
//             mat_A[89] * mat_B[821] +
//             mat_A[90] * mat_B[853] +
//             mat_A[91] * mat_B[885] +
//             mat_A[92] * mat_B[917] +
//             mat_A[93] * mat_B[949] +
//             mat_A[94] * mat_B[981] +
//             mat_A[95] * mat_B[1013];
//  mat_C[86] <= 
//             mat_A[64] * mat_B[22] +
//             mat_A[65] * mat_B[54] +
//             mat_A[66] * mat_B[86] +
//             mat_A[67] * mat_B[118] +
//             mat_A[68] * mat_B[150] +
//             mat_A[69] * mat_B[182] +
//             mat_A[70] * mat_B[214] +
//             mat_A[71] * mat_B[246] +
//             mat_A[72] * mat_B[278] +
//             mat_A[73] * mat_B[310] +
//             mat_A[74] * mat_B[342] +
//             mat_A[75] * mat_B[374] +
//             mat_A[76] * mat_B[406] +
//             mat_A[77] * mat_B[438] +
//             mat_A[78] * mat_B[470] +
//             mat_A[79] * mat_B[502] +
//             mat_A[80] * mat_B[534] +
//             mat_A[81] * mat_B[566] +
//             mat_A[82] * mat_B[598] +
//             mat_A[83] * mat_B[630] +
//             mat_A[84] * mat_B[662] +
//             mat_A[85] * mat_B[694] +
//             mat_A[86] * mat_B[726] +
//             mat_A[87] * mat_B[758] +
//             mat_A[88] * mat_B[790] +
//             mat_A[89] * mat_B[822] +
//             mat_A[90] * mat_B[854] +
//             mat_A[91] * mat_B[886] +
//             mat_A[92] * mat_B[918] +
//             mat_A[93] * mat_B[950] +
//             mat_A[94] * mat_B[982] +
//             mat_A[95] * mat_B[1014];
//  mat_C[87] <= 
//             mat_A[64] * mat_B[23] +
//             mat_A[65] * mat_B[55] +
//             mat_A[66] * mat_B[87] +
//             mat_A[67] * mat_B[119] +
//             mat_A[68] * mat_B[151] +
//             mat_A[69] * mat_B[183] +
//             mat_A[70] * mat_B[215] +
//             mat_A[71] * mat_B[247] +
//             mat_A[72] * mat_B[279] +
//             mat_A[73] * mat_B[311] +
//             mat_A[74] * mat_B[343] +
//             mat_A[75] * mat_B[375] +
//             mat_A[76] * mat_B[407] +
//             mat_A[77] * mat_B[439] +
//             mat_A[78] * mat_B[471] +
//             mat_A[79] * mat_B[503] +
//             mat_A[80] * mat_B[535] +
//             mat_A[81] * mat_B[567] +
//             mat_A[82] * mat_B[599] +
//             mat_A[83] * mat_B[631] +
//             mat_A[84] * mat_B[663] +
//             mat_A[85] * mat_B[695] +
//             mat_A[86] * mat_B[727] +
//             mat_A[87] * mat_B[759] +
//             mat_A[88] * mat_B[791] +
//             mat_A[89] * mat_B[823] +
//             mat_A[90] * mat_B[855] +
//             mat_A[91] * mat_B[887] +
//             mat_A[92] * mat_B[919] +
//             mat_A[93] * mat_B[951] +
//             mat_A[94] * mat_B[983] +
//             mat_A[95] * mat_B[1015];
//  mat_C[88] <= 
//             mat_A[64] * mat_B[24] +
//             mat_A[65] * mat_B[56] +
//             mat_A[66] * mat_B[88] +
//             mat_A[67] * mat_B[120] +
//             mat_A[68] * mat_B[152] +
//             mat_A[69] * mat_B[184] +
//             mat_A[70] * mat_B[216] +
//             mat_A[71] * mat_B[248] +
//             mat_A[72] * mat_B[280] +
//             mat_A[73] * mat_B[312] +
//             mat_A[74] * mat_B[344] +
//             mat_A[75] * mat_B[376] +
//             mat_A[76] * mat_B[408] +
//             mat_A[77] * mat_B[440] +
//             mat_A[78] * mat_B[472] +
//             mat_A[79] * mat_B[504] +
//             mat_A[80] * mat_B[536] +
//             mat_A[81] * mat_B[568] +
//             mat_A[82] * mat_B[600] +
//             mat_A[83] * mat_B[632] +
//             mat_A[84] * mat_B[664] +
//             mat_A[85] * mat_B[696] +
//             mat_A[86] * mat_B[728] +
//             mat_A[87] * mat_B[760] +
//             mat_A[88] * mat_B[792] +
//             mat_A[89] * mat_B[824] +
//             mat_A[90] * mat_B[856] +
//             mat_A[91] * mat_B[888] +
//             mat_A[92] * mat_B[920] +
//             mat_A[93] * mat_B[952] +
//             mat_A[94] * mat_B[984] +
//             mat_A[95] * mat_B[1016];
//  mat_C[89] <= 
//             mat_A[64] * mat_B[25] +
//             mat_A[65] * mat_B[57] +
//             mat_A[66] * mat_B[89] +
//             mat_A[67] * mat_B[121] +
//             mat_A[68] * mat_B[153] +
//             mat_A[69] * mat_B[185] +
//             mat_A[70] * mat_B[217] +
//             mat_A[71] * mat_B[249] +
//             mat_A[72] * mat_B[281] +
//             mat_A[73] * mat_B[313] +
//             mat_A[74] * mat_B[345] +
//             mat_A[75] * mat_B[377] +
//             mat_A[76] * mat_B[409] +
//             mat_A[77] * mat_B[441] +
//             mat_A[78] * mat_B[473] +
//             mat_A[79] * mat_B[505] +
//             mat_A[80] * mat_B[537] +
//             mat_A[81] * mat_B[569] +
//             mat_A[82] * mat_B[601] +
//             mat_A[83] * mat_B[633] +
//             mat_A[84] * mat_B[665] +
//             mat_A[85] * mat_B[697] +
//             mat_A[86] * mat_B[729] +
//             mat_A[87] * mat_B[761] +
//             mat_A[88] * mat_B[793] +
//             mat_A[89] * mat_B[825] +
//             mat_A[90] * mat_B[857] +
//             mat_A[91] * mat_B[889] +
//             mat_A[92] * mat_B[921] +
//             mat_A[93] * mat_B[953] +
//             mat_A[94] * mat_B[985] +
//             mat_A[95] * mat_B[1017];
//  mat_C[90] <= 
//             mat_A[64] * mat_B[26] +
//             mat_A[65] * mat_B[58] +
//             mat_A[66] * mat_B[90] +
//             mat_A[67] * mat_B[122] +
//             mat_A[68] * mat_B[154] +
//             mat_A[69] * mat_B[186] +
//             mat_A[70] * mat_B[218] +
//             mat_A[71] * mat_B[250] +
//             mat_A[72] * mat_B[282] +
//             mat_A[73] * mat_B[314] +
//             mat_A[74] * mat_B[346] +
//             mat_A[75] * mat_B[378] +
//             mat_A[76] * mat_B[410] +
//             mat_A[77] * mat_B[442] +
//             mat_A[78] * mat_B[474] +
//             mat_A[79] * mat_B[506] +
//             mat_A[80] * mat_B[538] +
//             mat_A[81] * mat_B[570] +
//             mat_A[82] * mat_B[602] +
//             mat_A[83] * mat_B[634] +
//             mat_A[84] * mat_B[666] +
//             mat_A[85] * mat_B[698] +
//             mat_A[86] * mat_B[730] +
//             mat_A[87] * mat_B[762] +
//             mat_A[88] * mat_B[794] +
//             mat_A[89] * mat_B[826] +
//             mat_A[90] * mat_B[858] +
//             mat_A[91] * mat_B[890] +
//             mat_A[92] * mat_B[922] +
//             mat_A[93] * mat_B[954] +
//             mat_A[94] * mat_B[986] +
//             mat_A[95] * mat_B[1018];
//  mat_C[91] <= 
//             mat_A[64] * mat_B[27] +
//             mat_A[65] * mat_B[59] +
//             mat_A[66] * mat_B[91] +
//             mat_A[67] * mat_B[123] +
//             mat_A[68] * mat_B[155] +
//             mat_A[69] * mat_B[187] +
//             mat_A[70] * mat_B[219] +
//             mat_A[71] * mat_B[251] +
//             mat_A[72] * mat_B[283] +
//             mat_A[73] * mat_B[315] +
//             mat_A[74] * mat_B[347] +
//             mat_A[75] * mat_B[379] +
//             mat_A[76] * mat_B[411] +
//             mat_A[77] * mat_B[443] +
//             mat_A[78] * mat_B[475] +
//             mat_A[79] * mat_B[507] +
//             mat_A[80] * mat_B[539] +
//             mat_A[81] * mat_B[571] +
//             mat_A[82] * mat_B[603] +
//             mat_A[83] * mat_B[635] +
//             mat_A[84] * mat_B[667] +
//             mat_A[85] * mat_B[699] +
//             mat_A[86] * mat_B[731] +
//             mat_A[87] * mat_B[763] +
//             mat_A[88] * mat_B[795] +
//             mat_A[89] * mat_B[827] +
//             mat_A[90] * mat_B[859] +
//             mat_A[91] * mat_B[891] +
//             mat_A[92] * mat_B[923] +
//             mat_A[93] * mat_B[955] +
//             mat_A[94] * mat_B[987] +
//             mat_A[95] * mat_B[1019];
//  mat_C[92] <= 
//             mat_A[64] * mat_B[28] +
//             mat_A[65] * mat_B[60] +
//             mat_A[66] * mat_B[92] +
//             mat_A[67] * mat_B[124] +
//             mat_A[68] * mat_B[156] +
//             mat_A[69] * mat_B[188] +
//             mat_A[70] * mat_B[220] +
//             mat_A[71] * mat_B[252] +
//             mat_A[72] * mat_B[284] +
//             mat_A[73] * mat_B[316] +
//             mat_A[74] * mat_B[348] +
//             mat_A[75] * mat_B[380] +
//             mat_A[76] * mat_B[412] +
//             mat_A[77] * mat_B[444] +
//             mat_A[78] * mat_B[476] +
//             mat_A[79] * mat_B[508] +
//             mat_A[80] * mat_B[540] +
//             mat_A[81] * mat_B[572] +
//             mat_A[82] * mat_B[604] +
//             mat_A[83] * mat_B[636] +
//             mat_A[84] * mat_B[668] +
//             mat_A[85] * mat_B[700] +
//             mat_A[86] * mat_B[732] +
//             mat_A[87] * mat_B[764] +
//             mat_A[88] * mat_B[796] +
//             mat_A[89] * mat_B[828] +
//             mat_A[90] * mat_B[860] +
//             mat_A[91] * mat_B[892] +
//             mat_A[92] * mat_B[924] +
//             mat_A[93] * mat_B[956] +
//             mat_A[94] * mat_B[988] +
//             mat_A[95] * mat_B[1020];
//  mat_C[93] <= 
//             mat_A[64] * mat_B[29] +
//             mat_A[65] * mat_B[61] +
//             mat_A[66] * mat_B[93] +
//             mat_A[67] * mat_B[125] +
//             mat_A[68] * mat_B[157] +
//             mat_A[69] * mat_B[189] +
//             mat_A[70] * mat_B[221] +
//             mat_A[71] * mat_B[253] +
//             mat_A[72] * mat_B[285] +
//             mat_A[73] * mat_B[317] +
//             mat_A[74] * mat_B[349] +
//             mat_A[75] * mat_B[381] +
//             mat_A[76] * mat_B[413] +
//             mat_A[77] * mat_B[445] +
//             mat_A[78] * mat_B[477] +
//             mat_A[79] * mat_B[509] +
//             mat_A[80] * mat_B[541] +
//             mat_A[81] * mat_B[573] +
//             mat_A[82] * mat_B[605] +
//             mat_A[83] * mat_B[637] +
//             mat_A[84] * mat_B[669] +
//             mat_A[85] * mat_B[701] +
//             mat_A[86] * mat_B[733] +
//             mat_A[87] * mat_B[765] +
//             mat_A[88] * mat_B[797] +
//             mat_A[89] * mat_B[829] +
//             mat_A[90] * mat_B[861] +
//             mat_A[91] * mat_B[893] +
//             mat_A[92] * mat_B[925] +
//             mat_A[93] * mat_B[957] +
//             mat_A[94] * mat_B[989] +
//             mat_A[95] * mat_B[1021];
//  mat_C[94] <= 
//             mat_A[64] * mat_B[30] +
//             mat_A[65] * mat_B[62] +
//             mat_A[66] * mat_B[94] +
//             mat_A[67] * mat_B[126] +
//             mat_A[68] * mat_B[158] +
//             mat_A[69] * mat_B[190] +
//             mat_A[70] * mat_B[222] +
//             mat_A[71] * mat_B[254] +
//             mat_A[72] * mat_B[286] +
//             mat_A[73] * mat_B[318] +
//             mat_A[74] * mat_B[350] +
//             mat_A[75] * mat_B[382] +
//             mat_A[76] * mat_B[414] +
//             mat_A[77] * mat_B[446] +
//             mat_A[78] * mat_B[478] +
//             mat_A[79] * mat_B[510] +
//             mat_A[80] * mat_B[542] +
//             mat_A[81] * mat_B[574] +
//             mat_A[82] * mat_B[606] +
//             mat_A[83] * mat_B[638] +
//             mat_A[84] * mat_B[670] +
//             mat_A[85] * mat_B[702] +
//             mat_A[86] * mat_B[734] +
//             mat_A[87] * mat_B[766] +
//             mat_A[88] * mat_B[798] +
//             mat_A[89] * mat_B[830] +
//             mat_A[90] * mat_B[862] +
//             mat_A[91] * mat_B[894] +
//             mat_A[92] * mat_B[926] +
//             mat_A[93] * mat_B[958] +
//             mat_A[94] * mat_B[990] +
//             mat_A[95] * mat_B[1022];
//  mat_C[95] <= 
//             mat_A[64] * mat_B[31] +
//             mat_A[65] * mat_B[63] +
//             mat_A[66] * mat_B[95] +
//             mat_A[67] * mat_B[127] +
//             mat_A[68] * mat_B[159] +
//             mat_A[69] * mat_B[191] +
//             mat_A[70] * mat_B[223] +
//             mat_A[71] * mat_B[255] +
//             mat_A[72] * mat_B[287] +
//             mat_A[73] * mat_B[319] +
//             mat_A[74] * mat_B[351] +
//             mat_A[75] * mat_B[383] +
//             mat_A[76] * mat_B[415] +
//             mat_A[77] * mat_B[447] +
//             mat_A[78] * mat_B[479] +
//             mat_A[79] * mat_B[511] +
//             mat_A[80] * mat_B[543] +
//             mat_A[81] * mat_B[575] +
//             mat_A[82] * mat_B[607] +
//             mat_A[83] * mat_B[639] +
//             mat_A[84] * mat_B[671] +
//             mat_A[85] * mat_B[703] +
//             mat_A[86] * mat_B[735] +
//             mat_A[87] * mat_B[767] +
//             mat_A[88] * mat_B[799] +
//             mat_A[89] * mat_B[831] +
//             mat_A[90] * mat_B[863] +
//             mat_A[91] * mat_B[895] +
//             mat_A[92] * mat_B[927] +
//             mat_A[93] * mat_B[959] +
//             mat_A[94] * mat_B[991] +
//             mat_A[95] * mat_B[1023];
//  mat_C[96] <= 
//             mat_A[96] * mat_B[0] +
//             mat_A[97] * mat_B[32] +
//             mat_A[98] * mat_B[64] +
//             mat_A[99] * mat_B[96] +
//             mat_A[100] * mat_B[128] +
//             mat_A[101] * mat_B[160] +
//             mat_A[102] * mat_B[192] +
//             mat_A[103] * mat_B[224] +
//             mat_A[104] * mat_B[256] +
//             mat_A[105] * mat_B[288] +
//             mat_A[106] * mat_B[320] +
//             mat_A[107] * mat_B[352] +
//             mat_A[108] * mat_B[384] +
//             mat_A[109] * mat_B[416] +
//             mat_A[110] * mat_B[448] +
//             mat_A[111] * mat_B[480] +
//             mat_A[112] * mat_B[512] +
//             mat_A[113] * mat_B[544] +
//             mat_A[114] * mat_B[576] +
//             mat_A[115] * mat_B[608] +
//             mat_A[116] * mat_B[640] +
//             mat_A[117] * mat_B[672] +
//             mat_A[118] * mat_B[704] +
//             mat_A[119] * mat_B[736] +
//             mat_A[120] * mat_B[768] +
//             mat_A[121] * mat_B[800] +
//             mat_A[122] * mat_B[832] +
//             mat_A[123] * mat_B[864] +
//             mat_A[124] * mat_B[896] +
//             mat_A[125] * mat_B[928] +
//             mat_A[126] * mat_B[960] +
//             mat_A[127] * mat_B[992];
//  mat_C[97] <= 
//             mat_A[96] * mat_B[1] +
//             mat_A[97] * mat_B[33] +
//             mat_A[98] * mat_B[65] +
//             mat_A[99] * mat_B[97] +
//             mat_A[100] * mat_B[129] +
//             mat_A[101] * mat_B[161] +
//             mat_A[102] * mat_B[193] +
//             mat_A[103] * mat_B[225] +
//             mat_A[104] * mat_B[257] +
//             mat_A[105] * mat_B[289] +
//             mat_A[106] * mat_B[321] +
//             mat_A[107] * mat_B[353] +
//             mat_A[108] * mat_B[385] +
//             mat_A[109] * mat_B[417] +
//             mat_A[110] * mat_B[449] +
//             mat_A[111] * mat_B[481] +
//             mat_A[112] * mat_B[513] +
//             mat_A[113] * mat_B[545] +
//             mat_A[114] * mat_B[577] +
//             mat_A[115] * mat_B[609] +
//             mat_A[116] * mat_B[641] +
//             mat_A[117] * mat_B[673] +
//             mat_A[118] * mat_B[705] +
//             mat_A[119] * mat_B[737] +
//             mat_A[120] * mat_B[769] +
//             mat_A[121] * mat_B[801] +
//             mat_A[122] * mat_B[833] +
//             mat_A[123] * mat_B[865] +
//             mat_A[124] * mat_B[897] +
//             mat_A[125] * mat_B[929] +
//             mat_A[126] * mat_B[961] +
//             mat_A[127] * mat_B[993];
//  mat_C[98] <= 
//             mat_A[96] * mat_B[2] +
//             mat_A[97] * mat_B[34] +
//             mat_A[98] * mat_B[66] +
//             mat_A[99] * mat_B[98] +
//             mat_A[100] * mat_B[130] +
//             mat_A[101] * mat_B[162] +
//             mat_A[102] * mat_B[194] +
//             mat_A[103] * mat_B[226] +
//             mat_A[104] * mat_B[258] +
//             mat_A[105] * mat_B[290] +
//             mat_A[106] * mat_B[322] +
//             mat_A[107] * mat_B[354] +
//             mat_A[108] * mat_B[386] +
//             mat_A[109] * mat_B[418] +
//             mat_A[110] * mat_B[450] +
//             mat_A[111] * mat_B[482] +
//             mat_A[112] * mat_B[514] +
//             mat_A[113] * mat_B[546] +
//             mat_A[114] * mat_B[578] +
//             mat_A[115] * mat_B[610] +
//             mat_A[116] * mat_B[642] +
//             mat_A[117] * mat_B[674] +
//             mat_A[118] * mat_B[706] +
//             mat_A[119] * mat_B[738] +
//             mat_A[120] * mat_B[770] +
//             mat_A[121] * mat_B[802] +
//             mat_A[122] * mat_B[834] +
//             mat_A[123] * mat_B[866] +
//             mat_A[124] * mat_B[898] +
//             mat_A[125] * mat_B[930] +
//             mat_A[126] * mat_B[962] +
//             mat_A[127] * mat_B[994];
//  mat_C[99] <= 
//             mat_A[96] * mat_B[3] +
//             mat_A[97] * mat_B[35] +
//             mat_A[98] * mat_B[67] +
//             mat_A[99] * mat_B[99] +
//             mat_A[100] * mat_B[131] +
//             mat_A[101] * mat_B[163] +
//             mat_A[102] * mat_B[195] +
//             mat_A[103] * mat_B[227] +
//             mat_A[104] * mat_B[259] +
//             mat_A[105] * mat_B[291] +
//             mat_A[106] * mat_B[323] +
//             mat_A[107] * mat_B[355] +
//             mat_A[108] * mat_B[387] +
//             mat_A[109] * mat_B[419] +
//             mat_A[110] * mat_B[451] +
//             mat_A[111] * mat_B[483] +
//             mat_A[112] * mat_B[515] +
//             mat_A[113] * mat_B[547] +
//             mat_A[114] * mat_B[579] +
//             mat_A[115] * mat_B[611] +
//             mat_A[116] * mat_B[643] +
//             mat_A[117] * mat_B[675] +
//             mat_A[118] * mat_B[707] +
//             mat_A[119] * mat_B[739] +
//             mat_A[120] * mat_B[771] +
//             mat_A[121] * mat_B[803] +
//             mat_A[122] * mat_B[835] +
//             mat_A[123] * mat_B[867] +
//             mat_A[124] * mat_B[899] +
//             mat_A[125] * mat_B[931] +
//             mat_A[126] * mat_B[963] +
//             mat_A[127] * mat_B[995];
//  mat_C[100] <= 
//             mat_A[96] * mat_B[4] +
//             mat_A[97] * mat_B[36] +
//             mat_A[98] * mat_B[68] +
//             mat_A[99] * mat_B[100] +
//             mat_A[100] * mat_B[132] +
//             mat_A[101] * mat_B[164] +
//             mat_A[102] * mat_B[196] +
//             mat_A[103] * mat_B[228] +
//             mat_A[104] * mat_B[260] +
//             mat_A[105] * mat_B[292] +
//             mat_A[106] * mat_B[324] +
//             mat_A[107] * mat_B[356] +
//             mat_A[108] * mat_B[388] +
//             mat_A[109] * mat_B[420] +
//             mat_A[110] * mat_B[452] +
//             mat_A[111] * mat_B[484] +
//             mat_A[112] * mat_B[516] +
//             mat_A[113] * mat_B[548] +
//             mat_A[114] * mat_B[580] +
//             mat_A[115] * mat_B[612] +
//             mat_A[116] * mat_B[644] +
//             mat_A[117] * mat_B[676] +
//             mat_A[118] * mat_B[708] +
//             mat_A[119] * mat_B[740] +
//             mat_A[120] * mat_B[772] +
//             mat_A[121] * mat_B[804] +
//             mat_A[122] * mat_B[836] +
//             mat_A[123] * mat_B[868] +
//             mat_A[124] * mat_B[900] +
//             mat_A[125] * mat_B[932] +
//             mat_A[126] * mat_B[964] +
//             mat_A[127] * mat_B[996];
//  mat_C[101] <= 
//             mat_A[96] * mat_B[5] +
//             mat_A[97] * mat_B[37] +
//             mat_A[98] * mat_B[69] +
//             mat_A[99] * mat_B[101] +
//             mat_A[100] * mat_B[133] +
//             mat_A[101] * mat_B[165] +
//             mat_A[102] * mat_B[197] +
//             mat_A[103] * mat_B[229] +
//             mat_A[104] * mat_B[261] +
//             mat_A[105] * mat_B[293] +
//             mat_A[106] * mat_B[325] +
//             mat_A[107] * mat_B[357] +
//             mat_A[108] * mat_B[389] +
//             mat_A[109] * mat_B[421] +
//             mat_A[110] * mat_B[453] +
//             mat_A[111] * mat_B[485] +
//             mat_A[112] * mat_B[517] +
//             mat_A[113] * mat_B[549] +
//             mat_A[114] * mat_B[581] +
//             mat_A[115] * mat_B[613] +
//             mat_A[116] * mat_B[645] +
//             mat_A[117] * mat_B[677] +
//             mat_A[118] * mat_B[709] +
//             mat_A[119] * mat_B[741] +
//             mat_A[120] * mat_B[773] +
//             mat_A[121] * mat_B[805] +
//             mat_A[122] * mat_B[837] +
//             mat_A[123] * mat_B[869] +
//             mat_A[124] * mat_B[901] +
//             mat_A[125] * mat_B[933] +
//             mat_A[126] * mat_B[965] +
//             mat_A[127] * mat_B[997];
//  mat_C[102] <= 
//             mat_A[96] * mat_B[6] +
//             mat_A[97] * mat_B[38] +
//             mat_A[98] * mat_B[70] +
//             mat_A[99] * mat_B[102] +
//             mat_A[100] * mat_B[134] +
//             mat_A[101] * mat_B[166] +
//             mat_A[102] * mat_B[198] +
//             mat_A[103] * mat_B[230] +
//             mat_A[104] * mat_B[262] +
//             mat_A[105] * mat_B[294] +
//             mat_A[106] * mat_B[326] +
//             mat_A[107] * mat_B[358] +
//             mat_A[108] * mat_B[390] +
//             mat_A[109] * mat_B[422] +
//             mat_A[110] * mat_B[454] +
//             mat_A[111] * mat_B[486] +
//             mat_A[112] * mat_B[518] +
//             mat_A[113] * mat_B[550] +
//             mat_A[114] * mat_B[582] +
//             mat_A[115] * mat_B[614] +
//             mat_A[116] * mat_B[646] +
//             mat_A[117] * mat_B[678] +
//             mat_A[118] * mat_B[710] +
//             mat_A[119] * mat_B[742] +
//             mat_A[120] * mat_B[774] +
//             mat_A[121] * mat_B[806] +
//             mat_A[122] * mat_B[838] +
//             mat_A[123] * mat_B[870] +
//             mat_A[124] * mat_B[902] +
//             mat_A[125] * mat_B[934] +
//             mat_A[126] * mat_B[966] +
//             mat_A[127] * mat_B[998];
//  mat_C[103] <= 
//             mat_A[96] * mat_B[7] +
//             mat_A[97] * mat_B[39] +
//             mat_A[98] * mat_B[71] +
//             mat_A[99] * mat_B[103] +
//             mat_A[100] * mat_B[135] +
//             mat_A[101] * mat_B[167] +
//             mat_A[102] * mat_B[199] +
//             mat_A[103] * mat_B[231] +
//             mat_A[104] * mat_B[263] +
//             mat_A[105] * mat_B[295] +
//             mat_A[106] * mat_B[327] +
//             mat_A[107] * mat_B[359] +
//             mat_A[108] * mat_B[391] +
//             mat_A[109] * mat_B[423] +
//             mat_A[110] * mat_B[455] +
//             mat_A[111] * mat_B[487] +
//             mat_A[112] * mat_B[519] +
//             mat_A[113] * mat_B[551] +
//             mat_A[114] * mat_B[583] +
//             mat_A[115] * mat_B[615] +
//             mat_A[116] * mat_B[647] +
//             mat_A[117] * mat_B[679] +
//             mat_A[118] * mat_B[711] +
//             mat_A[119] * mat_B[743] +
//             mat_A[120] * mat_B[775] +
//             mat_A[121] * mat_B[807] +
//             mat_A[122] * mat_B[839] +
//             mat_A[123] * mat_B[871] +
//             mat_A[124] * mat_B[903] +
//             mat_A[125] * mat_B[935] +
//             mat_A[126] * mat_B[967] +
//             mat_A[127] * mat_B[999];
//  mat_C[104] <= 
//             mat_A[96] * mat_B[8] +
//             mat_A[97] * mat_B[40] +
//             mat_A[98] * mat_B[72] +
//             mat_A[99] * mat_B[104] +
//             mat_A[100] * mat_B[136] +
//             mat_A[101] * mat_B[168] +
//             mat_A[102] * mat_B[200] +
//             mat_A[103] * mat_B[232] +
//             mat_A[104] * mat_B[264] +
//             mat_A[105] * mat_B[296] +
//             mat_A[106] * mat_B[328] +
//             mat_A[107] * mat_B[360] +
//             mat_A[108] * mat_B[392] +
//             mat_A[109] * mat_B[424] +
//             mat_A[110] * mat_B[456] +
//             mat_A[111] * mat_B[488] +
//             mat_A[112] * mat_B[520] +
//             mat_A[113] * mat_B[552] +
//             mat_A[114] * mat_B[584] +
//             mat_A[115] * mat_B[616] +
//             mat_A[116] * mat_B[648] +
//             mat_A[117] * mat_B[680] +
//             mat_A[118] * mat_B[712] +
//             mat_A[119] * mat_B[744] +
//             mat_A[120] * mat_B[776] +
//             mat_A[121] * mat_B[808] +
//             mat_A[122] * mat_B[840] +
//             mat_A[123] * mat_B[872] +
//             mat_A[124] * mat_B[904] +
//             mat_A[125] * mat_B[936] +
//             mat_A[126] * mat_B[968] +
//             mat_A[127] * mat_B[1000];
//  mat_C[105] <= 
//             mat_A[96] * mat_B[9] +
//             mat_A[97] * mat_B[41] +
//             mat_A[98] * mat_B[73] +
//             mat_A[99] * mat_B[105] +
//             mat_A[100] * mat_B[137] +
//             mat_A[101] * mat_B[169] +
//             mat_A[102] * mat_B[201] +
//             mat_A[103] * mat_B[233] +
//             mat_A[104] * mat_B[265] +
//             mat_A[105] * mat_B[297] +
//             mat_A[106] * mat_B[329] +
//             mat_A[107] * mat_B[361] +
//             mat_A[108] * mat_B[393] +
//             mat_A[109] * mat_B[425] +
//             mat_A[110] * mat_B[457] +
//             mat_A[111] * mat_B[489] +
//             mat_A[112] * mat_B[521] +
//             mat_A[113] * mat_B[553] +
//             mat_A[114] * mat_B[585] +
//             mat_A[115] * mat_B[617] +
//             mat_A[116] * mat_B[649] +
//             mat_A[117] * mat_B[681] +
//             mat_A[118] * mat_B[713] +
//             mat_A[119] * mat_B[745] +
//             mat_A[120] * mat_B[777] +
//             mat_A[121] * mat_B[809] +
//             mat_A[122] * mat_B[841] +
//             mat_A[123] * mat_B[873] +
//             mat_A[124] * mat_B[905] +
//             mat_A[125] * mat_B[937] +
//             mat_A[126] * mat_B[969] +
//             mat_A[127] * mat_B[1001];
//  mat_C[106] <= 
//             mat_A[96] * mat_B[10] +
//             mat_A[97] * mat_B[42] +
//             mat_A[98] * mat_B[74] +
//             mat_A[99] * mat_B[106] +
//             mat_A[100] * mat_B[138] +
//             mat_A[101] * mat_B[170] +
//             mat_A[102] * mat_B[202] +
//             mat_A[103] * mat_B[234] +
//             mat_A[104] * mat_B[266] +
//             mat_A[105] * mat_B[298] +
//             mat_A[106] * mat_B[330] +
//             mat_A[107] * mat_B[362] +
//             mat_A[108] * mat_B[394] +
//             mat_A[109] * mat_B[426] +
//             mat_A[110] * mat_B[458] +
//             mat_A[111] * mat_B[490] +
//             mat_A[112] * mat_B[522] +
//             mat_A[113] * mat_B[554] +
//             mat_A[114] * mat_B[586] +
//             mat_A[115] * mat_B[618] +
//             mat_A[116] * mat_B[650] +
//             mat_A[117] * mat_B[682] +
//             mat_A[118] * mat_B[714] +
//             mat_A[119] * mat_B[746] +
//             mat_A[120] * mat_B[778] +
//             mat_A[121] * mat_B[810] +
//             mat_A[122] * mat_B[842] +
//             mat_A[123] * mat_B[874] +
//             mat_A[124] * mat_B[906] +
//             mat_A[125] * mat_B[938] +
//             mat_A[126] * mat_B[970] +
//             mat_A[127] * mat_B[1002];
//  mat_C[107] <= 
//             mat_A[96] * mat_B[11] +
//             mat_A[97] * mat_B[43] +
//             mat_A[98] * mat_B[75] +
//             mat_A[99] * mat_B[107] +
//             mat_A[100] * mat_B[139] +
//             mat_A[101] * mat_B[171] +
//             mat_A[102] * mat_B[203] +
//             mat_A[103] * mat_B[235] +
//             mat_A[104] * mat_B[267] +
//             mat_A[105] * mat_B[299] +
//             mat_A[106] * mat_B[331] +
//             mat_A[107] * mat_B[363] +
//             mat_A[108] * mat_B[395] +
//             mat_A[109] * mat_B[427] +
//             mat_A[110] * mat_B[459] +
//             mat_A[111] * mat_B[491] +
//             mat_A[112] * mat_B[523] +
//             mat_A[113] * mat_B[555] +
//             mat_A[114] * mat_B[587] +
//             mat_A[115] * mat_B[619] +
//             mat_A[116] * mat_B[651] +
//             mat_A[117] * mat_B[683] +
//             mat_A[118] * mat_B[715] +
//             mat_A[119] * mat_B[747] +
//             mat_A[120] * mat_B[779] +
//             mat_A[121] * mat_B[811] +
//             mat_A[122] * mat_B[843] +
//             mat_A[123] * mat_B[875] +
//             mat_A[124] * mat_B[907] +
//             mat_A[125] * mat_B[939] +
//             mat_A[126] * mat_B[971] +
//             mat_A[127] * mat_B[1003];
//  mat_C[108] <= 
//             mat_A[96] * mat_B[12] +
//             mat_A[97] * mat_B[44] +
//             mat_A[98] * mat_B[76] +
//             mat_A[99] * mat_B[108] +
//             mat_A[100] * mat_B[140] +
//             mat_A[101] * mat_B[172] +
//             mat_A[102] * mat_B[204] +
//             mat_A[103] * mat_B[236] +
//             mat_A[104] * mat_B[268] +
//             mat_A[105] * mat_B[300] +
//             mat_A[106] * mat_B[332] +
//             mat_A[107] * mat_B[364] +
//             mat_A[108] * mat_B[396] +
//             mat_A[109] * mat_B[428] +
//             mat_A[110] * mat_B[460] +
//             mat_A[111] * mat_B[492] +
//             mat_A[112] * mat_B[524] +
//             mat_A[113] * mat_B[556] +
//             mat_A[114] * mat_B[588] +
//             mat_A[115] * mat_B[620] +
//             mat_A[116] * mat_B[652] +
//             mat_A[117] * mat_B[684] +
//             mat_A[118] * mat_B[716] +
//             mat_A[119] * mat_B[748] +
//             mat_A[120] * mat_B[780] +
//             mat_A[121] * mat_B[812] +
//             mat_A[122] * mat_B[844] +
//             mat_A[123] * mat_B[876] +
//             mat_A[124] * mat_B[908] +
//             mat_A[125] * mat_B[940] +
//             mat_A[126] * mat_B[972] +
//             mat_A[127] * mat_B[1004];
//  mat_C[109] <= 
//             mat_A[96] * mat_B[13] +
//             mat_A[97] * mat_B[45] +
//             mat_A[98] * mat_B[77] +
//             mat_A[99] * mat_B[109] +
//             mat_A[100] * mat_B[141] +
//             mat_A[101] * mat_B[173] +
//             mat_A[102] * mat_B[205] +
//             mat_A[103] * mat_B[237] +
//             mat_A[104] * mat_B[269] +
//             mat_A[105] * mat_B[301] +
//             mat_A[106] * mat_B[333] +
//             mat_A[107] * mat_B[365] +
//             mat_A[108] * mat_B[397] +
//             mat_A[109] * mat_B[429] +
//             mat_A[110] * mat_B[461] +
//             mat_A[111] * mat_B[493] +
//             mat_A[112] * mat_B[525] +
//             mat_A[113] * mat_B[557] +
//             mat_A[114] * mat_B[589] +
//             mat_A[115] * mat_B[621] +
//             mat_A[116] * mat_B[653] +
//             mat_A[117] * mat_B[685] +
//             mat_A[118] * mat_B[717] +
//             mat_A[119] * mat_B[749] +
//             mat_A[120] * mat_B[781] +
//             mat_A[121] * mat_B[813] +
//             mat_A[122] * mat_B[845] +
//             mat_A[123] * mat_B[877] +
//             mat_A[124] * mat_B[909] +
//             mat_A[125] * mat_B[941] +
//             mat_A[126] * mat_B[973] +
//             mat_A[127] * mat_B[1005];
//  mat_C[110] <= 
//             mat_A[96] * mat_B[14] +
//             mat_A[97] * mat_B[46] +
//             mat_A[98] * mat_B[78] +
//             mat_A[99] * mat_B[110] +
//             mat_A[100] * mat_B[142] +
//             mat_A[101] * mat_B[174] +
//             mat_A[102] * mat_B[206] +
//             mat_A[103] * mat_B[238] +
//             mat_A[104] * mat_B[270] +
//             mat_A[105] * mat_B[302] +
//             mat_A[106] * mat_B[334] +
//             mat_A[107] * mat_B[366] +
//             mat_A[108] * mat_B[398] +
//             mat_A[109] * mat_B[430] +
//             mat_A[110] * mat_B[462] +
//             mat_A[111] * mat_B[494] +
//             mat_A[112] * mat_B[526] +
//             mat_A[113] * mat_B[558] +
//             mat_A[114] * mat_B[590] +
//             mat_A[115] * mat_B[622] +
//             mat_A[116] * mat_B[654] +
//             mat_A[117] * mat_B[686] +
//             mat_A[118] * mat_B[718] +
//             mat_A[119] * mat_B[750] +
//             mat_A[120] * mat_B[782] +
//             mat_A[121] * mat_B[814] +
//             mat_A[122] * mat_B[846] +
//             mat_A[123] * mat_B[878] +
//             mat_A[124] * mat_B[910] +
//             mat_A[125] * mat_B[942] +
//             mat_A[126] * mat_B[974] +
//             mat_A[127] * mat_B[1006];
//  mat_C[111] <= 
//             mat_A[96] * mat_B[15] +
//             mat_A[97] * mat_B[47] +
//             mat_A[98] * mat_B[79] +
//             mat_A[99] * mat_B[111] +
//             mat_A[100] * mat_B[143] +
//             mat_A[101] * mat_B[175] +
//             mat_A[102] * mat_B[207] +
//             mat_A[103] * mat_B[239] +
//             mat_A[104] * mat_B[271] +
//             mat_A[105] * mat_B[303] +
//             mat_A[106] * mat_B[335] +
//             mat_A[107] * mat_B[367] +
//             mat_A[108] * mat_B[399] +
//             mat_A[109] * mat_B[431] +
//             mat_A[110] * mat_B[463] +
//             mat_A[111] * mat_B[495] +
//             mat_A[112] * mat_B[527] +
//             mat_A[113] * mat_B[559] +
//             mat_A[114] * mat_B[591] +
//             mat_A[115] * mat_B[623] +
//             mat_A[116] * mat_B[655] +
//             mat_A[117] * mat_B[687] +
//             mat_A[118] * mat_B[719] +
//             mat_A[119] * mat_B[751] +
//             mat_A[120] * mat_B[783] +
//             mat_A[121] * mat_B[815] +
//             mat_A[122] * mat_B[847] +
//             mat_A[123] * mat_B[879] +
//             mat_A[124] * mat_B[911] +
//             mat_A[125] * mat_B[943] +
//             mat_A[126] * mat_B[975] +
//             mat_A[127] * mat_B[1007];
//  mat_C[112] <= 
//             mat_A[96] * mat_B[16] +
//             mat_A[97] * mat_B[48] +
//             mat_A[98] * mat_B[80] +
//             mat_A[99] * mat_B[112] +
//             mat_A[100] * mat_B[144] +
//             mat_A[101] * mat_B[176] +
//             mat_A[102] * mat_B[208] +
//             mat_A[103] * mat_B[240] +
//             mat_A[104] * mat_B[272] +
//             mat_A[105] * mat_B[304] +
//             mat_A[106] * mat_B[336] +
//             mat_A[107] * mat_B[368] +
//             mat_A[108] * mat_B[400] +
//             mat_A[109] * mat_B[432] +
//             mat_A[110] * mat_B[464] +
//             mat_A[111] * mat_B[496] +
//             mat_A[112] * mat_B[528] +
//             mat_A[113] * mat_B[560] +
//             mat_A[114] * mat_B[592] +
//             mat_A[115] * mat_B[624] +
//             mat_A[116] * mat_B[656] +
//             mat_A[117] * mat_B[688] +
//             mat_A[118] * mat_B[720] +
//             mat_A[119] * mat_B[752] +
//             mat_A[120] * mat_B[784] +
//             mat_A[121] * mat_B[816] +
//             mat_A[122] * mat_B[848] +
//             mat_A[123] * mat_B[880] +
//             mat_A[124] * mat_B[912] +
//             mat_A[125] * mat_B[944] +
//             mat_A[126] * mat_B[976] +
//             mat_A[127] * mat_B[1008];
//  mat_C[113] <= 
//             mat_A[96] * mat_B[17] +
//             mat_A[97] * mat_B[49] +
//             mat_A[98] * mat_B[81] +
//             mat_A[99] * mat_B[113] +
//             mat_A[100] * mat_B[145] +
//             mat_A[101] * mat_B[177] +
//             mat_A[102] * mat_B[209] +
//             mat_A[103] * mat_B[241] +
//             mat_A[104] * mat_B[273] +
//             mat_A[105] * mat_B[305] +
//             mat_A[106] * mat_B[337] +
//             mat_A[107] * mat_B[369] +
//             mat_A[108] * mat_B[401] +
//             mat_A[109] * mat_B[433] +
//             mat_A[110] * mat_B[465] +
//             mat_A[111] * mat_B[497] +
//             mat_A[112] * mat_B[529] +
//             mat_A[113] * mat_B[561] +
//             mat_A[114] * mat_B[593] +
//             mat_A[115] * mat_B[625] +
//             mat_A[116] * mat_B[657] +
//             mat_A[117] * mat_B[689] +
//             mat_A[118] * mat_B[721] +
//             mat_A[119] * mat_B[753] +
//             mat_A[120] * mat_B[785] +
//             mat_A[121] * mat_B[817] +
//             mat_A[122] * mat_B[849] +
//             mat_A[123] * mat_B[881] +
//             mat_A[124] * mat_B[913] +
//             mat_A[125] * mat_B[945] +
//             mat_A[126] * mat_B[977] +
//             mat_A[127] * mat_B[1009];
//  mat_C[114] <= 
//             mat_A[96] * mat_B[18] +
//             mat_A[97] * mat_B[50] +
//             mat_A[98] * mat_B[82] +
//             mat_A[99] * mat_B[114] +
//             mat_A[100] * mat_B[146] +
//             mat_A[101] * mat_B[178] +
//             mat_A[102] * mat_B[210] +
//             mat_A[103] * mat_B[242] +
//             mat_A[104] * mat_B[274] +
//             mat_A[105] * mat_B[306] +
//             mat_A[106] * mat_B[338] +
//             mat_A[107] * mat_B[370] +
//             mat_A[108] * mat_B[402] +
//             mat_A[109] * mat_B[434] +
//             mat_A[110] * mat_B[466] +
//             mat_A[111] * mat_B[498] +
//             mat_A[112] * mat_B[530] +
//             mat_A[113] * mat_B[562] +
//             mat_A[114] * mat_B[594] +
//             mat_A[115] * mat_B[626] +
//             mat_A[116] * mat_B[658] +
//             mat_A[117] * mat_B[690] +
//             mat_A[118] * mat_B[722] +
//             mat_A[119] * mat_B[754] +
//             mat_A[120] * mat_B[786] +
//             mat_A[121] * mat_B[818] +
//             mat_A[122] * mat_B[850] +
//             mat_A[123] * mat_B[882] +
//             mat_A[124] * mat_B[914] +
//             mat_A[125] * mat_B[946] +
//             mat_A[126] * mat_B[978] +
//             mat_A[127] * mat_B[1010];
//  mat_C[115] <= 
//             mat_A[96] * mat_B[19] +
//             mat_A[97] * mat_B[51] +
//             mat_A[98] * mat_B[83] +
//             mat_A[99] * mat_B[115] +
//             mat_A[100] * mat_B[147] +
//             mat_A[101] * mat_B[179] +
//             mat_A[102] * mat_B[211] +
//             mat_A[103] * mat_B[243] +
//             mat_A[104] * mat_B[275] +
//             mat_A[105] * mat_B[307] +
//             mat_A[106] * mat_B[339] +
//             mat_A[107] * mat_B[371] +
//             mat_A[108] * mat_B[403] +
//             mat_A[109] * mat_B[435] +
//             mat_A[110] * mat_B[467] +
//             mat_A[111] * mat_B[499] +
//             mat_A[112] * mat_B[531] +
//             mat_A[113] * mat_B[563] +
//             mat_A[114] * mat_B[595] +
//             mat_A[115] * mat_B[627] +
//             mat_A[116] * mat_B[659] +
//             mat_A[117] * mat_B[691] +
//             mat_A[118] * mat_B[723] +
//             mat_A[119] * mat_B[755] +
//             mat_A[120] * mat_B[787] +
//             mat_A[121] * mat_B[819] +
//             mat_A[122] * mat_B[851] +
//             mat_A[123] * mat_B[883] +
//             mat_A[124] * mat_B[915] +
//             mat_A[125] * mat_B[947] +
//             mat_A[126] * mat_B[979] +
//             mat_A[127] * mat_B[1011];
//  mat_C[116] <= 
//             mat_A[96] * mat_B[20] +
//             mat_A[97] * mat_B[52] +
//             mat_A[98] * mat_B[84] +
//             mat_A[99] * mat_B[116] +
//             mat_A[100] * mat_B[148] +
//             mat_A[101] * mat_B[180] +
//             mat_A[102] * mat_B[212] +
//             mat_A[103] * mat_B[244] +
//             mat_A[104] * mat_B[276] +
//             mat_A[105] * mat_B[308] +
//             mat_A[106] * mat_B[340] +
//             mat_A[107] * mat_B[372] +
//             mat_A[108] * mat_B[404] +
//             mat_A[109] * mat_B[436] +
//             mat_A[110] * mat_B[468] +
//             mat_A[111] * mat_B[500] +
//             mat_A[112] * mat_B[532] +
//             mat_A[113] * mat_B[564] +
//             mat_A[114] * mat_B[596] +
//             mat_A[115] * mat_B[628] +
//             mat_A[116] * mat_B[660] +
//             mat_A[117] * mat_B[692] +
//             mat_A[118] * mat_B[724] +
//             mat_A[119] * mat_B[756] +
//             mat_A[120] * mat_B[788] +
//             mat_A[121] * mat_B[820] +
//             mat_A[122] * mat_B[852] +
//             mat_A[123] * mat_B[884] +
//             mat_A[124] * mat_B[916] +
//             mat_A[125] * mat_B[948] +
//             mat_A[126] * mat_B[980] +
//             mat_A[127] * mat_B[1012];
//  mat_C[117] <= 
//             mat_A[96] * mat_B[21] +
//             mat_A[97] * mat_B[53] +
//             mat_A[98] * mat_B[85] +
//             mat_A[99] * mat_B[117] +
//             mat_A[100] * mat_B[149] +
//             mat_A[101] * mat_B[181] +
//             mat_A[102] * mat_B[213] +
//             mat_A[103] * mat_B[245] +
//             mat_A[104] * mat_B[277] +
//             mat_A[105] * mat_B[309] +
//             mat_A[106] * mat_B[341] +
//             mat_A[107] * mat_B[373] +
//             mat_A[108] * mat_B[405] +
//             mat_A[109] * mat_B[437] +
//             mat_A[110] * mat_B[469] +
//             mat_A[111] * mat_B[501] +
//             mat_A[112] * mat_B[533] +
//             mat_A[113] * mat_B[565] +
//             mat_A[114] * mat_B[597] +
//             mat_A[115] * mat_B[629] +
//             mat_A[116] * mat_B[661] +
//             mat_A[117] * mat_B[693] +
//             mat_A[118] * mat_B[725] +
//             mat_A[119] * mat_B[757] +
//             mat_A[120] * mat_B[789] +
//             mat_A[121] * mat_B[821] +
//             mat_A[122] * mat_B[853] +
//             mat_A[123] * mat_B[885] +
//             mat_A[124] * mat_B[917] +
//             mat_A[125] * mat_B[949] +
//             mat_A[126] * mat_B[981] +
//             mat_A[127] * mat_B[1013];
//  mat_C[118] <= 
//             mat_A[96] * mat_B[22] +
//             mat_A[97] * mat_B[54] +
//             mat_A[98] * mat_B[86] +
//             mat_A[99] * mat_B[118] +
//             mat_A[100] * mat_B[150] +
//             mat_A[101] * mat_B[182] +
//             mat_A[102] * mat_B[214] +
//             mat_A[103] * mat_B[246] +
//             mat_A[104] * mat_B[278] +
//             mat_A[105] * mat_B[310] +
//             mat_A[106] * mat_B[342] +
//             mat_A[107] * mat_B[374] +
//             mat_A[108] * mat_B[406] +
//             mat_A[109] * mat_B[438] +
//             mat_A[110] * mat_B[470] +
//             mat_A[111] * mat_B[502] +
//             mat_A[112] * mat_B[534] +
//             mat_A[113] * mat_B[566] +
//             mat_A[114] * mat_B[598] +
//             mat_A[115] * mat_B[630] +
//             mat_A[116] * mat_B[662] +
//             mat_A[117] * mat_B[694] +
//             mat_A[118] * mat_B[726] +
//             mat_A[119] * mat_B[758] +
//             mat_A[120] * mat_B[790] +
//             mat_A[121] * mat_B[822] +
//             mat_A[122] * mat_B[854] +
//             mat_A[123] * mat_B[886] +
//             mat_A[124] * mat_B[918] +
//             mat_A[125] * mat_B[950] +
//             mat_A[126] * mat_B[982] +
//             mat_A[127] * mat_B[1014];
//  mat_C[119] <= 
//             mat_A[96] * mat_B[23] +
//             mat_A[97] * mat_B[55] +
//             mat_A[98] * mat_B[87] +
//             mat_A[99] * mat_B[119] +
//             mat_A[100] * mat_B[151] +
//             mat_A[101] * mat_B[183] +
//             mat_A[102] * mat_B[215] +
//             mat_A[103] * mat_B[247] +
//             mat_A[104] * mat_B[279] +
//             mat_A[105] * mat_B[311] +
//             mat_A[106] * mat_B[343] +
//             mat_A[107] * mat_B[375] +
//             mat_A[108] * mat_B[407] +
//             mat_A[109] * mat_B[439] +
//             mat_A[110] * mat_B[471] +
//             mat_A[111] * mat_B[503] +
//             mat_A[112] * mat_B[535] +
//             mat_A[113] * mat_B[567] +
//             mat_A[114] * mat_B[599] +
//             mat_A[115] * mat_B[631] +
//             mat_A[116] * mat_B[663] +
//             mat_A[117] * mat_B[695] +
//             mat_A[118] * mat_B[727] +
//             mat_A[119] * mat_B[759] +
//             mat_A[120] * mat_B[791] +
//             mat_A[121] * mat_B[823] +
//             mat_A[122] * mat_B[855] +
//             mat_A[123] * mat_B[887] +
//             mat_A[124] * mat_B[919] +
//             mat_A[125] * mat_B[951] +
//             mat_A[126] * mat_B[983] +
//             mat_A[127] * mat_B[1015];
//  mat_C[120] <= 
//             mat_A[96] * mat_B[24] +
//             mat_A[97] * mat_B[56] +
//             mat_A[98] * mat_B[88] +
//             mat_A[99] * mat_B[120] +
//             mat_A[100] * mat_B[152] +
//             mat_A[101] * mat_B[184] +
//             mat_A[102] * mat_B[216] +
//             mat_A[103] * mat_B[248] +
//             mat_A[104] * mat_B[280] +
//             mat_A[105] * mat_B[312] +
//             mat_A[106] * mat_B[344] +
//             mat_A[107] * mat_B[376] +
//             mat_A[108] * mat_B[408] +
//             mat_A[109] * mat_B[440] +
//             mat_A[110] * mat_B[472] +
//             mat_A[111] * mat_B[504] +
//             mat_A[112] * mat_B[536] +
//             mat_A[113] * mat_B[568] +
//             mat_A[114] * mat_B[600] +
//             mat_A[115] * mat_B[632] +
//             mat_A[116] * mat_B[664] +
//             mat_A[117] * mat_B[696] +
//             mat_A[118] * mat_B[728] +
//             mat_A[119] * mat_B[760] +
//             mat_A[120] * mat_B[792] +
//             mat_A[121] * mat_B[824] +
//             mat_A[122] * mat_B[856] +
//             mat_A[123] * mat_B[888] +
//             mat_A[124] * mat_B[920] +
//             mat_A[125] * mat_B[952] +
//             mat_A[126] * mat_B[984] +
//             mat_A[127] * mat_B[1016];
//  mat_C[121] <= 
//             mat_A[96] * mat_B[25] +
//             mat_A[97] * mat_B[57] +
//             mat_A[98] * mat_B[89] +
//             mat_A[99] * mat_B[121] +
//             mat_A[100] * mat_B[153] +
//             mat_A[101] * mat_B[185] +
//             mat_A[102] * mat_B[217] +
//             mat_A[103] * mat_B[249] +
//             mat_A[104] * mat_B[281] +
//             mat_A[105] * mat_B[313] +
//             mat_A[106] * mat_B[345] +
//             mat_A[107] * mat_B[377] +
//             mat_A[108] * mat_B[409] +
//             mat_A[109] * mat_B[441] +
//             mat_A[110] * mat_B[473] +
//             mat_A[111] * mat_B[505] +
//             mat_A[112] * mat_B[537] +
//             mat_A[113] * mat_B[569] +
//             mat_A[114] * mat_B[601] +
//             mat_A[115] * mat_B[633] +
//             mat_A[116] * mat_B[665] +
//             mat_A[117] * mat_B[697] +
//             mat_A[118] * mat_B[729] +
//             mat_A[119] * mat_B[761] +
//             mat_A[120] * mat_B[793] +
//             mat_A[121] * mat_B[825] +
//             mat_A[122] * mat_B[857] +
//             mat_A[123] * mat_B[889] +
//             mat_A[124] * mat_B[921] +
//             mat_A[125] * mat_B[953] +
//             mat_A[126] * mat_B[985] +
//             mat_A[127] * mat_B[1017];
//  mat_C[122] <= 
//             mat_A[96] * mat_B[26] +
//             mat_A[97] * mat_B[58] +
//             mat_A[98] * mat_B[90] +
//             mat_A[99] * mat_B[122] +
//             mat_A[100] * mat_B[154] +
//             mat_A[101] * mat_B[186] +
//             mat_A[102] * mat_B[218] +
//             mat_A[103] * mat_B[250] +
//             mat_A[104] * mat_B[282] +
//             mat_A[105] * mat_B[314] +
//             mat_A[106] * mat_B[346] +
//             mat_A[107] * mat_B[378] +
//             mat_A[108] * mat_B[410] +
//             mat_A[109] * mat_B[442] +
//             mat_A[110] * mat_B[474] +
//             mat_A[111] * mat_B[506] +
//             mat_A[112] * mat_B[538] +
//             mat_A[113] * mat_B[570] +
//             mat_A[114] * mat_B[602] +
//             mat_A[115] * mat_B[634] +
//             mat_A[116] * mat_B[666] +
//             mat_A[117] * mat_B[698] +
//             mat_A[118] * mat_B[730] +
//             mat_A[119] * mat_B[762] +
//             mat_A[120] * mat_B[794] +
//             mat_A[121] * mat_B[826] +
//             mat_A[122] * mat_B[858] +
//             mat_A[123] * mat_B[890] +
//             mat_A[124] * mat_B[922] +
//             mat_A[125] * mat_B[954] +
//             mat_A[126] * mat_B[986] +
//             mat_A[127] * mat_B[1018];
//  mat_C[123] <= 
//             mat_A[96] * mat_B[27] +
//             mat_A[97] * mat_B[59] +
//             mat_A[98] * mat_B[91] +
//             mat_A[99] * mat_B[123] +
//             mat_A[100] * mat_B[155] +
//             mat_A[101] * mat_B[187] +
//             mat_A[102] * mat_B[219] +
//             mat_A[103] * mat_B[251] +
//             mat_A[104] * mat_B[283] +
//             mat_A[105] * mat_B[315] +
//             mat_A[106] * mat_B[347] +
//             mat_A[107] * mat_B[379] +
//             mat_A[108] * mat_B[411] +
//             mat_A[109] * mat_B[443] +
//             mat_A[110] * mat_B[475] +
//             mat_A[111] * mat_B[507] +
//             mat_A[112] * mat_B[539] +
//             mat_A[113] * mat_B[571] +
//             mat_A[114] * mat_B[603] +
//             mat_A[115] * mat_B[635] +
//             mat_A[116] * mat_B[667] +
//             mat_A[117] * mat_B[699] +
//             mat_A[118] * mat_B[731] +
//             mat_A[119] * mat_B[763] +
//             mat_A[120] * mat_B[795] +
//             mat_A[121] * mat_B[827] +
//             mat_A[122] * mat_B[859] +
//             mat_A[123] * mat_B[891] +
//             mat_A[124] * mat_B[923] +
//             mat_A[125] * mat_B[955] +
//             mat_A[126] * mat_B[987] +
//             mat_A[127] * mat_B[1019];
//  mat_C[124] <= 
//             mat_A[96] * mat_B[28] +
//             mat_A[97] * mat_B[60] +
//             mat_A[98] * mat_B[92] +
//             mat_A[99] * mat_B[124] +
//             mat_A[100] * mat_B[156] +
//             mat_A[101] * mat_B[188] +
//             mat_A[102] * mat_B[220] +
//             mat_A[103] * mat_B[252] +
//             mat_A[104] * mat_B[284] +
//             mat_A[105] * mat_B[316] +
//             mat_A[106] * mat_B[348] +
//             mat_A[107] * mat_B[380] +
//             mat_A[108] * mat_B[412] +
//             mat_A[109] * mat_B[444] +
//             mat_A[110] * mat_B[476] +
//             mat_A[111] * mat_B[508] +
//             mat_A[112] * mat_B[540] +
//             mat_A[113] * mat_B[572] +
//             mat_A[114] * mat_B[604] +
//             mat_A[115] * mat_B[636] +
//             mat_A[116] * mat_B[668] +
//             mat_A[117] * mat_B[700] +
//             mat_A[118] * mat_B[732] +
//             mat_A[119] * mat_B[764] +
//             mat_A[120] * mat_B[796] +
//             mat_A[121] * mat_B[828] +
//             mat_A[122] * mat_B[860] +
//             mat_A[123] * mat_B[892] +
//             mat_A[124] * mat_B[924] +
//             mat_A[125] * mat_B[956] +
//             mat_A[126] * mat_B[988] +
//             mat_A[127] * mat_B[1020];
//  mat_C[125] <= 
//             mat_A[96] * mat_B[29] +
//             mat_A[97] * mat_B[61] +
//             mat_A[98] * mat_B[93] +
//             mat_A[99] * mat_B[125] +
//             mat_A[100] * mat_B[157] +
//             mat_A[101] * mat_B[189] +
//             mat_A[102] * mat_B[221] +
//             mat_A[103] * mat_B[253] +
//             mat_A[104] * mat_B[285] +
//             mat_A[105] * mat_B[317] +
//             mat_A[106] * mat_B[349] +
//             mat_A[107] * mat_B[381] +
//             mat_A[108] * mat_B[413] +
//             mat_A[109] * mat_B[445] +
//             mat_A[110] * mat_B[477] +
//             mat_A[111] * mat_B[509] +
//             mat_A[112] * mat_B[541] +
//             mat_A[113] * mat_B[573] +
//             mat_A[114] * mat_B[605] +
//             mat_A[115] * mat_B[637] +
//             mat_A[116] * mat_B[669] +
//             mat_A[117] * mat_B[701] +
//             mat_A[118] * mat_B[733] +
//             mat_A[119] * mat_B[765] +
//             mat_A[120] * mat_B[797] +
//             mat_A[121] * mat_B[829] +
//             mat_A[122] * mat_B[861] +
//             mat_A[123] * mat_B[893] +
//             mat_A[124] * mat_B[925] +
//             mat_A[125] * mat_B[957] +
//             mat_A[126] * mat_B[989] +
//             mat_A[127] * mat_B[1021];
//  mat_C[126] <= 
//             mat_A[96] * mat_B[30] +
//             mat_A[97] * mat_B[62] +
//             mat_A[98] * mat_B[94] +
//             mat_A[99] * mat_B[126] +
//             mat_A[100] * mat_B[158] +
//             mat_A[101] * mat_B[190] +
//             mat_A[102] * mat_B[222] +
//             mat_A[103] * mat_B[254] +
//             mat_A[104] * mat_B[286] +
//             mat_A[105] * mat_B[318] +
//             mat_A[106] * mat_B[350] +
//             mat_A[107] * mat_B[382] +
//             mat_A[108] * mat_B[414] +
//             mat_A[109] * mat_B[446] +
//             mat_A[110] * mat_B[478] +
//             mat_A[111] * mat_B[510] +
//             mat_A[112] * mat_B[542] +
//             mat_A[113] * mat_B[574] +
//             mat_A[114] * mat_B[606] +
//             mat_A[115] * mat_B[638] +
//             mat_A[116] * mat_B[670] +
//             mat_A[117] * mat_B[702] +
//             mat_A[118] * mat_B[734] +
//             mat_A[119] * mat_B[766] +
//             mat_A[120] * mat_B[798] +
//             mat_A[121] * mat_B[830] +
//             mat_A[122] * mat_B[862] +
//             mat_A[123] * mat_B[894] +
//             mat_A[124] * mat_B[926] +
//             mat_A[125] * mat_B[958] +
//             mat_A[126] * mat_B[990] +
//             mat_A[127] * mat_B[1022];
//  mat_C[127] <= 
//             mat_A[96] * mat_B[31] +
//             mat_A[97] * mat_B[63] +
//             mat_A[98] * mat_B[95] +
//             mat_A[99] * mat_B[127] +
//             mat_A[100] * mat_B[159] +
//             mat_A[101] * mat_B[191] +
//             mat_A[102] * mat_B[223] +
//             mat_A[103] * mat_B[255] +
//             mat_A[104] * mat_B[287] +
//             mat_A[105] * mat_B[319] +
//             mat_A[106] * mat_B[351] +
//             mat_A[107] * mat_B[383] +
//             mat_A[108] * mat_B[415] +
//             mat_A[109] * mat_B[447] +
//             mat_A[110] * mat_B[479] +
//             mat_A[111] * mat_B[511] +
//             mat_A[112] * mat_B[543] +
//             mat_A[113] * mat_B[575] +
//             mat_A[114] * mat_B[607] +
//             mat_A[115] * mat_B[639] +
//             mat_A[116] * mat_B[671] +
//             mat_A[117] * mat_B[703] +
//             mat_A[118] * mat_B[735] +
//             mat_A[119] * mat_B[767] +
//             mat_A[120] * mat_B[799] +
//             mat_A[121] * mat_B[831] +
//             mat_A[122] * mat_B[863] +
//             mat_A[123] * mat_B[895] +
//             mat_A[124] * mat_B[927] +
//             mat_A[125] * mat_B[959] +
//             mat_A[126] * mat_B[991] +
//             mat_A[127] * mat_B[1023];
//  mat_C[128] <= 
//             mat_A[128] * mat_B[0] +
//             mat_A[129] * mat_B[32] +
//             mat_A[130] * mat_B[64] +
//             mat_A[131] * mat_B[96] +
//             mat_A[132] * mat_B[128] +
//             mat_A[133] * mat_B[160] +
//             mat_A[134] * mat_B[192] +
//             mat_A[135] * mat_B[224] +
//             mat_A[136] * mat_B[256] +
//             mat_A[137] * mat_B[288] +
//             mat_A[138] * mat_B[320] +
//             mat_A[139] * mat_B[352] +
//             mat_A[140] * mat_B[384] +
//             mat_A[141] * mat_B[416] +
//             mat_A[142] * mat_B[448] +
//             mat_A[143] * mat_B[480] +
//             mat_A[144] * mat_B[512] +
//             mat_A[145] * mat_B[544] +
//             mat_A[146] * mat_B[576] +
//             mat_A[147] * mat_B[608] +
//             mat_A[148] * mat_B[640] +
//             mat_A[149] * mat_B[672] +
//             mat_A[150] * mat_B[704] +
//             mat_A[151] * mat_B[736] +
//             mat_A[152] * mat_B[768] +
//             mat_A[153] * mat_B[800] +
//             mat_A[154] * mat_B[832] +
//             mat_A[155] * mat_B[864] +
//             mat_A[156] * mat_B[896] +
//             mat_A[157] * mat_B[928] +
//             mat_A[158] * mat_B[960] +
//             mat_A[159] * mat_B[992];
//  mat_C[129] <= 
//             mat_A[128] * mat_B[1] +
//             mat_A[129] * mat_B[33] +
//             mat_A[130] * mat_B[65] +
//             mat_A[131] * mat_B[97] +
//             mat_A[132] * mat_B[129] +
//             mat_A[133] * mat_B[161] +
//             mat_A[134] * mat_B[193] +
//             mat_A[135] * mat_B[225] +
//             mat_A[136] * mat_B[257] +
//             mat_A[137] * mat_B[289] +
//             mat_A[138] * mat_B[321] +
//             mat_A[139] * mat_B[353] +
//             mat_A[140] * mat_B[385] +
//             mat_A[141] * mat_B[417] +
//             mat_A[142] * mat_B[449] +
//             mat_A[143] * mat_B[481] +
//             mat_A[144] * mat_B[513] +
//             mat_A[145] * mat_B[545] +
//             mat_A[146] * mat_B[577] +
//             mat_A[147] * mat_B[609] +
//             mat_A[148] * mat_B[641] +
//             mat_A[149] * mat_B[673] +
//             mat_A[150] * mat_B[705] +
//             mat_A[151] * mat_B[737] +
//             mat_A[152] * mat_B[769] +
//             mat_A[153] * mat_B[801] +
//             mat_A[154] * mat_B[833] +
//             mat_A[155] * mat_B[865] +
//             mat_A[156] * mat_B[897] +
//             mat_A[157] * mat_B[929] +
//             mat_A[158] * mat_B[961] +
//             mat_A[159] * mat_B[993];
//  mat_C[130] <= 
//             mat_A[128] * mat_B[2] +
//             mat_A[129] * mat_B[34] +
//             mat_A[130] * mat_B[66] +
//             mat_A[131] * mat_B[98] +
//             mat_A[132] * mat_B[130] +
//             mat_A[133] * mat_B[162] +
//             mat_A[134] * mat_B[194] +
//             mat_A[135] * mat_B[226] +
//             mat_A[136] * mat_B[258] +
//             mat_A[137] * mat_B[290] +
//             mat_A[138] * mat_B[322] +
//             mat_A[139] * mat_B[354] +
//             mat_A[140] * mat_B[386] +
//             mat_A[141] * mat_B[418] +
//             mat_A[142] * mat_B[450] +
//             mat_A[143] * mat_B[482] +
//             mat_A[144] * mat_B[514] +
//             mat_A[145] * mat_B[546] +
//             mat_A[146] * mat_B[578] +
//             mat_A[147] * mat_B[610] +
//             mat_A[148] * mat_B[642] +
//             mat_A[149] * mat_B[674] +
//             mat_A[150] * mat_B[706] +
//             mat_A[151] * mat_B[738] +
//             mat_A[152] * mat_B[770] +
//             mat_A[153] * mat_B[802] +
//             mat_A[154] * mat_B[834] +
//             mat_A[155] * mat_B[866] +
//             mat_A[156] * mat_B[898] +
//             mat_A[157] * mat_B[930] +
//             mat_A[158] * mat_B[962] +
//             mat_A[159] * mat_B[994];
//  mat_C[131] <= 
//             mat_A[128] * mat_B[3] +
//             mat_A[129] * mat_B[35] +
//             mat_A[130] * mat_B[67] +
//             mat_A[131] * mat_B[99] +
//             mat_A[132] * mat_B[131] +
//             mat_A[133] * mat_B[163] +
//             mat_A[134] * mat_B[195] +
//             mat_A[135] * mat_B[227] +
//             mat_A[136] * mat_B[259] +
//             mat_A[137] * mat_B[291] +
//             mat_A[138] * mat_B[323] +
//             mat_A[139] * mat_B[355] +
//             mat_A[140] * mat_B[387] +
//             mat_A[141] * mat_B[419] +
//             mat_A[142] * mat_B[451] +
//             mat_A[143] * mat_B[483] +
//             mat_A[144] * mat_B[515] +
//             mat_A[145] * mat_B[547] +
//             mat_A[146] * mat_B[579] +
//             mat_A[147] * mat_B[611] +
//             mat_A[148] * mat_B[643] +
//             mat_A[149] * mat_B[675] +
//             mat_A[150] * mat_B[707] +
//             mat_A[151] * mat_B[739] +
//             mat_A[152] * mat_B[771] +
//             mat_A[153] * mat_B[803] +
//             mat_A[154] * mat_B[835] +
//             mat_A[155] * mat_B[867] +
//             mat_A[156] * mat_B[899] +
//             mat_A[157] * mat_B[931] +
//             mat_A[158] * mat_B[963] +
//             mat_A[159] * mat_B[995];
//  mat_C[132] <= 
//             mat_A[128] * mat_B[4] +
//             mat_A[129] * mat_B[36] +
//             mat_A[130] * mat_B[68] +
//             mat_A[131] * mat_B[100] +
//             mat_A[132] * mat_B[132] +
//             mat_A[133] * mat_B[164] +
//             mat_A[134] * mat_B[196] +
//             mat_A[135] * mat_B[228] +
//             mat_A[136] * mat_B[260] +
//             mat_A[137] * mat_B[292] +
//             mat_A[138] * mat_B[324] +
//             mat_A[139] * mat_B[356] +
//             mat_A[140] * mat_B[388] +
//             mat_A[141] * mat_B[420] +
//             mat_A[142] * mat_B[452] +
//             mat_A[143] * mat_B[484] +
//             mat_A[144] * mat_B[516] +
//             mat_A[145] * mat_B[548] +
//             mat_A[146] * mat_B[580] +
//             mat_A[147] * mat_B[612] +
//             mat_A[148] * mat_B[644] +
//             mat_A[149] * mat_B[676] +
//             mat_A[150] * mat_B[708] +
//             mat_A[151] * mat_B[740] +
//             mat_A[152] * mat_B[772] +
//             mat_A[153] * mat_B[804] +
//             mat_A[154] * mat_B[836] +
//             mat_A[155] * mat_B[868] +
//             mat_A[156] * mat_B[900] +
//             mat_A[157] * mat_B[932] +
//             mat_A[158] * mat_B[964] +
//             mat_A[159] * mat_B[996];
//  mat_C[133] <= 
//             mat_A[128] * mat_B[5] +
//             mat_A[129] * mat_B[37] +
//             mat_A[130] * mat_B[69] +
//             mat_A[131] * mat_B[101] +
//             mat_A[132] * mat_B[133] +
//             mat_A[133] * mat_B[165] +
//             mat_A[134] * mat_B[197] +
//             mat_A[135] * mat_B[229] +
//             mat_A[136] * mat_B[261] +
//             mat_A[137] * mat_B[293] +
//             mat_A[138] * mat_B[325] +
//             mat_A[139] * mat_B[357] +
//             mat_A[140] * mat_B[389] +
//             mat_A[141] * mat_B[421] +
//             mat_A[142] * mat_B[453] +
//             mat_A[143] * mat_B[485] +
//             mat_A[144] * mat_B[517] +
//             mat_A[145] * mat_B[549] +
//             mat_A[146] * mat_B[581] +
//             mat_A[147] * mat_B[613] +
//             mat_A[148] * mat_B[645] +
//             mat_A[149] * mat_B[677] +
//             mat_A[150] * mat_B[709] +
//             mat_A[151] * mat_B[741] +
//             mat_A[152] * mat_B[773] +
//             mat_A[153] * mat_B[805] +
//             mat_A[154] * mat_B[837] +
//             mat_A[155] * mat_B[869] +
//             mat_A[156] * mat_B[901] +
//             mat_A[157] * mat_B[933] +
//             mat_A[158] * mat_B[965] +
//             mat_A[159] * mat_B[997];
//  mat_C[134] <= 
//             mat_A[128] * mat_B[6] +
//             mat_A[129] * mat_B[38] +
//             mat_A[130] * mat_B[70] +
//             mat_A[131] * mat_B[102] +
//             mat_A[132] * mat_B[134] +
//             mat_A[133] * mat_B[166] +
//             mat_A[134] * mat_B[198] +
//             mat_A[135] * mat_B[230] +
//             mat_A[136] * mat_B[262] +
//             mat_A[137] * mat_B[294] +
//             mat_A[138] * mat_B[326] +
//             mat_A[139] * mat_B[358] +
//             mat_A[140] * mat_B[390] +
//             mat_A[141] * mat_B[422] +
//             mat_A[142] * mat_B[454] +
//             mat_A[143] * mat_B[486] +
//             mat_A[144] * mat_B[518] +
//             mat_A[145] * mat_B[550] +
//             mat_A[146] * mat_B[582] +
//             mat_A[147] * mat_B[614] +
//             mat_A[148] * mat_B[646] +
//             mat_A[149] * mat_B[678] +
//             mat_A[150] * mat_B[710] +
//             mat_A[151] * mat_B[742] +
//             mat_A[152] * mat_B[774] +
//             mat_A[153] * mat_B[806] +
//             mat_A[154] * mat_B[838] +
//             mat_A[155] * mat_B[870] +
//             mat_A[156] * mat_B[902] +
//             mat_A[157] * mat_B[934] +
//             mat_A[158] * mat_B[966] +
//             mat_A[159] * mat_B[998];
//  mat_C[135] <= 
//             mat_A[128] * mat_B[7] +
//             mat_A[129] * mat_B[39] +
//             mat_A[130] * mat_B[71] +
//             mat_A[131] * mat_B[103] +
//             mat_A[132] * mat_B[135] +
//             mat_A[133] * mat_B[167] +
//             mat_A[134] * mat_B[199] +
//             mat_A[135] * mat_B[231] +
//             mat_A[136] * mat_B[263] +
//             mat_A[137] * mat_B[295] +
//             mat_A[138] * mat_B[327] +
//             mat_A[139] * mat_B[359] +
//             mat_A[140] * mat_B[391] +
//             mat_A[141] * mat_B[423] +
//             mat_A[142] * mat_B[455] +
//             mat_A[143] * mat_B[487] +
//             mat_A[144] * mat_B[519] +
//             mat_A[145] * mat_B[551] +
//             mat_A[146] * mat_B[583] +
//             mat_A[147] * mat_B[615] +
//             mat_A[148] * mat_B[647] +
//             mat_A[149] * mat_B[679] +
//             mat_A[150] * mat_B[711] +
//             mat_A[151] * mat_B[743] +
//             mat_A[152] * mat_B[775] +
//             mat_A[153] * mat_B[807] +
//             mat_A[154] * mat_B[839] +
//             mat_A[155] * mat_B[871] +
//             mat_A[156] * mat_B[903] +
//             mat_A[157] * mat_B[935] +
//             mat_A[158] * mat_B[967] +
//             mat_A[159] * mat_B[999];
//  mat_C[136] <= 
//             mat_A[128] * mat_B[8] +
//             mat_A[129] * mat_B[40] +
//             mat_A[130] * mat_B[72] +
//             mat_A[131] * mat_B[104] +
//             mat_A[132] * mat_B[136] +
//             mat_A[133] * mat_B[168] +
//             mat_A[134] * mat_B[200] +
//             mat_A[135] * mat_B[232] +
//             mat_A[136] * mat_B[264] +
//             mat_A[137] * mat_B[296] +
//             mat_A[138] * mat_B[328] +
//             mat_A[139] * mat_B[360] +
//             mat_A[140] * mat_B[392] +
//             mat_A[141] * mat_B[424] +
//             mat_A[142] * mat_B[456] +
//             mat_A[143] * mat_B[488] +
//             mat_A[144] * mat_B[520] +
//             mat_A[145] * mat_B[552] +
//             mat_A[146] * mat_B[584] +
//             mat_A[147] * mat_B[616] +
//             mat_A[148] * mat_B[648] +
//             mat_A[149] * mat_B[680] +
//             mat_A[150] * mat_B[712] +
//             mat_A[151] * mat_B[744] +
//             mat_A[152] * mat_B[776] +
//             mat_A[153] * mat_B[808] +
//             mat_A[154] * mat_B[840] +
//             mat_A[155] * mat_B[872] +
//             mat_A[156] * mat_B[904] +
//             mat_A[157] * mat_B[936] +
//             mat_A[158] * mat_B[968] +
//             mat_A[159] * mat_B[1000];
//  mat_C[137] <= 
//             mat_A[128] * mat_B[9] +
//             mat_A[129] * mat_B[41] +
//             mat_A[130] * mat_B[73] +
//             mat_A[131] * mat_B[105] +
//             mat_A[132] * mat_B[137] +
//             mat_A[133] * mat_B[169] +
//             mat_A[134] * mat_B[201] +
//             mat_A[135] * mat_B[233] +
//             mat_A[136] * mat_B[265] +
//             mat_A[137] * mat_B[297] +
//             mat_A[138] * mat_B[329] +
//             mat_A[139] * mat_B[361] +
//             mat_A[140] * mat_B[393] +
//             mat_A[141] * mat_B[425] +
//             mat_A[142] * mat_B[457] +
//             mat_A[143] * mat_B[489] +
//             mat_A[144] * mat_B[521] +
//             mat_A[145] * mat_B[553] +
//             mat_A[146] * mat_B[585] +
//             mat_A[147] * mat_B[617] +
//             mat_A[148] * mat_B[649] +
//             mat_A[149] * mat_B[681] +
//             mat_A[150] * mat_B[713] +
//             mat_A[151] * mat_B[745] +
//             mat_A[152] * mat_B[777] +
//             mat_A[153] * mat_B[809] +
//             mat_A[154] * mat_B[841] +
//             mat_A[155] * mat_B[873] +
//             mat_A[156] * mat_B[905] +
//             mat_A[157] * mat_B[937] +
//             mat_A[158] * mat_B[969] +
//             mat_A[159] * mat_B[1001];
//  mat_C[138] <= 
//             mat_A[128] * mat_B[10] +
//             mat_A[129] * mat_B[42] +
//             mat_A[130] * mat_B[74] +
//             mat_A[131] * mat_B[106] +
//             mat_A[132] * mat_B[138] +
//             mat_A[133] * mat_B[170] +
//             mat_A[134] * mat_B[202] +
//             mat_A[135] * mat_B[234] +
//             mat_A[136] * mat_B[266] +
//             mat_A[137] * mat_B[298] +
//             mat_A[138] * mat_B[330] +
//             mat_A[139] * mat_B[362] +
//             mat_A[140] * mat_B[394] +
//             mat_A[141] * mat_B[426] +
//             mat_A[142] * mat_B[458] +
//             mat_A[143] * mat_B[490] +
//             mat_A[144] * mat_B[522] +
//             mat_A[145] * mat_B[554] +
//             mat_A[146] * mat_B[586] +
//             mat_A[147] * mat_B[618] +
//             mat_A[148] * mat_B[650] +
//             mat_A[149] * mat_B[682] +
//             mat_A[150] * mat_B[714] +
//             mat_A[151] * mat_B[746] +
//             mat_A[152] * mat_B[778] +
//             mat_A[153] * mat_B[810] +
//             mat_A[154] * mat_B[842] +
//             mat_A[155] * mat_B[874] +
//             mat_A[156] * mat_B[906] +
//             mat_A[157] * mat_B[938] +
//             mat_A[158] * mat_B[970] +
//             mat_A[159] * mat_B[1002];
//  mat_C[139] <= 
//             mat_A[128] * mat_B[11] +
//             mat_A[129] * mat_B[43] +
//             mat_A[130] * mat_B[75] +
//             mat_A[131] * mat_B[107] +
//             mat_A[132] * mat_B[139] +
//             mat_A[133] * mat_B[171] +
//             mat_A[134] * mat_B[203] +
//             mat_A[135] * mat_B[235] +
//             mat_A[136] * mat_B[267] +
//             mat_A[137] * mat_B[299] +
//             mat_A[138] * mat_B[331] +
//             mat_A[139] * mat_B[363] +
//             mat_A[140] * mat_B[395] +
//             mat_A[141] * mat_B[427] +
//             mat_A[142] * mat_B[459] +
//             mat_A[143] * mat_B[491] +
//             mat_A[144] * mat_B[523] +
//             mat_A[145] * mat_B[555] +
//             mat_A[146] * mat_B[587] +
//             mat_A[147] * mat_B[619] +
//             mat_A[148] * mat_B[651] +
//             mat_A[149] * mat_B[683] +
//             mat_A[150] * mat_B[715] +
//             mat_A[151] * mat_B[747] +
//             mat_A[152] * mat_B[779] +
//             mat_A[153] * mat_B[811] +
//             mat_A[154] * mat_B[843] +
//             mat_A[155] * mat_B[875] +
//             mat_A[156] * mat_B[907] +
//             mat_A[157] * mat_B[939] +
//             mat_A[158] * mat_B[971] +
//             mat_A[159] * mat_B[1003];
//  mat_C[140] <= 
//             mat_A[128] * mat_B[12] +
//             mat_A[129] * mat_B[44] +
//             mat_A[130] * mat_B[76] +
//             mat_A[131] * mat_B[108] +
//             mat_A[132] * mat_B[140] +
//             mat_A[133] * mat_B[172] +
//             mat_A[134] * mat_B[204] +
//             mat_A[135] * mat_B[236] +
//             mat_A[136] * mat_B[268] +
//             mat_A[137] * mat_B[300] +
//             mat_A[138] * mat_B[332] +
//             mat_A[139] * mat_B[364] +
//             mat_A[140] * mat_B[396] +
//             mat_A[141] * mat_B[428] +
//             mat_A[142] * mat_B[460] +
//             mat_A[143] * mat_B[492] +
//             mat_A[144] * mat_B[524] +
//             mat_A[145] * mat_B[556] +
//             mat_A[146] * mat_B[588] +
//             mat_A[147] * mat_B[620] +
//             mat_A[148] * mat_B[652] +
//             mat_A[149] * mat_B[684] +
//             mat_A[150] * mat_B[716] +
//             mat_A[151] * mat_B[748] +
//             mat_A[152] * mat_B[780] +
//             mat_A[153] * mat_B[812] +
//             mat_A[154] * mat_B[844] +
//             mat_A[155] * mat_B[876] +
//             mat_A[156] * mat_B[908] +
//             mat_A[157] * mat_B[940] +
//             mat_A[158] * mat_B[972] +
//             mat_A[159] * mat_B[1004];
//  mat_C[141] <= 
//             mat_A[128] * mat_B[13] +
//             mat_A[129] * mat_B[45] +
//             mat_A[130] * mat_B[77] +
//             mat_A[131] * mat_B[109] +
//             mat_A[132] * mat_B[141] +
//             mat_A[133] * mat_B[173] +
//             mat_A[134] * mat_B[205] +
//             mat_A[135] * mat_B[237] +
//             mat_A[136] * mat_B[269] +
//             mat_A[137] * mat_B[301] +
//             mat_A[138] * mat_B[333] +
//             mat_A[139] * mat_B[365] +
//             mat_A[140] * mat_B[397] +
//             mat_A[141] * mat_B[429] +
//             mat_A[142] * mat_B[461] +
//             mat_A[143] * mat_B[493] +
//             mat_A[144] * mat_B[525] +
//             mat_A[145] * mat_B[557] +
//             mat_A[146] * mat_B[589] +
//             mat_A[147] * mat_B[621] +
//             mat_A[148] * mat_B[653] +
//             mat_A[149] * mat_B[685] +
//             mat_A[150] * mat_B[717] +
//             mat_A[151] * mat_B[749] +
//             mat_A[152] * mat_B[781] +
//             mat_A[153] * mat_B[813] +
//             mat_A[154] * mat_B[845] +
//             mat_A[155] * mat_B[877] +
//             mat_A[156] * mat_B[909] +
//             mat_A[157] * mat_B[941] +
//             mat_A[158] * mat_B[973] +
//             mat_A[159] * mat_B[1005];
//  mat_C[142] <= 
//             mat_A[128] * mat_B[14] +
//             mat_A[129] * mat_B[46] +
//             mat_A[130] * mat_B[78] +
//             mat_A[131] * mat_B[110] +
//             mat_A[132] * mat_B[142] +
//             mat_A[133] * mat_B[174] +
//             mat_A[134] * mat_B[206] +
//             mat_A[135] * mat_B[238] +
//             mat_A[136] * mat_B[270] +
//             mat_A[137] * mat_B[302] +
//             mat_A[138] * mat_B[334] +
//             mat_A[139] * mat_B[366] +
//             mat_A[140] * mat_B[398] +
//             mat_A[141] * mat_B[430] +
//             mat_A[142] * mat_B[462] +
//             mat_A[143] * mat_B[494] +
//             mat_A[144] * mat_B[526] +
//             mat_A[145] * mat_B[558] +
//             mat_A[146] * mat_B[590] +
//             mat_A[147] * mat_B[622] +
//             mat_A[148] * mat_B[654] +
//             mat_A[149] * mat_B[686] +
//             mat_A[150] * mat_B[718] +
//             mat_A[151] * mat_B[750] +
//             mat_A[152] * mat_B[782] +
//             mat_A[153] * mat_B[814] +
//             mat_A[154] * mat_B[846] +
//             mat_A[155] * mat_B[878] +
//             mat_A[156] * mat_B[910] +
//             mat_A[157] * mat_B[942] +
//             mat_A[158] * mat_B[974] +
//             mat_A[159] * mat_B[1006];
//  mat_C[143] <= 
//             mat_A[128] * mat_B[15] +
//             mat_A[129] * mat_B[47] +
//             mat_A[130] * mat_B[79] +
//             mat_A[131] * mat_B[111] +
//             mat_A[132] * mat_B[143] +
//             mat_A[133] * mat_B[175] +
//             mat_A[134] * mat_B[207] +
//             mat_A[135] * mat_B[239] +
//             mat_A[136] * mat_B[271] +
//             mat_A[137] * mat_B[303] +
//             mat_A[138] * mat_B[335] +
//             mat_A[139] * mat_B[367] +
//             mat_A[140] * mat_B[399] +
//             mat_A[141] * mat_B[431] +
//             mat_A[142] * mat_B[463] +
//             mat_A[143] * mat_B[495] +
//             mat_A[144] * mat_B[527] +
//             mat_A[145] * mat_B[559] +
//             mat_A[146] * mat_B[591] +
//             mat_A[147] * mat_B[623] +
//             mat_A[148] * mat_B[655] +
//             mat_A[149] * mat_B[687] +
//             mat_A[150] * mat_B[719] +
//             mat_A[151] * mat_B[751] +
//             mat_A[152] * mat_B[783] +
//             mat_A[153] * mat_B[815] +
//             mat_A[154] * mat_B[847] +
//             mat_A[155] * mat_B[879] +
//             mat_A[156] * mat_B[911] +
//             mat_A[157] * mat_B[943] +
//             mat_A[158] * mat_B[975] +
//             mat_A[159] * mat_B[1007];
//  mat_C[144] <= 
//             mat_A[128] * mat_B[16] +
//             mat_A[129] * mat_B[48] +
//             mat_A[130] * mat_B[80] +
//             mat_A[131] * mat_B[112] +
//             mat_A[132] * mat_B[144] +
//             mat_A[133] * mat_B[176] +
//             mat_A[134] * mat_B[208] +
//             mat_A[135] * mat_B[240] +
//             mat_A[136] * mat_B[272] +
//             mat_A[137] * mat_B[304] +
//             mat_A[138] * mat_B[336] +
//             mat_A[139] * mat_B[368] +
//             mat_A[140] * mat_B[400] +
//             mat_A[141] * mat_B[432] +
//             mat_A[142] * mat_B[464] +
//             mat_A[143] * mat_B[496] +
//             mat_A[144] * mat_B[528] +
//             mat_A[145] * mat_B[560] +
//             mat_A[146] * mat_B[592] +
//             mat_A[147] * mat_B[624] +
//             mat_A[148] * mat_B[656] +
//             mat_A[149] * mat_B[688] +
//             mat_A[150] * mat_B[720] +
//             mat_A[151] * mat_B[752] +
//             mat_A[152] * mat_B[784] +
//             mat_A[153] * mat_B[816] +
//             mat_A[154] * mat_B[848] +
//             mat_A[155] * mat_B[880] +
//             mat_A[156] * mat_B[912] +
//             mat_A[157] * mat_B[944] +
//             mat_A[158] * mat_B[976] +
//             mat_A[159] * mat_B[1008];
//  mat_C[145] <= 
//             mat_A[128] * mat_B[17] +
//             mat_A[129] * mat_B[49] +
//             mat_A[130] * mat_B[81] +
//             mat_A[131] * mat_B[113] +
//             mat_A[132] * mat_B[145] +
//             mat_A[133] * mat_B[177] +
//             mat_A[134] * mat_B[209] +
//             mat_A[135] * mat_B[241] +
//             mat_A[136] * mat_B[273] +
//             mat_A[137] * mat_B[305] +
//             mat_A[138] * mat_B[337] +
//             mat_A[139] * mat_B[369] +
//             mat_A[140] * mat_B[401] +
//             mat_A[141] * mat_B[433] +
//             mat_A[142] * mat_B[465] +
//             mat_A[143] * mat_B[497] +
//             mat_A[144] * mat_B[529] +
//             mat_A[145] * mat_B[561] +
//             mat_A[146] * mat_B[593] +
//             mat_A[147] * mat_B[625] +
//             mat_A[148] * mat_B[657] +
//             mat_A[149] * mat_B[689] +
//             mat_A[150] * mat_B[721] +
//             mat_A[151] * mat_B[753] +
//             mat_A[152] * mat_B[785] +
//             mat_A[153] * mat_B[817] +
//             mat_A[154] * mat_B[849] +
//             mat_A[155] * mat_B[881] +
//             mat_A[156] * mat_B[913] +
//             mat_A[157] * mat_B[945] +
//             mat_A[158] * mat_B[977] +
//             mat_A[159] * mat_B[1009];
//  mat_C[146] <= 
//             mat_A[128] * mat_B[18] +
//             mat_A[129] * mat_B[50] +
//             mat_A[130] * mat_B[82] +
//             mat_A[131] * mat_B[114] +
//             mat_A[132] * mat_B[146] +
//             mat_A[133] * mat_B[178] +
//             mat_A[134] * mat_B[210] +
//             mat_A[135] * mat_B[242] +
//             mat_A[136] * mat_B[274] +
//             mat_A[137] * mat_B[306] +
//             mat_A[138] * mat_B[338] +
//             mat_A[139] * mat_B[370] +
//             mat_A[140] * mat_B[402] +
//             mat_A[141] * mat_B[434] +
//             mat_A[142] * mat_B[466] +
//             mat_A[143] * mat_B[498] +
//             mat_A[144] * mat_B[530] +
//             mat_A[145] * mat_B[562] +
//             mat_A[146] * mat_B[594] +
//             mat_A[147] * mat_B[626] +
//             mat_A[148] * mat_B[658] +
//             mat_A[149] * mat_B[690] +
//             mat_A[150] * mat_B[722] +
//             mat_A[151] * mat_B[754] +
//             mat_A[152] * mat_B[786] +
//             mat_A[153] * mat_B[818] +
//             mat_A[154] * mat_B[850] +
//             mat_A[155] * mat_B[882] +
//             mat_A[156] * mat_B[914] +
//             mat_A[157] * mat_B[946] +
//             mat_A[158] * mat_B[978] +
//             mat_A[159] * mat_B[1010];
//  mat_C[147] <= 
//             mat_A[128] * mat_B[19] +
//             mat_A[129] * mat_B[51] +
//             mat_A[130] * mat_B[83] +
//             mat_A[131] * mat_B[115] +
//             mat_A[132] * mat_B[147] +
//             mat_A[133] * mat_B[179] +
//             mat_A[134] * mat_B[211] +
//             mat_A[135] * mat_B[243] +
//             mat_A[136] * mat_B[275] +
//             mat_A[137] * mat_B[307] +
//             mat_A[138] * mat_B[339] +
//             mat_A[139] * mat_B[371] +
//             mat_A[140] * mat_B[403] +
//             mat_A[141] * mat_B[435] +
//             mat_A[142] * mat_B[467] +
//             mat_A[143] * mat_B[499] +
//             mat_A[144] * mat_B[531] +
//             mat_A[145] * mat_B[563] +
//             mat_A[146] * mat_B[595] +
//             mat_A[147] * mat_B[627] +
//             mat_A[148] * mat_B[659] +
//             mat_A[149] * mat_B[691] +
//             mat_A[150] * mat_B[723] +
//             mat_A[151] * mat_B[755] +
//             mat_A[152] * mat_B[787] +
//             mat_A[153] * mat_B[819] +
//             mat_A[154] * mat_B[851] +
//             mat_A[155] * mat_B[883] +
//             mat_A[156] * mat_B[915] +
//             mat_A[157] * mat_B[947] +
//             mat_A[158] * mat_B[979] +
//             mat_A[159] * mat_B[1011];
//  mat_C[148] <= 
//             mat_A[128] * mat_B[20] +
//             mat_A[129] * mat_B[52] +
//             mat_A[130] * mat_B[84] +
//             mat_A[131] * mat_B[116] +
//             mat_A[132] * mat_B[148] +
//             mat_A[133] * mat_B[180] +
//             mat_A[134] * mat_B[212] +
//             mat_A[135] * mat_B[244] +
//             mat_A[136] * mat_B[276] +
//             mat_A[137] * mat_B[308] +
//             mat_A[138] * mat_B[340] +
//             mat_A[139] * mat_B[372] +
//             mat_A[140] * mat_B[404] +
//             mat_A[141] * mat_B[436] +
//             mat_A[142] * mat_B[468] +
//             mat_A[143] * mat_B[500] +
//             mat_A[144] * mat_B[532] +
//             mat_A[145] * mat_B[564] +
//             mat_A[146] * mat_B[596] +
//             mat_A[147] * mat_B[628] +
//             mat_A[148] * mat_B[660] +
//             mat_A[149] * mat_B[692] +
//             mat_A[150] * mat_B[724] +
//             mat_A[151] * mat_B[756] +
//             mat_A[152] * mat_B[788] +
//             mat_A[153] * mat_B[820] +
//             mat_A[154] * mat_B[852] +
//             mat_A[155] * mat_B[884] +
//             mat_A[156] * mat_B[916] +
//             mat_A[157] * mat_B[948] +
//             mat_A[158] * mat_B[980] +
//             mat_A[159] * mat_B[1012];
//  mat_C[149] <= 
//             mat_A[128] * mat_B[21] +
//             mat_A[129] * mat_B[53] +
//             mat_A[130] * mat_B[85] +
//             mat_A[131] * mat_B[117] +
//             mat_A[132] * mat_B[149] +
//             mat_A[133] * mat_B[181] +
//             mat_A[134] * mat_B[213] +
//             mat_A[135] * mat_B[245] +
//             mat_A[136] * mat_B[277] +
//             mat_A[137] * mat_B[309] +
//             mat_A[138] * mat_B[341] +
//             mat_A[139] * mat_B[373] +
//             mat_A[140] * mat_B[405] +
//             mat_A[141] * mat_B[437] +
//             mat_A[142] * mat_B[469] +
//             mat_A[143] * mat_B[501] +
//             mat_A[144] * mat_B[533] +
//             mat_A[145] * mat_B[565] +
//             mat_A[146] * mat_B[597] +
//             mat_A[147] * mat_B[629] +
//             mat_A[148] * mat_B[661] +
//             mat_A[149] * mat_B[693] +
//             mat_A[150] * mat_B[725] +
//             mat_A[151] * mat_B[757] +
//             mat_A[152] * mat_B[789] +
//             mat_A[153] * mat_B[821] +
//             mat_A[154] * mat_B[853] +
//             mat_A[155] * mat_B[885] +
//             mat_A[156] * mat_B[917] +
//             mat_A[157] * mat_B[949] +
//             mat_A[158] * mat_B[981] +
//             mat_A[159] * mat_B[1013];
//  mat_C[150] <= 
//             mat_A[128] * mat_B[22] +
//             mat_A[129] * mat_B[54] +
//             mat_A[130] * mat_B[86] +
//             mat_A[131] * mat_B[118] +
//             mat_A[132] * mat_B[150] +
//             mat_A[133] * mat_B[182] +
//             mat_A[134] * mat_B[214] +
//             mat_A[135] * mat_B[246] +
//             mat_A[136] * mat_B[278] +
//             mat_A[137] * mat_B[310] +
//             mat_A[138] * mat_B[342] +
//             mat_A[139] * mat_B[374] +
//             mat_A[140] * mat_B[406] +
//             mat_A[141] * mat_B[438] +
//             mat_A[142] * mat_B[470] +
//             mat_A[143] * mat_B[502] +
//             mat_A[144] * mat_B[534] +
//             mat_A[145] * mat_B[566] +
//             mat_A[146] * mat_B[598] +
//             mat_A[147] * mat_B[630] +
//             mat_A[148] * mat_B[662] +
//             mat_A[149] * mat_B[694] +
//             mat_A[150] * mat_B[726] +
//             mat_A[151] * mat_B[758] +
//             mat_A[152] * mat_B[790] +
//             mat_A[153] * mat_B[822] +
//             mat_A[154] * mat_B[854] +
//             mat_A[155] * mat_B[886] +
//             mat_A[156] * mat_B[918] +
//             mat_A[157] * mat_B[950] +
//             mat_A[158] * mat_B[982] +
//             mat_A[159] * mat_B[1014];
//  mat_C[151] <= 
//             mat_A[128] * mat_B[23] +
//             mat_A[129] * mat_B[55] +
//             mat_A[130] * mat_B[87] +
//             mat_A[131] * mat_B[119] +
//             mat_A[132] * mat_B[151] +
//             mat_A[133] * mat_B[183] +
//             mat_A[134] * mat_B[215] +
//             mat_A[135] * mat_B[247] +
//             mat_A[136] * mat_B[279] +
//             mat_A[137] * mat_B[311] +
//             mat_A[138] * mat_B[343] +
//             mat_A[139] * mat_B[375] +
//             mat_A[140] * mat_B[407] +
//             mat_A[141] * mat_B[439] +
//             mat_A[142] * mat_B[471] +
//             mat_A[143] * mat_B[503] +
//             mat_A[144] * mat_B[535] +
//             mat_A[145] * mat_B[567] +
//             mat_A[146] * mat_B[599] +
//             mat_A[147] * mat_B[631] +
//             mat_A[148] * mat_B[663] +
//             mat_A[149] * mat_B[695] +
//             mat_A[150] * mat_B[727] +
//             mat_A[151] * mat_B[759] +
//             mat_A[152] * mat_B[791] +
//             mat_A[153] * mat_B[823] +
//             mat_A[154] * mat_B[855] +
//             mat_A[155] * mat_B[887] +
//             mat_A[156] * mat_B[919] +
//             mat_A[157] * mat_B[951] +
//             mat_A[158] * mat_B[983] +
//             mat_A[159] * mat_B[1015];
//  mat_C[152] <= 
//             mat_A[128] * mat_B[24] +
//             mat_A[129] * mat_B[56] +
//             mat_A[130] * mat_B[88] +
//             mat_A[131] * mat_B[120] +
//             mat_A[132] * mat_B[152] +
//             mat_A[133] * mat_B[184] +
//             mat_A[134] * mat_B[216] +
//             mat_A[135] * mat_B[248] +
//             mat_A[136] * mat_B[280] +
//             mat_A[137] * mat_B[312] +
//             mat_A[138] * mat_B[344] +
//             mat_A[139] * mat_B[376] +
//             mat_A[140] * mat_B[408] +
//             mat_A[141] * mat_B[440] +
//             mat_A[142] * mat_B[472] +
//             mat_A[143] * mat_B[504] +
//             mat_A[144] * mat_B[536] +
//             mat_A[145] * mat_B[568] +
//             mat_A[146] * mat_B[600] +
//             mat_A[147] * mat_B[632] +
//             mat_A[148] * mat_B[664] +
//             mat_A[149] * mat_B[696] +
//             mat_A[150] * mat_B[728] +
//             mat_A[151] * mat_B[760] +
//             mat_A[152] * mat_B[792] +
//             mat_A[153] * mat_B[824] +
//             mat_A[154] * mat_B[856] +
//             mat_A[155] * mat_B[888] +
//             mat_A[156] * mat_B[920] +
//             mat_A[157] * mat_B[952] +
//             mat_A[158] * mat_B[984] +
//             mat_A[159] * mat_B[1016];
//  mat_C[153] <= 
//             mat_A[128] * mat_B[25] +
//             mat_A[129] * mat_B[57] +
//             mat_A[130] * mat_B[89] +
//             mat_A[131] * mat_B[121] +
//             mat_A[132] * mat_B[153] +
//             mat_A[133] * mat_B[185] +
//             mat_A[134] * mat_B[217] +
//             mat_A[135] * mat_B[249] +
//             mat_A[136] * mat_B[281] +
//             mat_A[137] * mat_B[313] +
//             mat_A[138] * mat_B[345] +
//             mat_A[139] * mat_B[377] +
//             mat_A[140] * mat_B[409] +
//             mat_A[141] * mat_B[441] +
//             mat_A[142] * mat_B[473] +
//             mat_A[143] * mat_B[505] +
//             mat_A[144] * mat_B[537] +
//             mat_A[145] * mat_B[569] +
//             mat_A[146] * mat_B[601] +
//             mat_A[147] * mat_B[633] +
//             mat_A[148] * mat_B[665] +
//             mat_A[149] * mat_B[697] +
//             mat_A[150] * mat_B[729] +
//             mat_A[151] * mat_B[761] +
//             mat_A[152] * mat_B[793] +
//             mat_A[153] * mat_B[825] +
//             mat_A[154] * mat_B[857] +
//             mat_A[155] * mat_B[889] +
//             mat_A[156] * mat_B[921] +
//             mat_A[157] * mat_B[953] +
//             mat_A[158] * mat_B[985] +
//             mat_A[159] * mat_B[1017];
//  mat_C[154] <= 
//             mat_A[128] * mat_B[26] +
//             mat_A[129] * mat_B[58] +
//             mat_A[130] * mat_B[90] +
//             mat_A[131] * mat_B[122] +
//             mat_A[132] * mat_B[154] +
//             mat_A[133] * mat_B[186] +
//             mat_A[134] * mat_B[218] +
//             mat_A[135] * mat_B[250] +
//             mat_A[136] * mat_B[282] +
//             mat_A[137] * mat_B[314] +
//             mat_A[138] * mat_B[346] +
//             mat_A[139] * mat_B[378] +
//             mat_A[140] * mat_B[410] +
//             mat_A[141] * mat_B[442] +
//             mat_A[142] * mat_B[474] +
//             mat_A[143] * mat_B[506] +
//             mat_A[144] * mat_B[538] +
//             mat_A[145] * mat_B[570] +
//             mat_A[146] * mat_B[602] +
//             mat_A[147] * mat_B[634] +
//             mat_A[148] * mat_B[666] +
//             mat_A[149] * mat_B[698] +
//             mat_A[150] * mat_B[730] +
//             mat_A[151] * mat_B[762] +
//             mat_A[152] * mat_B[794] +
//             mat_A[153] * mat_B[826] +
//             mat_A[154] * mat_B[858] +
//             mat_A[155] * mat_B[890] +
//             mat_A[156] * mat_B[922] +
//             mat_A[157] * mat_B[954] +
//             mat_A[158] * mat_B[986] +
//             mat_A[159] * mat_B[1018];
//  mat_C[155] <= 
//             mat_A[128] * mat_B[27] +
//             mat_A[129] * mat_B[59] +
//             mat_A[130] * mat_B[91] +
//             mat_A[131] * mat_B[123] +
//             mat_A[132] * mat_B[155] +
//             mat_A[133] * mat_B[187] +
//             mat_A[134] * mat_B[219] +
//             mat_A[135] * mat_B[251] +
//             mat_A[136] * mat_B[283] +
//             mat_A[137] * mat_B[315] +
//             mat_A[138] * mat_B[347] +
//             mat_A[139] * mat_B[379] +
//             mat_A[140] * mat_B[411] +
//             mat_A[141] * mat_B[443] +
//             mat_A[142] * mat_B[475] +
//             mat_A[143] * mat_B[507] +
//             mat_A[144] * mat_B[539] +
//             mat_A[145] * mat_B[571] +
//             mat_A[146] * mat_B[603] +
//             mat_A[147] * mat_B[635] +
//             mat_A[148] * mat_B[667] +
//             mat_A[149] * mat_B[699] +
//             mat_A[150] * mat_B[731] +
//             mat_A[151] * mat_B[763] +
//             mat_A[152] * mat_B[795] +
//             mat_A[153] * mat_B[827] +
//             mat_A[154] * mat_B[859] +
//             mat_A[155] * mat_B[891] +
//             mat_A[156] * mat_B[923] +
//             mat_A[157] * mat_B[955] +
//             mat_A[158] * mat_B[987] +
//             mat_A[159] * mat_B[1019];
//  mat_C[156] <= 
//             mat_A[128] * mat_B[28] +
//             mat_A[129] * mat_B[60] +
//             mat_A[130] * mat_B[92] +
//             mat_A[131] * mat_B[124] +
//             mat_A[132] * mat_B[156] +
//             mat_A[133] * mat_B[188] +
//             mat_A[134] * mat_B[220] +
//             mat_A[135] * mat_B[252] +
//             mat_A[136] * mat_B[284] +
//             mat_A[137] * mat_B[316] +
//             mat_A[138] * mat_B[348] +
//             mat_A[139] * mat_B[380] +
//             mat_A[140] * mat_B[412] +
//             mat_A[141] * mat_B[444] +
//             mat_A[142] * mat_B[476] +
//             mat_A[143] * mat_B[508] +
//             mat_A[144] * mat_B[540] +
//             mat_A[145] * mat_B[572] +
//             mat_A[146] * mat_B[604] +
//             mat_A[147] * mat_B[636] +
//             mat_A[148] * mat_B[668] +
//             mat_A[149] * mat_B[700] +
//             mat_A[150] * mat_B[732] +
//             mat_A[151] * mat_B[764] +
//             mat_A[152] * mat_B[796] +
//             mat_A[153] * mat_B[828] +
//             mat_A[154] * mat_B[860] +
//             mat_A[155] * mat_B[892] +
//             mat_A[156] * mat_B[924] +
//             mat_A[157] * mat_B[956] +
//             mat_A[158] * mat_B[988] +
//             mat_A[159] * mat_B[1020];
//  mat_C[157] <= 
//             mat_A[128] * mat_B[29] +
//             mat_A[129] * mat_B[61] +
//             mat_A[130] * mat_B[93] +
//             mat_A[131] * mat_B[125] +
//             mat_A[132] * mat_B[157] +
//             mat_A[133] * mat_B[189] +
//             mat_A[134] * mat_B[221] +
//             mat_A[135] * mat_B[253] +
//             mat_A[136] * mat_B[285] +
//             mat_A[137] * mat_B[317] +
//             mat_A[138] * mat_B[349] +
//             mat_A[139] * mat_B[381] +
//             mat_A[140] * mat_B[413] +
//             mat_A[141] * mat_B[445] +
//             mat_A[142] * mat_B[477] +
//             mat_A[143] * mat_B[509] +
//             mat_A[144] * mat_B[541] +
//             mat_A[145] * mat_B[573] +
//             mat_A[146] * mat_B[605] +
//             mat_A[147] * mat_B[637] +
//             mat_A[148] * mat_B[669] +
//             mat_A[149] * mat_B[701] +
//             mat_A[150] * mat_B[733] +
//             mat_A[151] * mat_B[765] +
//             mat_A[152] * mat_B[797] +
//             mat_A[153] * mat_B[829] +
//             mat_A[154] * mat_B[861] +
//             mat_A[155] * mat_B[893] +
//             mat_A[156] * mat_B[925] +
//             mat_A[157] * mat_B[957] +
//             mat_A[158] * mat_B[989] +
//             mat_A[159] * mat_B[1021];
//  mat_C[158] <= 
//             mat_A[128] * mat_B[30] +
//             mat_A[129] * mat_B[62] +
//             mat_A[130] * mat_B[94] +
//             mat_A[131] * mat_B[126] +
//             mat_A[132] * mat_B[158] +
//             mat_A[133] * mat_B[190] +
//             mat_A[134] * mat_B[222] +
//             mat_A[135] * mat_B[254] +
//             mat_A[136] * mat_B[286] +
//             mat_A[137] * mat_B[318] +
//             mat_A[138] * mat_B[350] +
//             mat_A[139] * mat_B[382] +
//             mat_A[140] * mat_B[414] +
//             mat_A[141] * mat_B[446] +
//             mat_A[142] * mat_B[478] +
//             mat_A[143] * mat_B[510] +
//             mat_A[144] * mat_B[542] +
//             mat_A[145] * mat_B[574] +
//             mat_A[146] * mat_B[606] +
//             mat_A[147] * mat_B[638] +
//             mat_A[148] * mat_B[670] +
//             mat_A[149] * mat_B[702] +
//             mat_A[150] * mat_B[734] +
//             mat_A[151] * mat_B[766] +
//             mat_A[152] * mat_B[798] +
//             mat_A[153] * mat_B[830] +
//             mat_A[154] * mat_B[862] +
//             mat_A[155] * mat_B[894] +
//             mat_A[156] * mat_B[926] +
//             mat_A[157] * mat_B[958] +
//             mat_A[158] * mat_B[990] +
//             mat_A[159] * mat_B[1022];
//  mat_C[159] <= 
//             mat_A[128] * mat_B[31] +
//             mat_A[129] * mat_B[63] +
//             mat_A[130] * mat_B[95] +
//             mat_A[131] * mat_B[127] +
//             mat_A[132] * mat_B[159] +
//             mat_A[133] * mat_B[191] +
//             mat_A[134] * mat_B[223] +
//             mat_A[135] * mat_B[255] +
//             mat_A[136] * mat_B[287] +
//             mat_A[137] * mat_B[319] +
//             mat_A[138] * mat_B[351] +
//             mat_A[139] * mat_B[383] +
//             mat_A[140] * mat_B[415] +
//             mat_A[141] * mat_B[447] +
//             mat_A[142] * mat_B[479] +
//             mat_A[143] * mat_B[511] +
//             mat_A[144] * mat_B[543] +
//             mat_A[145] * mat_B[575] +
//             mat_A[146] * mat_B[607] +
//             mat_A[147] * mat_B[639] +
//             mat_A[148] * mat_B[671] +
//             mat_A[149] * mat_B[703] +
//             mat_A[150] * mat_B[735] +
//             mat_A[151] * mat_B[767] +
//             mat_A[152] * mat_B[799] +
//             mat_A[153] * mat_B[831] +
//             mat_A[154] * mat_B[863] +
//             mat_A[155] * mat_B[895] +
//             mat_A[156] * mat_B[927] +
//             mat_A[157] * mat_B[959] +
//             mat_A[158] * mat_B[991] +
//             mat_A[159] * mat_B[1023];
//  mat_C[160] <= 
//             mat_A[160] * mat_B[0] +
//             mat_A[161] * mat_B[32] +
//             mat_A[162] * mat_B[64] +
//             mat_A[163] * mat_B[96] +
//             mat_A[164] * mat_B[128] +
//             mat_A[165] * mat_B[160] +
//             mat_A[166] * mat_B[192] +
//             mat_A[167] * mat_B[224] +
//             mat_A[168] * mat_B[256] +
//             mat_A[169] * mat_B[288] +
//             mat_A[170] * mat_B[320] +
//             mat_A[171] * mat_B[352] +
//             mat_A[172] * mat_B[384] +
//             mat_A[173] * mat_B[416] +
//             mat_A[174] * mat_B[448] +
//             mat_A[175] * mat_B[480] +
//             mat_A[176] * mat_B[512] +
//             mat_A[177] * mat_B[544] +
//             mat_A[178] * mat_B[576] +
//             mat_A[179] * mat_B[608] +
//             mat_A[180] * mat_B[640] +
//             mat_A[181] * mat_B[672] +
//             mat_A[182] * mat_B[704] +
//             mat_A[183] * mat_B[736] +
//             mat_A[184] * mat_B[768] +
//             mat_A[185] * mat_B[800] +
//             mat_A[186] * mat_B[832] +
//             mat_A[187] * mat_B[864] +
//             mat_A[188] * mat_B[896] +
//             mat_A[189] * mat_B[928] +
//             mat_A[190] * mat_B[960] +
//             mat_A[191] * mat_B[992];
//  mat_C[161] <= 
//             mat_A[160] * mat_B[1] +
//             mat_A[161] * mat_B[33] +
//             mat_A[162] * mat_B[65] +
//             mat_A[163] * mat_B[97] +
//             mat_A[164] * mat_B[129] +
//             mat_A[165] * mat_B[161] +
//             mat_A[166] * mat_B[193] +
//             mat_A[167] * mat_B[225] +
//             mat_A[168] * mat_B[257] +
//             mat_A[169] * mat_B[289] +
//             mat_A[170] * mat_B[321] +
//             mat_A[171] * mat_B[353] +
//             mat_A[172] * mat_B[385] +
//             mat_A[173] * mat_B[417] +
//             mat_A[174] * mat_B[449] +
//             mat_A[175] * mat_B[481] +
//             mat_A[176] * mat_B[513] +
//             mat_A[177] * mat_B[545] +
//             mat_A[178] * mat_B[577] +
//             mat_A[179] * mat_B[609] +
//             mat_A[180] * mat_B[641] +
//             mat_A[181] * mat_B[673] +
//             mat_A[182] * mat_B[705] +
//             mat_A[183] * mat_B[737] +
//             mat_A[184] * mat_B[769] +
//             mat_A[185] * mat_B[801] +
//             mat_A[186] * mat_B[833] +
//             mat_A[187] * mat_B[865] +
//             mat_A[188] * mat_B[897] +
//             mat_A[189] * mat_B[929] +
//             mat_A[190] * mat_B[961] +
//             mat_A[191] * mat_B[993];
//  mat_C[162] <= 
//             mat_A[160] * mat_B[2] +
//             mat_A[161] * mat_B[34] +
//             mat_A[162] * mat_B[66] +
//             mat_A[163] * mat_B[98] +
//             mat_A[164] * mat_B[130] +
//             mat_A[165] * mat_B[162] +
//             mat_A[166] * mat_B[194] +
//             mat_A[167] * mat_B[226] +
//             mat_A[168] * mat_B[258] +
//             mat_A[169] * mat_B[290] +
//             mat_A[170] * mat_B[322] +
//             mat_A[171] * mat_B[354] +
//             mat_A[172] * mat_B[386] +
//             mat_A[173] * mat_B[418] +
//             mat_A[174] * mat_B[450] +
//             mat_A[175] * mat_B[482] +
//             mat_A[176] * mat_B[514] +
//             mat_A[177] * mat_B[546] +
//             mat_A[178] * mat_B[578] +
//             mat_A[179] * mat_B[610] +
//             mat_A[180] * mat_B[642] +
//             mat_A[181] * mat_B[674] +
//             mat_A[182] * mat_B[706] +
//             mat_A[183] * mat_B[738] +
//             mat_A[184] * mat_B[770] +
//             mat_A[185] * mat_B[802] +
//             mat_A[186] * mat_B[834] +
//             mat_A[187] * mat_B[866] +
//             mat_A[188] * mat_B[898] +
//             mat_A[189] * mat_B[930] +
//             mat_A[190] * mat_B[962] +
//             mat_A[191] * mat_B[994];
//  mat_C[163] <= 
//             mat_A[160] * mat_B[3] +
//             mat_A[161] * mat_B[35] +
//             mat_A[162] * mat_B[67] +
//             mat_A[163] * mat_B[99] +
//             mat_A[164] * mat_B[131] +
//             mat_A[165] * mat_B[163] +
//             mat_A[166] * mat_B[195] +
//             mat_A[167] * mat_B[227] +
//             mat_A[168] * mat_B[259] +
//             mat_A[169] * mat_B[291] +
//             mat_A[170] * mat_B[323] +
//             mat_A[171] * mat_B[355] +
//             mat_A[172] * mat_B[387] +
//             mat_A[173] * mat_B[419] +
//             mat_A[174] * mat_B[451] +
//             mat_A[175] * mat_B[483] +
//             mat_A[176] * mat_B[515] +
//             mat_A[177] * mat_B[547] +
//             mat_A[178] * mat_B[579] +
//             mat_A[179] * mat_B[611] +
//             mat_A[180] * mat_B[643] +
//             mat_A[181] * mat_B[675] +
//             mat_A[182] * mat_B[707] +
//             mat_A[183] * mat_B[739] +
//             mat_A[184] * mat_B[771] +
//             mat_A[185] * mat_B[803] +
//             mat_A[186] * mat_B[835] +
//             mat_A[187] * mat_B[867] +
//             mat_A[188] * mat_B[899] +
//             mat_A[189] * mat_B[931] +
//             mat_A[190] * mat_B[963] +
//             mat_A[191] * mat_B[995];
//  mat_C[164] <= 
//             mat_A[160] * mat_B[4] +
//             mat_A[161] * mat_B[36] +
//             mat_A[162] * mat_B[68] +
//             mat_A[163] * mat_B[100] +
//             mat_A[164] * mat_B[132] +
//             mat_A[165] * mat_B[164] +
//             mat_A[166] * mat_B[196] +
//             mat_A[167] * mat_B[228] +
//             mat_A[168] * mat_B[260] +
//             mat_A[169] * mat_B[292] +
//             mat_A[170] * mat_B[324] +
//             mat_A[171] * mat_B[356] +
//             mat_A[172] * mat_B[388] +
//             mat_A[173] * mat_B[420] +
//             mat_A[174] * mat_B[452] +
//             mat_A[175] * mat_B[484] +
//             mat_A[176] * mat_B[516] +
//             mat_A[177] * mat_B[548] +
//             mat_A[178] * mat_B[580] +
//             mat_A[179] * mat_B[612] +
//             mat_A[180] * mat_B[644] +
//             mat_A[181] * mat_B[676] +
//             mat_A[182] * mat_B[708] +
//             mat_A[183] * mat_B[740] +
//             mat_A[184] * mat_B[772] +
//             mat_A[185] * mat_B[804] +
//             mat_A[186] * mat_B[836] +
//             mat_A[187] * mat_B[868] +
//             mat_A[188] * mat_B[900] +
//             mat_A[189] * mat_B[932] +
//             mat_A[190] * mat_B[964] +
//             mat_A[191] * mat_B[996];
//  mat_C[165] <= 
//             mat_A[160] * mat_B[5] +
//             mat_A[161] * mat_B[37] +
//             mat_A[162] * mat_B[69] +
//             mat_A[163] * mat_B[101] +
//             mat_A[164] * mat_B[133] +
//             mat_A[165] * mat_B[165] +
//             mat_A[166] * mat_B[197] +
//             mat_A[167] * mat_B[229] +
//             mat_A[168] * mat_B[261] +
//             mat_A[169] * mat_B[293] +
//             mat_A[170] * mat_B[325] +
//             mat_A[171] * mat_B[357] +
//             mat_A[172] * mat_B[389] +
//             mat_A[173] * mat_B[421] +
//             mat_A[174] * mat_B[453] +
//             mat_A[175] * mat_B[485] +
//             mat_A[176] * mat_B[517] +
//             mat_A[177] * mat_B[549] +
//             mat_A[178] * mat_B[581] +
//             mat_A[179] * mat_B[613] +
//             mat_A[180] * mat_B[645] +
//             mat_A[181] * mat_B[677] +
//             mat_A[182] * mat_B[709] +
//             mat_A[183] * mat_B[741] +
//             mat_A[184] * mat_B[773] +
//             mat_A[185] * mat_B[805] +
//             mat_A[186] * mat_B[837] +
//             mat_A[187] * mat_B[869] +
//             mat_A[188] * mat_B[901] +
//             mat_A[189] * mat_B[933] +
//             mat_A[190] * mat_B[965] +
//             mat_A[191] * mat_B[997];
//  mat_C[166] <= 
//             mat_A[160] * mat_B[6] +
//             mat_A[161] * mat_B[38] +
//             mat_A[162] * mat_B[70] +
//             mat_A[163] * mat_B[102] +
//             mat_A[164] * mat_B[134] +
//             mat_A[165] * mat_B[166] +
//             mat_A[166] * mat_B[198] +
//             mat_A[167] * mat_B[230] +
//             mat_A[168] * mat_B[262] +
//             mat_A[169] * mat_B[294] +
//             mat_A[170] * mat_B[326] +
//             mat_A[171] * mat_B[358] +
//             mat_A[172] * mat_B[390] +
//             mat_A[173] * mat_B[422] +
//             mat_A[174] * mat_B[454] +
//             mat_A[175] * mat_B[486] +
//             mat_A[176] * mat_B[518] +
//             mat_A[177] * mat_B[550] +
//             mat_A[178] * mat_B[582] +
//             mat_A[179] * mat_B[614] +
//             mat_A[180] * mat_B[646] +
//             mat_A[181] * mat_B[678] +
//             mat_A[182] * mat_B[710] +
//             mat_A[183] * mat_B[742] +
//             mat_A[184] * mat_B[774] +
//             mat_A[185] * mat_B[806] +
//             mat_A[186] * mat_B[838] +
//             mat_A[187] * mat_B[870] +
//             mat_A[188] * mat_B[902] +
//             mat_A[189] * mat_B[934] +
//             mat_A[190] * mat_B[966] +
//             mat_A[191] * mat_B[998];
//  mat_C[167] <= 
//             mat_A[160] * mat_B[7] +
//             mat_A[161] * mat_B[39] +
//             mat_A[162] * mat_B[71] +
//             mat_A[163] * mat_B[103] +
//             mat_A[164] * mat_B[135] +
//             mat_A[165] * mat_B[167] +
//             mat_A[166] * mat_B[199] +
//             mat_A[167] * mat_B[231] +
//             mat_A[168] * mat_B[263] +
//             mat_A[169] * mat_B[295] +
//             mat_A[170] * mat_B[327] +
//             mat_A[171] * mat_B[359] +
//             mat_A[172] * mat_B[391] +
//             mat_A[173] * mat_B[423] +
//             mat_A[174] * mat_B[455] +
//             mat_A[175] * mat_B[487] +
//             mat_A[176] * mat_B[519] +
//             mat_A[177] * mat_B[551] +
//             mat_A[178] * mat_B[583] +
//             mat_A[179] * mat_B[615] +
//             mat_A[180] * mat_B[647] +
//             mat_A[181] * mat_B[679] +
//             mat_A[182] * mat_B[711] +
//             mat_A[183] * mat_B[743] +
//             mat_A[184] * mat_B[775] +
//             mat_A[185] * mat_B[807] +
//             mat_A[186] * mat_B[839] +
//             mat_A[187] * mat_B[871] +
//             mat_A[188] * mat_B[903] +
//             mat_A[189] * mat_B[935] +
//             mat_A[190] * mat_B[967] +
//             mat_A[191] * mat_B[999];
//  mat_C[168] <= 
//             mat_A[160] * mat_B[8] +
//             mat_A[161] * mat_B[40] +
//             mat_A[162] * mat_B[72] +
//             mat_A[163] * mat_B[104] +
//             mat_A[164] * mat_B[136] +
//             mat_A[165] * mat_B[168] +
//             mat_A[166] * mat_B[200] +
//             mat_A[167] * mat_B[232] +
//             mat_A[168] * mat_B[264] +
//             mat_A[169] * mat_B[296] +
//             mat_A[170] * mat_B[328] +
//             mat_A[171] * mat_B[360] +
//             mat_A[172] * mat_B[392] +
//             mat_A[173] * mat_B[424] +
//             mat_A[174] * mat_B[456] +
//             mat_A[175] * mat_B[488] +
//             mat_A[176] * mat_B[520] +
//             mat_A[177] * mat_B[552] +
//             mat_A[178] * mat_B[584] +
//             mat_A[179] * mat_B[616] +
//             mat_A[180] * mat_B[648] +
//             mat_A[181] * mat_B[680] +
//             mat_A[182] * mat_B[712] +
//             mat_A[183] * mat_B[744] +
//             mat_A[184] * mat_B[776] +
//             mat_A[185] * mat_B[808] +
//             mat_A[186] * mat_B[840] +
//             mat_A[187] * mat_B[872] +
//             mat_A[188] * mat_B[904] +
//             mat_A[189] * mat_B[936] +
//             mat_A[190] * mat_B[968] +
//             mat_A[191] * mat_B[1000];
//  mat_C[169] <= 
//             mat_A[160] * mat_B[9] +
//             mat_A[161] * mat_B[41] +
//             mat_A[162] * mat_B[73] +
//             mat_A[163] * mat_B[105] +
//             mat_A[164] * mat_B[137] +
//             mat_A[165] * mat_B[169] +
//             mat_A[166] * mat_B[201] +
//             mat_A[167] * mat_B[233] +
//             mat_A[168] * mat_B[265] +
//             mat_A[169] * mat_B[297] +
//             mat_A[170] * mat_B[329] +
//             mat_A[171] * mat_B[361] +
//             mat_A[172] * mat_B[393] +
//             mat_A[173] * mat_B[425] +
//             mat_A[174] * mat_B[457] +
//             mat_A[175] * mat_B[489] +
//             mat_A[176] * mat_B[521] +
//             mat_A[177] * mat_B[553] +
//             mat_A[178] * mat_B[585] +
//             mat_A[179] * mat_B[617] +
//             mat_A[180] * mat_B[649] +
//             mat_A[181] * mat_B[681] +
//             mat_A[182] * mat_B[713] +
//             mat_A[183] * mat_B[745] +
//             mat_A[184] * mat_B[777] +
//             mat_A[185] * mat_B[809] +
//             mat_A[186] * mat_B[841] +
//             mat_A[187] * mat_B[873] +
//             mat_A[188] * mat_B[905] +
//             mat_A[189] * mat_B[937] +
//             mat_A[190] * mat_B[969] +
//             mat_A[191] * mat_B[1001];
//  mat_C[170] <= 
//             mat_A[160] * mat_B[10] +
//             mat_A[161] * mat_B[42] +
//             mat_A[162] * mat_B[74] +
//             mat_A[163] * mat_B[106] +
//             mat_A[164] * mat_B[138] +
//             mat_A[165] * mat_B[170] +
//             mat_A[166] * mat_B[202] +
//             mat_A[167] * mat_B[234] +
//             mat_A[168] * mat_B[266] +
//             mat_A[169] * mat_B[298] +
//             mat_A[170] * mat_B[330] +
//             mat_A[171] * mat_B[362] +
//             mat_A[172] * mat_B[394] +
//             mat_A[173] * mat_B[426] +
//             mat_A[174] * mat_B[458] +
//             mat_A[175] * mat_B[490] +
//             mat_A[176] * mat_B[522] +
//             mat_A[177] * mat_B[554] +
//             mat_A[178] * mat_B[586] +
//             mat_A[179] * mat_B[618] +
//             mat_A[180] * mat_B[650] +
//             mat_A[181] * mat_B[682] +
//             mat_A[182] * mat_B[714] +
//             mat_A[183] * mat_B[746] +
//             mat_A[184] * mat_B[778] +
//             mat_A[185] * mat_B[810] +
//             mat_A[186] * mat_B[842] +
//             mat_A[187] * mat_B[874] +
//             mat_A[188] * mat_B[906] +
//             mat_A[189] * mat_B[938] +
//             mat_A[190] * mat_B[970] +
//             mat_A[191] * mat_B[1002];
//  mat_C[171] <= 
//             mat_A[160] * mat_B[11] +
//             mat_A[161] * mat_B[43] +
//             mat_A[162] * mat_B[75] +
//             mat_A[163] * mat_B[107] +
//             mat_A[164] * mat_B[139] +
//             mat_A[165] * mat_B[171] +
//             mat_A[166] * mat_B[203] +
//             mat_A[167] * mat_B[235] +
//             mat_A[168] * mat_B[267] +
//             mat_A[169] * mat_B[299] +
//             mat_A[170] * mat_B[331] +
//             mat_A[171] * mat_B[363] +
//             mat_A[172] * mat_B[395] +
//             mat_A[173] * mat_B[427] +
//             mat_A[174] * mat_B[459] +
//             mat_A[175] * mat_B[491] +
//             mat_A[176] * mat_B[523] +
//             mat_A[177] * mat_B[555] +
//             mat_A[178] * mat_B[587] +
//             mat_A[179] * mat_B[619] +
//             mat_A[180] * mat_B[651] +
//             mat_A[181] * mat_B[683] +
//             mat_A[182] * mat_B[715] +
//             mat_A[183] * mat_B[747] +
//             mat_A[184] * mat_B[779] +
//             mat_A[185] * mat_B[811] +
//             mat_A[186] * mat_B[843] +
//             mat_A[187] * mat_B[875] +
//             mat_A[188] * mat_B[907] +
//             mat_A[189] * mat_B[939] +
//             mat_A[190] * mat_B[971] +
//             mat_A[191] * mat_B[1003];
//  mat_C[172] <= 
//             mat_A[160] * mat_B[12] +
//             mat_A[161] * mat_B[44] +
//             mat_A[162] * mat_B[76] +
//             mat_A[163] * mat_B[108] +
//             mat_A[164] * mat_B[140] +
//             mat_A[165] * mat_B[172] +
//             mat_A[166] * mat_B[204] +
//             mat_A[167] * mat_B[236] +
//             mat_A[168] * mat_B[268] +
//             mat_A[169] * mat_B[300] +
//             mat_A[170] * mat_B[332] +
//             mat_A[171] * mat_B[364] +
//             mat_A[172] * mat_B[396] +
//             mat_A[173] * mat_B[428] +
//             mat_A[174] * mat_B[460] +
//             mat_A[175] * mat_B[492] +
//             mat_A[176] * mat_B[524] +
//             mat_A[177] * mat_B[556] +
//             mat_A[178] * mat_B[588] +
//             mat_A[179] * mat_B[620] +
//             mat_A[180] * mat_B[652] +
//             mat_A[181] * mat_B[684] +
//             mat_A[182] * mat_B[716] +
//             mat_A[183] * mat_B[748] +
//             mat_A[184] * mat_B[780] +
//             mat_A[185] * mat_B[812] +
//             mat_A[186] * mat_B[844] +
//             mat_A[187] * mat_B[876] +
//             mat_A[188] * mat_B[908] +
//             mat_A[189] * mat_B[940] +
//             mat_A[190] * mat_B[972] +
//             mat_A[191] * mat_B[1004];
//  mat_C[173] <= 
//             mat_A[160] * mat_B[13] +
//             mat_A[161] * mat_B[45] +
//             mat_A[162] * mat_B[77] +
//             mat_A[163] * mat_B[109] +
//             mat_A[164] * mat_B[141] +
//             mat_A[165] * mat_B[173] +
//             mat_A[166] * mat_B[205] +
//             mat_A[167] * mat_B[237] +
//             mat_A[168] * mat_B[269] +
//             mat_A[169] * mat_B[301] +
//             mat_A[170] * mat_B[333] +
//             mat_A[171] * mat_B[365] +
//             mat_A[172] * mat_B[397] +
//             mat_A[173] * mat_B[429] +
//             mat_A[174] * mat_B[461] +
//             mat_A[175] * mat_B[493] +
//             mat_A[176] * mat_B[525] +
//             mat_A[177] * mat_B[557] +
//             mat_A[178] * mat_B[589] +
//             mat_A[179] * mat_B[621] +
//             mat_A[180] * mat_B[653] +
//             mat_A[181] * mat_B[685] +
//             mat_A[182] * mat_B[717] +
//             mat_A[183] * mat_B[749] +
//             mat_A[184] * mat_B[781] +
//             mat_A[185] * mat_B[813] +
//             mat_A[186] * mat_B[845] +
//             mat_A[187] * mat_B[877] +
//             mat_A[188] * mat_B[909] +
//             mat_A[189] * mat_B[941] +
//             mat_A[190] * mat_B[973] +
//             mat_A[191] * mat_B[1005];
//  mat_C[174] <= 
//             mat_A[160] * mat_B[14] +
//             mat_A[161] * mat_B[46] +
//             mat_A[162] * mat_B[78] +
//             mat_A[163] * mat_B[110] +
//             mat_A[164] * mat_B[142] +
//             mat_A[165] * mat_B[174] +
//             mat_A[166] * mat_B[206] +
//             mat_A[167] * mat_B[238] +
//             mat_A[168] * mat_B[270] +
//             mat_A[169] * mat_B[302] +
//             mat_A[170] * mat_B[334] +
//             mat_A[171] * mat_B[366] +
//             mat_A[172] * mat_B[398] +
//             mat_A[173] * mat_B[430] +
//             mat_A[174] * mat_B[462] +
//             mat_A[175] * mat_B[494] +
//             mat_A[176] * mat_B[526] +
//             mat_A[177] * mat_B[558] +
//             mat_A[178] * mat_B[590] +
//             mat_A[179] * mat_B[622] +
//             mat_A[180] * mat_B[654] +
//             mat_A[181] * mat_B[686] +
//             mat_A[182] * mat_B[718] +
//             mat_A[183] * mat_B[750] +
//             mat_A[184] * mat_B[782] +
//             mat_A[185] * mat_B[814] +
//             mat_A[186] * mat_B[846] +
//             mat_A[187] * mat_B[878] +
//             mat_A[188] * mat_B[910] +
//             mat_A[189] * mat_B[942] +
//             mat_A[190] * mat_B[974] +
//             mat_A[191] * mat_B[1006];
//  mat_C[175] <= 
//             mat_A[160] * mat_B[15] +
//             mat_A[161] * mat_B[47] +
//             mat_A[162] * mat_B[79] +
//             mat_A[163] * mat_B[111] +
//             mat_A[164] * mat_B[143] +
//             mat_A[165] * mat_B[175] +
//             mat_A[166] * mat_B[207] +
//             mat_A[167] * mat_B[239] +
//             mat_A[168] * mat_B[271] +
//             mat_A[169] * mat_B[303] +
//             mat_A[170] * mat_B[335] +
//             mat_A[171] * mat_B[367] +
//             mat_A[172] * mat_B[399] +
//             mat_A[173] * mat_B[431] +
//             mat_A[174] * mat_B[463] +
//             mat_A[175] * mat_B[495] +
//             mat_A[176] * mat_B[527] +
//             mat_A[177] * mat_B[559] +
//             mat_A[178] * mat_B[591] +
//             mat_A[179] * mat_B[623] +
//             mat_A[180] * mat_B[655] +
//             mat_A[181] * mat_B[687] +
//             mat_A[182] * mat_B[719] +
//             mat_A[183] * mat_B[751] +
//             mat_A[184] * mat_B[783] +
//             mat_A[185] * mat_B[815] +
//             mat_A[186] * mat_B[847] +
//             mat_A[187] * mat_B[879] +
//             mat_A[188] * mat_B[911] +
//             mat_A[189] * mat_B[943] +
//             mat_A[190] * mat_B[975] +
//             mat_A[191] * mat_B[1007];
//  mat_C[176] <= 
//             mat_A[160] * mat_B[16] +
//             mat_A[161] * mat_B[48] +
//             mat_A[162] * mat_B[80] +
//             mat_A[163] * mat_B[112] +
//             mat_A[164] * mat_B[144] +
//             mat_A[165] * mat_B[176] +
//             mat_A[166] * mat_B[208] +
//             mat_A[167] * mat_B[240] +
//             mat_A[168] * mat_B[272] +
//             mat_A[169] * mat_B[304] +
//             mat_A[170] * mat_B[336] +
//             mat_A[171] * mat_B[368] +
//             mat_A[172] * mat_B[400] +
//             mat_A[173] * mat_B[432] +
//             mat_A[174] * mat_B[464] +
//             mat_A[175] * mat_B[496] +
//             mat_A[176] * mat_B[528] +
//             mat_A[177] * mat_B[560] +
//             mat_A[178] * mat_B[592] +
//             mat_A[179] * mat_B[624] +
//             mat_A[180] * mat_B[656] +
//             mat_A[181] * mat_B[688] +
//             mat_A[182] * mat_B[720] +
//             mat_A[183] * mat_B[752] +
//             mat_A[184] * mat_B[784] +
//             mat_A[185] * mat_B[816] +
//             mat_A[186] * mat_B[848] +
//             mat_A[187] * mat_B[880] +
//             mat_A[188] * mat_B[912] +
//             mat_A[189] * mat_B[944] +
//             mat_A[190] * mat_B[976] +
//             mat_A[191] * mat_B[1008];
//  mat_C[177] <= 
//             mat_A[160] * mat_B[17] +
//             mat_A[161] * mat_B[49] +
//             mat_A[162] * mat_B[81] +
//             mat_A[163] * mat_B[113] +
//             mat_A[164] * mat_B[145] +
//             mat_A[165] * mat_B[177] +
//             mat_A[166] * mat_B[209] +
//             mat_A[167] * mat_B[241] +
//             mat_A[168] * mat_B[273] +
//             mat_A[169] * mat_B[305] +
//             mat_A[170] * mat_B[337] +
//             mat_A[171] * mat_B[369] +
//             mat_A[172] * mat_B[401] +
//             mat_A[173] * mat_B[433] +
//             mat_A[174] * mat_B[465] +
//             mat_A[175] * mat_B[497] +
//             mat_A[176] * mat_B[529] +
//             mat_A[177] * mat_B[561] +
//             mat_A[178] * mat_B[593] +
//             mat_A[179] * mat_B[625] +
//             mat_A[180] * mat_B[657] +
//             mat_A[181] * mat_B[689] +
//             mat_A[182] * mat_B[721] +
//             mat_A[183] * mat_B[753] +
//             mat_A[184] * mat_B[785] +
//             mat_A[185] * mat_B[817] +
//             mat_A[186] * mat_B[849] +
//             mat_A[187] * mat_B[881] +
//             mat_A[188] * mat_B[913] +
//             mat_A[189] * mat_B[945] +
//             mat_A[190] * mat_B[977] +
//             mat_A[191] * mat_B[1009];
//  mat_C[178] <= 
//             mat_A[160] * mat_B[18] +
//             mat_A[161] * mat_B[50] +
//             mat_A[162] * mat_B[82] +
//             mat_A[163] * mat_B[114] +
//             mat_A[164] * mat_B[146] +
//             mat_A[165] * mat_B[178] +
//             mat_A[166] * mat_B[210] +
//             mat_A[167] * mat_B[242] +
//             mat_A[168] * mat_B[274] +
//             mat_A[169] * mat_B[306] +
//             mat_A[170] * mat_B[338] +
//             mat_A[171] * mat_B[370] +
//             mat_A[172] * mat_B[402] +
//             mat_A[173] * mat_B[434] +
//             mat_A[174] * mat_B[466] +
//             mat_A[175] * mat_B[498] +
//             mat_A[176] * mat_B[530] +
//             mat_A[177] * mat_B[562] +
//             mat_A[178] * mat_B[594] +
//             mat_A[179] * mat_B[626] +
//             mat_A[180] * mat_B[658] +
//             mat_A[181] * mat_B[690] +
//             mat_A[182] * mat_B[722] +
//             mat_A[183] * mat_B[754] +
//             mat_A[184] * mat_B[786] +
//             mat_A[185] * mat_B[818] +
//             mat_A[186] * mat_B[850] +
//             mat_A[187] * mat_B[882] +
//             mat_A[188] * mat_B[914] +
//             mat_A[189] * mat_B[946] +
//             mat_A[190] * mat_B[978] +
//             mat_A[191] * mat_B[1010];
//  mat_C[179] <= 
//             mat_A[160] * mat_B[19] +
//             mat_A[161] * mat_B[51] +
//             mat_A[162] * mat_B[83] +
//             mat_A[163] * mat_B[115] +
//             mat_A[164] * mat_B[147] +
//             mat_A[165] * mat_B[179] +
//             mat_A[166] * mat_B[211] +
//             mat_A[167] * mat_B[243] +
//             mat_A[168] * mat_B[275] +
//             mat_A[169] * mat_B[307] +
//             mat_A[170] * mat_B[339] +
//             mat_A[171] * mat_B[371] +
//             mat_A[172] * mat_B[403] +
//             mat_A[173] * mat_B[435] +
//             mat_A[174] * mat_B[467] +
//             mat_A[175] * mat_B[499] +
//             mat_A[176] * mat_B[531] +
//             mat_A[177] * mat_B[563] +
//             mat_A[178] * mat_B[595] +
//             mat_A[179] * mat_B[627] +
//             mat_A[180] * mat_B[659] +
//             mat_A[181] * mat_B[691] +
//             mat_A[182] * mat_B[723] +
//             mat_A[183] * mat_B[755] +
//             mat_A[184] * mat_B[787] +
//             mat_A[185] * mat_B[819] +
//             mat_A[186] * mat_B[851] +
//             mat_A[187] * mat_B[883] +
//             mat_A[188] * mat_B[915] +
//             mat_A[189] * mat_B[947] +
//             mat_A[190] * mat_B[979] +
//             mat_A[191] * mat_B[1011];
//  mat_C[180] <= 
//             mat_A[160] * mat_B[20] +
//             mat_A[161] * mat_B[52] +
//             mat_A[162] * mat_B[84] +
//             mat_A[163] * mat_B[116] +
//             mat_A[164] * mat_B[148] +
//             mat_A[165] * mat_B[180] +
//             mat_A[166] * mat_B[212] +
//             mat_A[167] * mat_B[244] +
//             mat_A[168] * mat_B[276] +
//             mat_A[169] * mat_B[308] +
//             mat_A[170] * mat_B[340] +
//             mat_A[171] * mat_B[372] +
//             mat_A[172] * mat_B[404] +
//             mat_A[173] * mat_B[436] +
//             mat_A[174] * mat_B[468] +
//             mat_A[175] * mat_B[500] +
//             mat_A[176] * mat_B[532] +
//             mat_A[177] * mat_B[564] +
//             mat_A[178] * mat_B[596] +
//             mat_A[179] * mat_B[628] +
//             mat_A[180] * mat_B[660] +
//             mat_A[181] * mat_B[692] +
//             mat_A[182] * mat_B[724] +
//             mat_A[183] * mat_B[756] +
//             mat_A[184] * mat_B[788] +
//             mat_A[185] * mat_B[820] +
//             mat_A[186] * mat_B[852] +
//             mat_A[187] * mat_B[884] +
//             mat_A[188] * mat_B[916] +
//             mat_A[189] * mat_B[948] +
//             mat_A[190] * mat_B[980] +
//             mat_A[191] * mat_B[1012];
//  mat_C[181] <= 
//             mat_A[160] * mat_B[21] +
//             mat_A[161] * mat_B[53] +
//             mat_A[162] * mat_B[85] +
//             mat_A[163] * mat_B[117] +
//             mat_A[164] * mat_B[149] +
//             mat_A[165] * mat_B[181] +
//             mat_A[166] * mat_B[213] +
//             mat_A[167] * mat_B[245] +
//             mat_A[168] * mat_B[277] +
//             mat_A[169] * mat_B[309] +
//             mat_A[170] * mat_B[341] +
//             mat_A[171] * mat_B[373] +
//             mat_A[172] * mat_B[405] +
//             mat_A[173] * mat_B[437] +
//             mat_A[174] * mat_B[469] +
//             mat_A[175] * mat_B[501] +
//             mat_A[176] * mat_B[533] +
//             mat_A[177] * mat_B[565] +
//             mat_A[178] * mat_B[597] +
//             mat_A[179] * mat_B[629] +
//             mat_A[180] * mat_B[661] +
//             mat_A[181] * mat_B[693] +
//             mat_A[182] * mat_B[725] +
//             mat_A[183] * mat_B[757] +
//             mat_A[184] * mat_B[789] +
//             mat_A[185] * mat_B[821] +
//             mat_A[186] * mat_B[853] +
//             mat_A[187] * mat_B[885] +
//             mat_A[188] * mat_B[917] +
//             mat_A[189] * mat_B[949] +
//             mat_A[190] * mat_B[981] +
//             mat_A[191] * mat_B[1013];
//  mat_C[182] <= 
//             mat_A[160] * mat_B[22] +
//             mat_A[161] * mat_B[54] +
//             mat_A[162] * mat_B[86] +
//             mat_A[163] * mat_B[118] +
//             mat_A[164] * mat_B[150] +
//             mat_A[165] * mat_B[182] +
//             mat_A[166] * mat_B[214] +
//             mat_A[167] * mat_B[246] +
//             mat_A[168] * mat_B[278] +
//             mat_A[169] * mat_B[310] +
//             mat_A[170] * mat_B[342] +
//             mat_A[171] * mat_B[374] +
//             mat_A[172] * mat_B[406] +
//             mat_A[173] * mat_B[438] +
//             mat_A[174] * mat_B[470] +
//             mat_A[175] * mat_B[502] +
//             mat_A[176] * mat_B[534] +
//             mat_A[177] * mat_B[566] +
//             mat_A[178] * mat_B[598] +
//             mat_A[179] * mat_B[630] +
//             mat_A[180] * mat_B[662] +
//             mat_A[181] * mat_B[694] +
//             mat_A[182] * mat_B[726] +
//             mat_A[183] * mat_B[758] +
//             mat_A[184] * mat_B[790] +
//             mat_A[185] * mat_B[822] +
//             mat_A[186] * mat_B[854] +
//             mat_A[187] * mat_B[886] +
//             mat_A[188] * mat_B[918] +
//             mat_A[189] * mat_B[950] +
//             mat_A[190] * mat_B[982] +
//             mat_A[191] * mat_B[1014];
//  mat_C[183] <= 
//             mat_A[160] * mat_B[23] +
//             mat_A[161] * mat_B[55] +
//             mat_A[162] * mat_B[87] +
//             mat_A[163] * mat_B[119] +
//             mat_A[164] * mat_B[151] +
//             mat_A[165] * mat_B[183] +
//             mat_A[166] * mat_B[215] +
//             mat_A[167] * mat_B[247] +
//             mat_A[168] * mat_B[279] +
//             mat_A[169] * mat_B[311] +
//             mat_A[170] * mat_B[343] +
//             mat_A[171] * mat_B[375] +
//             mat_A[172] * mat_B[407] +
//             mat_A[173] * mat_B[439] +
//             mat_A[174] * mat_B[471] +
//             mat_A[175] * mat_B[503] +
//             mat_A[176] * mat_B[535] +
//             mat_A[177] * mat_B[567] +
//             mat_A[178] * mat_B[599] +
//             mat_A[179] * mat_B[631] +
//             mat_A[180] * mat_B[663] +
//             mat_A[181] * mat_B[695] +
//             mat_A[182] * mat_B[727] +
//             mat_A[183] * mat_B[759] +
//             mat_A[184] * mat_B[791] +
//             mat_A[185] * mat_B[823] +
//             mat_A[186] * mat_B[855] +
//             mat_A[187] * mat_B[887] +
//             mat_A[188] * mat_B[919] +
//             mat_A[189] * mat_B[951] +
//             mat_A[190] * mat_B[983] +
//             mat_A[191] * mat_B[1015];
//  mat_C[184] <= 
//             mat_A[160] * mat_B[24] +
//             mat_A[161] * mat_B[56] +
//             mat_A[162] * mat_B[88] +
//             mat_A[163] * mat_B[120] +
//             mat_A[164] * mat_B[152] +
//             mat_A[165] * mat_B[184] +
//             mat_A[166] * mat_B[216] +
//             mat_A[167] * mat_B[248] +
//             mat_A[168] * mat_B[280] +
//             mat_A[169] * mat_B[312] +
//             mat_A[170] * mat_B[344] +
//             mat_A[171] * mat_B[376] +
//             mat_A[172] * mat_B[408] +
//             mat_A[173] * mat_B[440] +
//             mat_A[174] * mat_B[472] +
//             mat_A[175] * mat_B[504] +
//             mat_A[176] * mat_B[536] +
//             mat_A[177] * mat_B[568] +
//             mat_A[178] * mat_B[600] +
//             mat_A[179] * mat_B[632] +
//             mat_A[180] * mat_B[664] +
//             mat_A[181] * mat_B[696] +
//             mat_A[182] * mat_B[728] +
//             mat_A[183] * mat_B[760] +
//             mat_A[184] * mat_B[792] +
//             mat_A[185] * mat_B[824] +
//             mat_A[186] * mat_B[856] +
//             mat_A[187] * mat_B[888] +
//             mat_A[188] * mat_B[920] +
//             mat_A[189] * mat_B[952] +
//             mat_A[190] * mat_B[984] +
//             mat_A[191] * mat_B[1016];
//  mat_C[185] <= 
//             mat_A[160] * mat_B[25] +
//             mat_A[161] * mat_B[57] +
//             mat_A[162] * mat_B[89] +
//             mat_A[163] * mat_B[121] +
//             mat_A[164] * mat_B[153] +
//             mat_A[165] * mat_B[185] +
//             mat_A[166] * mat_B[217] +
//             mat_A[167] * mat_B[249] +
//             mat_A[168] * mat_B[281] +
//             mat_A[169] * mat_B[313] +
//             mat_A[170] * mat_B[345] +
//             mat_A[171] * mat_B[377] +
//             mat_A[172] * mat_B[409] +
//             mat_A[173] * mat_B[441] +
//             mat_A[174] * mat_B[473] +
//             mat_A[175] * mat_B[505] +
//             mat_A[176] * mat_B[537] +
//             mat_A[177] * mat_B[569] +
//             mat_A[178] * mat_B[601] +
//             mat_A[179] * mat_B[633] +
//             mat_A[180] * mat_B[665] +
//             mat_A[181] * mat_B[697] +
//             mat_A[182] * mat_B[729] +
//             mat_A[183] * mat_B[761] +
//             mat_A[184] * mat_B[793] +
//             mat_A[185] * mat_B[825] +
//             mat_A[186] * mat_B[857] +
//             mat_A[187] * mat_B[889] +
//             mat_A[188] * mat_B[921] +
//             mat_A[189] * mat_B[953] +
//             mat_A[190] * mat_B[985] +
//             mat_A[191] * mat_B[1017];
//  mat_C[186] <= 
//             mat_A[160] * mat_B[26] +
//             mat_A[161] * mat_B[58] +
//             mat_A[162] * mat_B[90] +
//             mat_A[163] * mat_B[122] +
//             mat_A[164] * mat_B[154] +
//             mat_A[165] * mat_B[186] +
//             mat_A[166] * mat_B[218] +
//             mat_A[167] * mat_B[250] +
//             mat_A[168] * mat_B[282] +
//             mat_A[169] * mat_B[314] +
//             mat_A[170] * mat_B[346] +
//             mat_A[171] * mat_B[378] +
//             mat_A[172] * mat_B[410] +
//             mat_A[173] * mat_B[442] +
//             mat_A[174] * mat_B[474] +
//             mat_A[175] * mat_B[506] +
//             mat_A[176] * mat_B[538] +
//             mat_A[177] * mat_B[570] +
//             mat_A[178] * mat_B[602] +
//             mat_A[179] * mat_B[634] +
//             mat_A[180] * mat_B[666] +
//             mat_A[181] * mat_B[698] +
//             mat_A[182] * mat_B[730] +
//             mat_A[183] * mat_B[762] +
//             mat_A[184] * mat_B[794] +
//             mat_A[185] * mat_B[826] +
//             mat_A[186] * mat_B[858] +
//             mat_A[187] * mat_B[890] +
//             mat_A[188] * mat_B[922] +
//             mat_A[189] * mat_B[954] +
//             mat_A[190] * mat_B[986] +
//             mat_A[191] * mat_B[1018];
//  mat_C[187] <= 
//             mat_A[160] * mat_B[27] +
//             mat_A[161] * mat_B[59] +
//             mat_A[162] * mat_B[91] +
//             mat_A[163] * mat_B[123] +
//             mat_A[164] * mat_B[155] +
//             mat_A[165] * mat_B[187] +
//             mat_A[166] * mat_B[219] +
//             mat_A[167] * mat_B[251] +
//             mat_A[168] * mat_B[283] +
//             mat_A[169] * mat_B[315] +
//             mat_A[170] * mat_B[347] +
//             mat_A[171] * mat_B[379] +
//             mat_A[172] * mat_B[411] +
//             mat_A[173] * mat_B[443] +
//             mat_A[174] * mat_B[475] +
//             mat_A[175] * mat_B[507] +
//             mat_A[176] * mat_B[539] +
//             mat_A[177] * mat_B[571] +
//             mat_A[178] * mat_B[603] +
//             mat_A[179] * mat_B[635] +
//             mat_A[180] * mat_B[667] +
//             mat_A[181] * mat_B[699] +
//             mat_A[182] * mat_B[731] +
//             mat_A[183] * mat_B[763] +
//             mat_A[184] * mat_B[795] +
//             mat_A[185] * mat_B[827] +
//             mat_A[186] * mat_B[859] +
//             mat_A[187] * mat_B[891] +
//             mat_A[188] * mat_B[923] +
//             mat_A[189] * mat_B[955] +
//             mat_A[190] * mat_B[987] +
//             mat_A[191] * mat_B[1019];
//  mat_C[188] <= 
//             mat_A[160] * mat_B[28] +
//             mat_A[161] * mat_B[60] +
//             mat_A[162] * mat_B[92] +
//             mat_A[163] * mat_B[124] +
//             mat_A[164] * mat_B[156] +
//             mat_A[165] * mat_B[188] +
//             mat_A[166] * mat_B[220] +
//             mat_A[167] * mat_B[252] +
//             mat_A[168] * mat_B[284] +
//             mat_A[169] * mat_B[316] +
//             mat_A[170] * mat_B[348] +
//             mat_A[171] * mat_B[380] +
//             mat_A[172] * mat_B[412] +
//             mat_A[173] * mat_B[444] +
//             mat_A[174] * mat_B[476] +
//             mat_A[175] * mat_B[508] +
//             mat_A[176] * mat_B[540] +
//             mat_A[177] * mat_B[572] +
//             mat_A[178] * mat_B[604] +
//             mat_A[179] * mat_B[636] +
//             mat_A[180] * mat_B[668] +
//             mat_A[181] * mat_B[700] +
//             mat_A[182] * mat_B[732] +
//             mat_A[183] * mat_B[764] +
//             mat_A[184] * mat_B[796] +
//             mat_A[185] * mat_B[828] +
//             mat_A[186] * mat_B[860] +
//             mat_A[187] * mat_B[892] +
//             mat_A[188] * mat_B[924] +
//             mat_A[189] * mat_B[956] +
//             mat_A[190] * mat_B[988] +
//             mat_A[191] * mat_B[1020];
//  mat_C[189] <= 
//             mat_A[160] * mat_B[29] +
//             mat_A[161] * mat_B[61] +
//             mat_A[162] * mat_B[93] +
//             mat_A[163] * mat_B[125] +
//             mat_A[164] * mat_B[157] +
//             mat_A[165] * mat_B[189] +
//             mat_A[166] * mat_B[221] +
//             mat_A[167] * mat_B[253] +
//             mat_A[168] * mat_B[285] +
//             mat_A[169] * mat_B[317] +
//             mat_A[170] * mat_B[349] +
//             mat_A[171] * mat_B[381] +
//             mat_A[172] * mat_B[413] +
//             mat_A[173] * mat_B[445] +
//             mat_A[174] * mat_B[477] +
//             mat_A[175] * mat_B[509] +
//             mat_A[176] * mat_B[541] +
//             mat_A[177] * mat_B[573] +
//             mat_A[178] * mat_B[605] +
//             mat_A[179] * mat_B[637] +
//             mat_A[180] * mat_B[669] +
//             mat_A[181] * mat_B[701] +
//             mat_A[182] * mat_B[733] +
//             mat_A[183] * mat_B[765] +
//             mat_A[184] * mat_B[797] +
//             mat_A[185] * mat_B[829] +
//             mat_A[186] * mat_B[861] +
//             mat_A[187] * mat_B[893] +
//             mat_A[188] * mat_B[925] +
//             mat_A[189] * mat_B[957] +
//             mat_A[190] * mat_B[989] +
//             mat_A[191] * mat_B[1021];
//  mat_C[190] <= 
//             mat_A[160] * mat_B[30] +
//             mat_A[161] * mat_B[62] +
//             mat_A[162] * mat_B[94] +
//             mat_A[163] * mat_B[126] +
//             mat_A[164] * mat_B[158] +
//             mat_A[165] * mat_B[190] +
//             mat_A[166] * mat_B[222] +
//             mat_A[167] * mat_B[254] +
//             mat_A[168] * mat_B[286] +
//             mat_A[169] * mat_B[318] +
//             mat_A[170] * mat_B[350] +
//             mat_A[171] * mat_B[382] +
//             mat_A[172] * mat_B[414] +
//             mat_A[173] * mat_B[446] +
//             mat_A[174] * mat_B[478] +
//             mat_A[175] * mat_B[510] +
//             mat_A[176] * mat_B[542] +
//             mat_A[177] * mat_B[574] +
//             mat_A[178] * mat_B[606] +
//             mat_A[179] * mat_B[638] +
//             mat_A[180] * mat_B[670] +
//             mat_A[181] * mat_B[702] +
//             mat_A[182] * mat_B[734] +
//             mat_A[183] * mat_B[766] +
//             mat_A[184] * mat_B[798] +
//             mat_A[185] * mat_B[830] +
//             mat_A[186] * mat_B[862] +
//             mat_A[187] * mat_B[894] +
//             mat_A[188] * mat_B[926] +
//             mat_A[189] * mat_B[958] +
//             mat_A[190] * mat_B[990] +
//             mat_A[191] * mat_B[1022];
//  mat_C[191] <= 
//             mat_A[160] * mat_B[31] +
//             mat_A[161] * mat_B[63] +
//             mat_A[162] * mat_B[95] +
//             mat_A[163] * mat_B[127] +
//             mat_A[164] * mat_B[159] +
//             mat_A[165] * mat_B[191] +
//             mat_A[166] * mat_B[223] +
//             mat_A[167] * mat_B[255] +
//             mat_A[168] * mat_B[287] +
//             mat_A[169] * mat_B[319] +
//             mat_A[170] * mat_B[351] +
//             mat_A[171] * mat_B[383] +
//             mat_A[172] * mat_B[415] +
//             mat_A[173] * mat_B[447] +
//             mat_A[174] * mat_B[479] +
//             mat_A[175] * mat_B[511] +
//             mat_A[176] * mat_B[543] +
//             mat_A[177] * mat_B[575] +
//             mat_A[178] * mat_B[607] +
//             mat_A[179] * mat_B[639] +
//             mat_A[180] * mat_B[671] +
//             mat_A[181] * mat_B[703] +
//             mat_A[182] * mat_B[735] +
//             mat_A[183] * mat_B[767] +
//             mat_A[184] * mat_B[799] +
//             mat_A[185] * mat_B[831] +
//             mat_A[186] * mat_B[863] +
//             mat_A[187] * mat_B[895] +
//             mat_A[188] * mat_B[927] +
//             mat_A[189] * mat_B[959] +
//             mat_A[190] * mat_B[991] +
//             mat_A[191] * mat_B[1023];
//  mat_C[192] <= 
//             mat_A[192] * mat_B[0] +
//             mat_A[193] * mat_B[32] +
//             mat_A[194] * mat_B[64] +
//             mat_A[195] * mat_B[96] +
//             mat_A[196] * mat_B[128] +
//             mat_A[197] * mat_B[160] +
//             mat_A[198] * mat_B[192] +
//             mat_A[199] * mat_B[224] +
//             mat_A[200] * mat_B[256] +
//             mat_A[201] * mat_B[288] +
//             mat_A[202] * mat_B[320] +
//             mat_A[203] * mat_B[352] +
//             mat_A[204] * mat_B[384] +
//             mat_A[205] * mat_B[416] +
//             mat_A[206] * mat_B[448] +
//             mat_A[207] * mat_B[480] +
//             mat_A[208] * mat_B[512] +
//             mat_A[209] * mat_B[544] +
//             mat_A[210] * mat_B[576] +
//             mat_A[211] * mat_B[608] +
//             mat_A[212] * mat_B[640] +
//             mat_A[213] * mat_B[672] +
//             mat_A[214] * mat_B[704] +
//             mat_A[215] * mat_B[736] +
//             mat_A[216] * mat_B[768] +
//             mat_A[217] * mat_B[800] +
//             mat_A[218] * mat_B[832] +
//             mat_A[219] * mat_B[864] +
//             mat_A[220] * mat_B[896] +
//             mat_A[221] * mat_B[928] +
//             mat_A[222] * mat_B[960] +
//             mat_A[223] * mat_B[992];
//  mat_C[193] <= 
//             mat_A[192] * mat_B[1] +
//             mat_A[193] * mat_B[33] +
//             mat_A[194] * mat_B[65] +
//             mat_A[195] * mat_B[97] +
//             mat_A[196] * mat_B[129] +
//             mat_A[197] * mat_B[161] +
//             mat_A[198] * mat_B[193] +
//             mat_A[199] * mat_B[225] +
//             mat_A[200] * mat_B[257] +
//             mat_A[201] * mat_B[289] +
//             mat_A[202] * mat_B[321] +
//             mat_A[203] * mat_B[353] +
//             mat_A[204] * mat_B[385] +
//             mat_A[205] * mat_B[417] +
//             mat_A[206] * mat_B[449] +
//             mat_A[207] * mat_B[481] +
//             mat_A[208] * mat_B[513] +
//             mat_A[209] * mat_B[545] +
//             mat_A[210] * mat_B[577] +
//             mat_A[211] * mat_B[609] +
//             mat_A[212] * mat_B[641] +
//             mat_A[213] * mat_B[673] +
//             mat_A[214] * mat_B[705] +
//             mat_A[215] * mat_B[737] +
//             mat_A[216] * mat_B[769] +
//             mat_A[217] * mat_B[801] +
//             mat_A[218] * mat_B[833] +
//             mat_A[219] * mat_B[865] +
//             mat_A[220] * mat_B[897] +
//             mat_A[221] * mat_B[929] +
//             mat_A[222] * mat_B[961] +
//             mat_A[223] * mat_B[993];
//  mat_C[194] <= 
//             mat_A[192] * mat_B[2] +
//             mat_A[193] * mat_B[34] +
//             mat_A[194] * mat_B[66] +
//             mat_A[195] * mat_B[98] +
//             mat_A[196] * mat_B[130] +
//             mat_A[197] * mat_B[162] +
//             mat_A[198] * mat_B[194] +
//             mat_A[199] * mat_B[226] +
//             mat_A[200] * mat_B[258] +
//             mat_A[201] * mat_B[290] +
//             mat_A[202] * mat_B[322] +
//             mat_A[203] * mat_B[354] +
//             mat_A[204] * mat_B[386] +
//             mat_A[205] * mat_B[418] +
//             mat_A[206] * mat_B[450] +
//             mat_A[207] * mat_B[482] +
//             mat_A[208] * mat_B[514] +
//             mat_A[209] * mat_B[546] +
//             mat_A[210] * mat_B[578] +
//             mat_A[211] * mat_B[610] +
//             mat_A[212] * mat_B[642] +
//             mat_A[213] * mat_B[674] +
//             mat_A[214] * mat_B[706] +
//             mat_A[215] * mat_B[738] +
//             mat_A[216] * mat_B[770] +
//             mat_A[217] * mat_B[802] +
//             mat_A[218] * mat_B[834] +
//             mat_A[219] * mat_B[866] +
//             mat_A[220] * mat_B[898] +
//             mat_A[221] * mat_B[930] +
//             mat_A[222] * mat_B[962] +
//             mat_A[223] * mat_B[994];
//  mat_C[195] <= 
//             mat_A[192] * mat_B[3] +
//             mat_A[193] * mat_B[35] +
//             mat_A[194] * mat_B[67] +
//             mat_A[195] * mat_B[99] +
//             mat_A[196] * mat_B[131] +
//             mat_A[197] * mat_B[163] +
//             mat_A[198] * mat_B[195] +
//             mat_A[199] * mat_B[227] +
//             mat_A[200] * mat_B[259] +
//             mat_A[201] * mat_B[291] +
//             mat_A[202] * mat_B[323] +
//             mat_A[203] * mat_B[355] +
//             mat_A[204] * mat_B[387] +
//             mat_A[205] * mat_B[419] +
//             mat_A[206] * mat_B[451] +
//             mat_A[207] * mat_B[483] +
//             mat_A[208] * mat_B[515] +
//             mat_A[209] * mat_B[547] +
//             mat_A[210] * mat_B[579] +
//             mat_A[211] * mat_B[611] +
//             mat_A[212] * mat_B[643] +
//             mat_A[213] * mat_B[675] +
//             mat_A[214] * mat_B[707] +
//             mat_A[215] * mat_B[739] +
//             mat_A[216] * mat_B[771] +
//             mat_A[217] * mat_B[803] +
//             mat_A[218] * mat_B[835] +
//             mat_A[219] * mat_B[867] +
//             mat_A[220] * mat_B[899] +
//             mat_A[221] * mat_B[931] +
//             mat_A[222] * mat_B[963] +
//             mat_A[223] * mat_B[995];
//  mat_C[196] <= 
//             mat_A[192] * mat_B[4] +
//             mat_A[193] * mat_B[36] +
//             mat_A[194] * mat_B[68] +
//             mat_A[195] * mat_B[100] +
//             mat_A[196] * mat_B[132] +
//             mat_A[197] * mat_B[164] +
//             mat_A[198] * mat_B[196] +
//             mat_A[199] * mat_B[228] +
//             mat_A[200] * mat_B[260] +
//             mat_A[201] * mat_B[292] +
//             mat_A[202] * mat_B[324] +
//             mat_A[203] * mat_B[356] +
//             mat_A[204] * mat_B[388] +
//             mat_A[205] * mat_B[420] +
//             mat_A[206] * mat_B[452] +
//             mat_A[207] * mat_B[484] +
//             mat_A[208] * mat_B[516] +
//             mat_A[209] * mat_B[548] +
//             mat_A[210] * mat_B[580] +
//             mat_A[211] * mat_B[612] +
//             mat_A[212] * mat_B[644] +
//             mat_A[213] * mat_B[676] +
//             mat_A[214] * mat_B[708] +
//             mat_A[215] * mat_B[740] +
//             mat_A[216] * mat_B[772] +
//             mat_A[217] * mat_B[804] +
//             mat_A[218] * mat_B[836] +
//             mat_A[219] * mat_B[868] +
//             mat_A[220] * mat_B[900] +
//             mat_A[221] * mat_B[932] +
//             mat_A[222] * mat_B[964] +
//             mat_A[223] * mat_B[996];
//  mat_C[197] <= 
//             mat_A[192] * mat_B[5] +
//             mat_A[193] * mat_B[37] +
//             mat_A[194] * mat_B[69] +
//             mat_A[195] * mat_B[101] +
//             mat_A[196] * mat_B[133] +
//             mat_A[197] * mat_B[165] +
//             mat_A[198] * mat_B[197] +
//             mat_A[199] * mat_B[229] +
//             mat_A[200] * mat_B[261] +
//             mat_A[201] * mat_B[293] +
//             mat_A[202] * mat_B[325] +
//             mat_A[203] * mat_B[357] +
//             mat_A[204] * mat_B[389] +
//             mat_A[205] * mat_B[421] +
//             mat_A[206] * mat_B[453] +
//             mat_A[207] * mat_B[485] +
//             mat_A[208] * mat_B[517] +
//             mat_A[209] * mat_B[549] +
//             mat_A[210] * mat_B[581] +
//             mat_A[211] * mat_B[613] +
//             mat_A[212] * mat_B[645] +
//             mat_A[213] * mat_B[677] +
//             mat_A[214] * mat_B[709] +
//             mat_A[215] * mat_B[741] +
//             mat_A[216] * mat_B[773] +
//             mat_A[217] * mat_B[805] +
//             mat_A[218] * mat_B[837] +
//             mat_A[219] * mat_B[869] +
//             mat_A[220] * mat_B[901] +
//             mat_A[221] * mat_B[933] +
//             mat_A[222] * mat_B[965] +
//             mat_A[223] * mat_B[997];
//  mat_C[198] <= 
//             mat_A[192] * mat_B[6] +
//             mat_A[193] * mat_B[38] +
//             mat_A[194] * mat_B[70] +
//             mat_A[195] * mat_B[102] +
//             mat_A[196] * mat_B[134] +
//             mat_A[197] * mat_B[166] +
//             mat_A[198] * mat_B[198] +
//             mat_A[199] * mat_B[230] +
//             mat_A[200] * mat_B[262] +
//             mat_A[201] * mat_B[294] +
//             mat_A[202] * mat_B[326] +
//             mat_A[203] * mat_B[358] +
//             mat_A[204] * mat_B[390] +
//             mat_A[205] * mat_B[422] +
//             mat_A[206] * mat_B[454] +
//             mat_A[207] * mat_B[486] +
//             mat_A[208] * mat_B[518] +
//             mat_A[209] * mat_B[550] +
//             mat_A[210] * mat_B[582] +
//             mat_A[211] * mat_B[614] +
//             mat_A[212] * mat_B[646] +
//             mat_A[213] * mat_B[678] +
//             mat_A[214] * mat_B[710] +
//             mat_A[215] * mat_B[742] +
//             mat_A[216] * mat_B[774] +
//             mat_A[217] * mat_B[806] +
//             mat_A[218] * mat_B[838] +
//             mat_A[219] * mat_B[870] +
//             mat_A[220] * mat_B[902] +
//             mat_A[221] * mat_B[934] +
//             mat_A[222] * mat_B[966] +
//             mat_A[223] * mat_B[998];
//  mat_C[199] <= 
//             mat_A[192] * mat_B[7] +
//             mat_A[193] * mat_B[39] +
//             mat_A[194] * mat_B[71] +
//             mat_A[195] * mat_B[103] +
//             mat_A[196] * mat_B[135] +
//             mat_A[197] * mat_B[167] +
//             mat_A[198] * mat_B[199] +
//             mat_A[199] * mat_B[231] +
//             mat_A[200] * mat_B[263] +
//             mat_A[201] * mat_B[295] +
//             mat_A[202] * mat_B[327] +
//             mat_A[203] * mat_B[359] +
//             mat_A[204] * mat_B[391] +
//             mat_A[205] * mat_B[423] +
//             mat_A[206] * mat_B[455] +
//             mat_A[207] * mat_B[487] +
//             mat_A[208] * mat_B[519] +
//             mat_A[209] * mat_B[551] +
//             mat_A[210] * mat_B[583] +
//             mat_A[211] * mat_B[615] +
//             mat_A[212] * mat_B[647] +
//             mat_A[213] * mat_B[679] +
//             mat_A[214] * mat_B[711] +
//             mat_A[215] * mat_B[743] +
//             mat_A[216] * mat_B[775] +
//             mat_A[217] * mat_B[807] +
//             mat_A[218] * mat_B[839] +
//             mat_A[219] * mat_B[871] +
//             mat_A[220] * mat_B[903] +
//             mat_A[221] * mat_B[935] +
//             mat_A[222] * mat_B[967] +
//             mat_A[223] * mat_B[999];
//  mat_C[200] <= 
//             mat_A[192] * mat_B[8] +
//             mat_A[193] * mat_B[40] +
//             mat_A[194] * mat_B[72] +
//             mat_A[195] * mat_B[104] +
//             mat_A[196] * mat_B[136] +
//             mat_A[197] * mat_B[168] +
//             mat_A[198] * mat_B[200] +
//             mat_A[199] * mat_B[232] +
//             mat_A[200] * mat_B[264] +
//             mat_A[201] * mat_B[296] +
//             mat_A[202] * mat_B[328] +
//             mat_A[203] * mat_B[360] +
//             mat_A[204] * mat_B[392] +
//             mat_A[205] * mat_B[424] +
//             mat_A[206] * mat_B[456] +
//             mat_A[207] * mat_B[488] +
//             mat_A[208] * mat_B[520] +
//             mat_A[209] * mat_B[552] +
//             mat_A[210] * mat_B[584] +
//             mat_A[211] * mat_B[616] +
//             mat_A[212] * mat_B[648] +
//             mat_A[213] * mat_B[680] +
//             mat_A[214] * mat_B[712] +
//             mat_A[215] * mat_B[744] +
//             mat_A[216] * mat_B[776] +
//             mat_A[217] * mat_B[808] +
//             mat_A[218] * mat_B[840] +
//             mat_A[219] * mat_B[872] +
//             mat_A[220] * mat_B[904] +
//             mat_A[221] * mat_B[936] +
//             mat_A[222] * mat_B[968] +
//             mat_A[223] * mat_B[1000];
//  mat_C[201] <= 
//             mat_A[192] * mat_B[9] +
//             mat_A[193] * mat_B[41] +
//             mat_A[194] * mat_B[73] +
//             mat_A[195] * mat_B[105] +
//             mat_A[196] * mat_B[137] +
//             mat_A[197] * mat_B[169] +
//             mat_A[198] * mat_B[201] +
//             mat_A[199] * mat_B[233] +
//             mat_A[200] * mat_B[265] +
//             mat_A[201] * mat_B[297] +
//             mat_A[202] * mat_B[329] +
//             mat_A[203] * mat_B[361] +
//             mat_A[204] * mat_B[393] +
//             mat_A[205] * mat_B[425] +
//             mat_A[206] * mat_B[457] +
//             mat_A[207] * mat_B[489] +
//             mat_A[208] * mat_B[521] +
//             mat_A[209] * mat_B[553] +
//             mat_A[210] * mat_B[585] +
//             mat_A[211] * mat_B[617] +
//             mat_A[212] * mat_B[649] +
//             mat_A[213] * mat_B[681] +
//             mat_A[214] * mat_B[713] +
//             mat_A[215] * mat_B[745] +
//             mat_A[216] * mat_B[777] +
//             mat_A[217] * mat_B[809] +
//             mat_A[218] * mat_B[841] +
//             mat_A[219] * mat_B[873] +
//             mat_A[220] * mat_B[905] +
//             mat_A[221] * mat_B[937] +
//             mat_A[222] * mat_B[969] +
//             mat_A[223] * mat_B[1001];
//  mat_C[202] <= 
//             mat_A[192] * mat_B[10] +
//             mat_A[193] * mat_B[42] +
//             mat_A[194] * mat_B[74] +
//             mat_A[195] * mat_B[106] +
//             mat_A[196] * mat_B[138] +
//             mat_A[197] * mat_B[170] +
//             mat_A[198] * mat_B[202] +
//             mat_A[199] * mat_B[234] +
//             mat_A[200] * mat_B[266] +
//             mat_A[201] * mat_B[298] +
//             mat_A[202] * mat_B[330] +
//             mat_A[203] * mat_B[362] +
//             mat_A[204] * mat_B[394] +
//             mat_A[205] * mat_B[426] +
//             mat_A[206] * mat_B[458] +
//             mat_A[207] * mat_B[490] +
//             mat_A[208] * mat_B[522] +
//             mat_A[209] * mat_B[554] +
//             mat_A[210] * mat_B[586] +
//             mat_A[211] * mat_B[618] +
//             mat_A[212] * mat_B[650] +
//             mat_A[213] * mat_B[682] +
//             mat_A[214] * mat_B[714] +
//             mat_A[215] * mat_B[746] +
//             mat_A[216] * mat_B[778] +
//             mat_A[217] * mat_B[810] +
//             mat_A[218] * mat_B[842] +
//             mat_A[219] * mat_B[874] +
//             mat_A[220] * mat_B[906] +
//             mat_A[221] * mat_B[938] +
//             mat_A[222] * mat_B[970] +
//             mat_A[223] * mat_B[1002];
//  mat_C[203] <= 
//             mat_A[192] * mat_B[11] +
//             mat_A[193] * mat_B[43] +
//             mat_A[194] * mat_B[75] +
//             mat_A[195] * mat_B[107] +
//             mat_A[196] * mat_B[139] +
//             mat_A[197] * mat_B[171] +
//             mat_A[198] * mat_B[203] +
//             mat_A[199] * mat_B[235] +
//             mat_A[200] * mat_B[267] +
//             mat_A[201] * mat_B[299] +
//             mat_A[202] * mat_B[331] +
//             mat_A[203] * mat_B[363] +
//             mat_A[204] * mat_B[395] +
//             mat_A[205] * mat_B[427] +
//             mat_A[206] * mat_B[459] +
//             mat_A[207] * mat_B[491] +
//             mat_A[208] * mat_B[523] +
//             mat_A[209] * mat_B[555] +
//             mat_A[210] * mat_B[587] +
//             mat_A[211] * mat_B[619] +
//             mat_A[212] * mat_B[651] +
//             mat_A[213] * mat_B[683] +
//             mat_A[214] * mat_B[715] +
//             mat_A[215] * mat_B[747] +
//             mat_A[216] * mat_B[779] +
//             mat_A[217] * mat_B[811] +
//             mat_A[218] * mat_B[843] +
//             mat_A[219] * mat_B[875] +
//             mat_A[220] * mat_B[907] +
//             mat_A[221] * mat_B[939] +
//             mat_A[222] * mat_B[971] +
//             mat_A[223] * mat_B[1003];
//  mat_C[204] <= 
//             mat_A[192] * mat_B[12] +
//             mat_A[193] * mat_B[44] +
//             mat_A[194] * mat_B[76] +
//             mat_A[195] * mat_B[108] +
//             mat_A[196] * mat_B[140] +
//             mat_A[197] * mat_B[172] +
//             mat_A[198] * mat_B[204] +
//             mat_A[199] * mat_B[236] +
//             mat_A[200] * mat_B[268] +
//             mat_A[201] * mat_B[300] +
//             mat_A[202] * mat_B[332] +
//             mat_A[203] * mat_B[364] +
//             mat_A[204] * mat_B[396] +
//             mat_A[205] * mat_B[428] +
//             mat_A[206] * mat_B[460] +
//             mat_A[207] * mat_B[492] +
//             mat_A[208] * mat_B[524] +
//             mat_A[209] * mat_B[556] +
//             mat_A[210] * mat_B[588] +
//             mat_A[211] * mat_B[620] +
//             mat_A[212] * mat_B[652] +
//             mat_A[213] * mat_B[684] +
//             mat_A[214] * mat_B[716] +
//             mat_A[215] * mat_B[748] +
//             mat_A[216] * mat_B[780] +
//             mat_A[217] * mat_B[812] +
//             mat_A[218] * mat_B[844] +
//             mat_A[219] * mat_B[876] +
//             mat_A[220] * mat_B[908] +
//             mat_A[221] * mat_B[940] +
//             mat_A[222] * mat_B[972] +
//             mat_A[223] * mat_B[1004];
//  mat_C[205] <= 
//             mat_A[192] * mat_B[13] +
//             mat_A[193] * mat_B[45] +
//             mat_A[194] * mat_B[77] +
//             mat_A[195] * mat_B[109] +
//             mat_A[196] * mat_B[141] +
//             mat_A[197] * mat_B[173] +
//             mat_A[198] * mat_B[205] +
//             mat_A[199] * mat_B[237] +
//             mat_A[200] * mat_B[269] +
//             mat_A[201] * mat_B[301] +
//             mat_A[202] * mat_B[333] +
//             mat_A[203] * mat_B[365] +
//             mat_A[204] * mat_B[397] +
//             mat_A[205] * mat_B[429] +
//             mat_A[206] * mat_B[461] +
//             mat_A[207] * mat_B[493] +
//             mat_A[208] * mat_B[525] +
//             mat_A[209] * mat_B[557] +
//             mat_A[210] * mat_B[589] +
//             mat_A[211] * mat_B[621] +
//             mat_A[212] * mat_B[653] +
//             mat_A[213] * mat_B[685] +
//             mat_A[214] * mat_B[717] +
//             mat_A[215] * mat_B[749] +
//             mat_A[216] * mat_B[781] +
//             mat_A[217] * mat_B[813] +
//             mat_A[218] * mat_B[845] +
//             mat_A[219] * mat_B[877] +
//             mat_A[220] * mat_B[909] +
//             mat_A[221] * mat_B[941] +
//             mat_A[222] * mat_B[973] +
//             mat_A[223] * mat_B[1005];
//  mat_C[206] <= 
//             mat_A[192] * mat_B[14] +
//             mat_A[193] * mat_B[46] +
//             mat_A[194] * mat_B[78] +
//             mat_A[195] * mat_B[110] +
//             mat_A[196] * mat_B[142] +
//             mat_A[197] * mat_B[174] +
//             mat_A[198] * mat_B[206] +
//             mat_A[199] * mat_B[238] +
//             mat_A[200] * mat_B[270] +
//             mat_A[201] * mat_B[302] +
//             mat_A[202] * mat_B[334] +
//             mat_A[203] * mat_B[366] +
//             mat_A[204] * mat_B[398] +
//             mat_A[205] * mat_B[430] +
//             mat_A[206] * mat_B[462] +
//             mat_A[207] * mat_B[494] +
//             mat_A[208] * mat_B[526] +
//             mat_A[209] * mat_B[558] +
//             mat_A[210] * mat_B[590] +
//             mat_A[211] * mat_B[622] +
//             mat_A[212] * mat_B[654] +
//             mat_A[213] * mat_B[686] +
//             mat_A[214] * mat_B[718] +
//             mat_A[215] * mat_B[750] +
//             mat_A[216] * mat_B[782] +
//             mat_A[217] * mat_B[814] +
//             mat_A[218] * mat_B[846] +
//             mat_A[219] * mat_B[878] +
//             mat_A[220] * mat_B[910] +
//             mat_A[221] * mat_B[942] +
//             mat_A[222] * mat_B[974] +
//             mat_A[223] * mat_B[1006];
//  mat_C[207] <= 
//             mat_A[192] * mat_B[15] +
//             mat_A[193] * mat_B[47] +
//             mat_A[194] * mat_B[79] +
//             mat_A[195] * mat_B[111] +
//             mat_A[196] * mat_B[143] +
//             mat_A[197] * mat_B[175] +
//             mat_A[198] * mat_B[207] +
//             mat_A[199] * mat_B[239] +
//             mat_A[200] * mat_B[271] +
//             mat_A[201] * mat_B[303] +
//             mat_A[202] * mat_B[335] +
//             mat_A[203] * mat_B[367] +
//             mat_A[204] * mat_B[399] +
//             mat_A[205] * mat_B[431] +
//             mat_A[206] * mat_B[463] +
//             mat_A[207] * mat_B[495] +
//             mat_A[208] * mat_B[527] +
//             mat_A[209] * mat_B[559] +
//             mat_A[210] * mat_B[591] +
//             mat_A[211] * mat_B[623] +
//             mat_A[212] * mat_B[655] +
//             mat_A[213] * mat_B[687] +
//             mat_A[214] * mat_B[719] +
//             mat_A[215] * mat_B[751] +
//             mat_A[216] * mat_B[783] +
//             mat_A[217] * mat_B[815] +
//             mat_A[218] * mat_B[847] +
//             mat_A[219] * mat_B[879] +
//             mat_A[220] * mat_B[911] +
//             mat_A[221] * mat_B[943] +
//             mat_A[222] * mat_B[975] +
//             mat_A[223] * mat_B[1007];
//  mat_C[208] <= 
//             mat_A[192] * mat_B[16] +
//             mat_A[193] * mat_B[48] +
//             mat_A[194] * mat_B[80] +
//             mat_A[195] * mat_B[112] +
//             mat_A[196] * mat_B[144] +
//             mat_A[197] * mat_B[176] +
//             mat_A[198] * mat_B[208] +
//             mat_A[199] * mat_B[240] +
//             mat_A[200] * mat_B[272] +
//             mat_A[201] * mat_B[304] +
//             mat_A[202] * mat_B[336] +
//             mat_A[203] * mat_B[368] +
//             mat_A[204] * mat_B[400] +
//             mat_A[205] * mat_B[432] +
//             mat_A[206] * mat_B[464] +
//             mat_A[207] * mat_B[496] +
//             mat_A[208] * mat_B[528] +
//             mat_A[209] * mat_B[560] +
//             mat_A[210] * mat_B[592] +
//             mat_A[211] * mat_B[624] +
//             mat_A[212] * mat_B[656] +
//             mat_A[213] * mat_B[688] +
//             mat_A[214] * mat_B[720] +
//             mat_A[215] * mat_B[752] +
//             mat_A[216] * mat_B[784] +
//             mat_A[217] * mat_B[816] +
//             mat_A[218] * mat_B[848] +
//             mat_A[219] * mat_B[880] +
//             mat_A[220] * mat_B[912] +
//             mat_A[221] * mat_B[944] +
//             mat_A[222] * mat_B[976] +
//             mat_A[223] * mat_B[1008];
//  mat_C[209] <= 
//             mat_A[192] * mat_B[17] +
//             mat_A[193] * mat_B[49] +
//             mat_A[194] * mat_B[81] +
//             mat_A[195] * mat_B[113] +
//             mat_A[196] * mat_B[145] +
//             mat_A[197] * mat_B[177] +
//             mat_A[198] * mat_B[209] +
//             mat_A[199] * mat_B[241] +
//             mat_A[200] * mat_B[273] +
//             mat_A[201] * mat_B[305] +
//             mat_A[202] * mat_B[337] +
//             mat_A[203] * mat_B[369] +
//             mat_A[204] * mat_B[401] +
//             mat_A[205] * mat_B[433] +
//             mat_A[206] * mat_B[465] +
//             mat_A[207] * mat_B[497] +
//             mat_A[208] * mat_B[529] +
//             mat_A[209] * mat_B[561] +
//             mat_A[210] * mat_B[593] +
//             mat_A[211] * mat_B[625] +
//             mat_A[212] * mat_B[657] +
//             mat_A[213] * mat_B[689] +
//             mat_A[214] * mat_B[721] +
//             mat_A[215] * mat_B[753] +
//             mat_A[216] * mat_B[785] +
//             mat_A[217] * mat_B[817] +
//             mat_A[218] * mat_B[849] +
//             mat_A[219] * mat_B[881] +
//             mat_A[220] * mat_B[913] +
//             mat_A[221] * mat_B[945] +
//             mat_A[222] * mat_B[977] +
//             mat_A[223] * mat_B[1009];
//  mat_C[210] <= 
//             mat_A[192] * mat_B[18] +
//             mat_A[193] * mat_B[50] +
//             mat_A[194] * mat_B[82] +
//             mat_A[195] * mat_B[114] +
//             mat_A[196] * mat_B[146] +
//             mat_A[197] * mat_B[178] +
//             mat_A[198] * mat_B[210] +
//             mat_A[199] * mat_B[242] +
//             mat_A[200] * mat_B[274] +
//             mat_A[201] * mat_B[306] +
//             mat_A[202] * mat_B[338] +
//             mat_A[203] * mat_B[370] +
//             mat_A[204] * mat_B[402] +
//             mat_A[205] * mat_B[434] +
//             mat_A[206] * mat_B[466] +
//             mat_A[207] * mat_B[498] +
//             mat_A[208] * mat_B[530] +
//             mat_A[209] * mat_B[562] +
//             mat_A[210] * mat_B[594] +
//             mat_A[211] * mat_B[626] +
//             mat_A[212] * mat_B[658] +
//             mat_A[213] * mat_B[690] +
//             mat_A[214] * mat_B[722] +
//             mat_A[215] * mat_B[754] +
//             mat_A[216] * mat_B[786] +
//             mat_A[217] * mat_B[818] +
//             mat_A[218] * mat_B[850] +
//             mat_A[219] * mat_B[882] +
//             mat_A[220] * mat_B[914] +
//             mat_A[221] * mat_B[946] +
//             mat_A[222] * mat_B[978] +
//             mat_A[223] * mat_B[1010];
//  mat_C[211] <= 
//             mat_A[192] * mat_B[19] +
//             mat_A[193] * mat_B[51] +
//             mat_A[194] * mat_B[83] +
//             mat_A[195] * mat_B[115] +
//             mat_A[196] * mat_B[147] +
//             mat_A[197] * mat_B[179] +
//             mat_A[198] * mat_B[211] +
//             mat_A[199] * mat_B[243] +
//             mat_A[200] * mat_B[275] +
//             mat_A[201] * mat_B[307] +
//             mat_A[202] * mat_B[339] +
//             mat_A[203] * mat_B[371] +
//             mat_A[204] * mat_B[403] +
//             mat_A[205] * mat_B[435] +
//             mat_A[206] * mat_B[467] +
//             mat_A[207] * mat_B[499] +
//             mat_A[208] * mat_B[531] +
//             mat_A[209] * mat_B[563] +
//             mat_A[210] * mat_B[595] +
//             mat_A[211] * mat_B[627] +
//             mat_A[212] * mat_B[659] +
//             mat_A[213] * mat_B[691] +
//             mat_A[214] * mat_B[723] +
//             mat_A[215] * mat_B[755] +
//             mat_A[216] * mat_B[787] +
//             mat_A[217] * mat_B[819] +
//             mat_A[218] * mat_B[851] +
//             mat_A[219] * mat_B[883] +
//             mat_A[220] * mat_B[915] +
//             mat_A[221] * mat_B[947] +
//             mat_A[222] * mat_B[979] +
//             mat_A[223] * mat_B[1011];
//  mat_C[212] <= 
//             mat_A[192] * mat_B[20] +
//             mat_A[193] * mat_B[52] +
//             mat_A[194] * mat_B[84] +
//             mat_A[195] * mat_B[116] +
//             mat_A[196] * mat_B[148] +
//             mat_A[197] * mat_B[180] +
//             mat_A[198] * mat_B[212] +
//             mat_A[199] * mat_B[244] +
//             mat_A[200] * mat_B[276] +
//             mat_A[201] * mat_B[308] +
//             mat_A[202] * mat_B[340] +
//             mat_A[203] * mat_B[372] +
//             mat_A[204] * mat_B[404] +
//             mat_A[205] * mat_B[436] +
//             mat_A[206] * mat_B[468] +
//             mat_A[207] * mat_B[500] +
//             mat_A[208] * mat_B[532] +
//             mat_A[209] * mat_B[564] +
//             mat_A[210] * mat_B[596] +
//             mat_A[211] * mat_B[628] +
//             mat_A[212] * mat_B[660] +
//             mat_A[213] * mat_B[692] +
//             mat_A[214] * mat_B[724] +
//             mat_A[215] * mat_B[756] +
//             mat_A[216] * mat_B[788] +
//             mat_A[217] * mat_B[820] +
//             mat_A[218] * mat_B[852] +
//             mat_A[219] * mat_B[884] +
//             mat_A[220] * mat_B[916] +
//             mat_A[221] * mat_B[948] +
//             mat_A[222] * mat_B[980] +
//             mat_A[223] * mat_B[1012];
//  mat_C[213] <= 
//             mat_A[192] * mat_B[21] +
//             mat_A[193] * mat_B[53] +
//             mat_A[194] * mat_B[85] +
//             mat_A[195] * mat_B[117] +
//             mat_A[196] * mat_B[149] +
//             mat_A[197] * mat_B[181] +
//             mat_A[198] * mat_B[213] +
//             mat_A[199] * mat_B[245] +
//             mat_A[200] * mat_B[277] +
//             mat_A[201] * mat_B[309] +
//             mat_A[202] * mat_B[341] +
//             mat_A[203] * mat_B[373] +
//             mat_A[204] * mat_B[405] +
//             mat_A[205] * mat_B[437] +
//             mat_A[206] * mat_B[469] +
//             mat_A[207] * mat_B[501] +
//             mat_A[208] * mat_B[533] +
//             mat_A[209] * mat_B[565] +
//             mat_A[210] * mat_B[597] +
//             mat_A[211] * mat_B[629] +
//             mat_A[212] * mat_B[661] +
//             mat_A[213] * mat_B[693] +
//             mat_A[214] * mat_B[725] +
//             mat_A[215] * mat_B[757] +
//             mat_A[216] * mat_B[789] +
//             mat_A[217] * mat_B[821] +
//             mat_A[218] * mat_B[853] +
//             mat_A[219] * mat_B[885] +
//             mat_A[220] * mat_B[917] +
//             mat_A[221] * mat_B[949] +
//             mat_A[222] * mat_B[981] +
//             mat_A[223] * mat_B[1013];
//  mat_C[214] <= 
//             mat_A[192] * mat_B[22] +
//             mat_A[193] * mat_B[54] +
//             mat_A[194] * mat_B[86] +
//             mat_A[195] * mat_B[118] +
//             mat_A[196] * mat_B[150] +
//             mat_A[197] * mat_B[182] +
//             mat_A[198] * mat_B[214] +
//             mat_A[199] * mat_B[246] +
//             mat_A[200] * mat_B[278] +
//             mat_A[201] * mat_B[310] +
//             mat_A[202] * mat_B[342] +
//             mat_A[203] * mat_B[374] +
//             mat_A[204] * mat_B[406] +
//             mat_A[205] * mat_B[438] +
//             mat_A[206] * mat_B[470] +
//             mat_A[207] * mat_B[502] +
//             mat_A[208] * mat_B[534] +
//             mat_A[209] * mat_B[566] +
//             mat_A[210] * mat_B[598] +
//             mat_A[211] * mat_B[630] +
//             mat_A[212] * mat_B[662] +
//             mat_A[213] * mat_B[694] +
//             mat_A[214] * mat_B[726] +
//             mat_A[215] * mat_B[758] +
//             mat_A[216] * mat_B[790] +
//             mat_A[217] * mat_B[822] +
//             mat_A[218] * mat_B[854] +
//             mat_A[219] * mat_B[886] +
//             mat_A[220] * mat_B[918] +
//             mat_A[221] * mat_B[950] +
//             mat_A[222] * mat_B[982] +
//             mat_A[223] * mat_B[1014];
//  mat_C[215] <= 
//             mat_A[192] * mat_B[23] +
//             mat_A[193] * mat_B[55] +
//             mat_A[194] * mat_B[87] +
//             mat_A[195] * mat_B[119] +
//             mat_A[196] * mat_B[151] +
//             mat_A[197] * mat_B[183] +
//             mat_A[198] * mat_B[215] +
//             mat_A[199] * mat_B[247] +
//             mat_A[200] * mat_B[279] +
//             mat_A[201] * mat_B[311] +
//             mat_A[202] * mat_B[343] +
//             mat_A[203] * mat_B[375] +
//             mat_A[204] * mat_B[407] +
//             mat_A[205] * mat_B[439] +
//             mat_A[206] * mat_B[471] +
//             mat_A[207] * mat_B[503] +
//             mat_A[208] * mat_B[535] +
//             mat_A[209] * mat_B[567] +
//             mat_A[210] * mat_B[599] +
//             mat_A[211] * mat_B[631] +
//             mat_A[212] * mat_B[663] +
//             mat_A[213] * mat_B[695] +
//             mat_A[214] * mat_B[727] +
//             mat_A[215] * mat_B[759] +
//             mat_A[216] * mat_B[791] +
//             mat_A[217] * mat_B[823] +
//             mat_A[218] * mat_B[855] +
//             mat_A[219] * mat_B[887] +
//             mat_A[220] * mat_B[919] +
//             mat_A[221] * mat_B[951] +
//             mat_A[222] * mat_B[983] +
//             mat_A[223] * mat_B[1015];
//  mat_C[216] <= 
//             mat_A[192] * mat_B[24] +
//             mat_A[193] * mat_B[56] +
//             mat_A[194] * mat_B[88] +
//             mat_A[195] * mat_B[120] +
//             mat_A[196] * mat_B[152] +
//             mat_A[197] * mat_B[184] +
//             mat_A[198] * mat_B[216] +
//             mat_A[199] * mat_B[248] +
//             mat_A[200] * mat_B[280] +
//             mat_A[201] * mat_B[312] +
//             mat_A[202] * mat_B[344] +
//             mat_A[203] * mat_B[376] +
//             mat_A[204] * mat_B[408] +
//             mat_A[205] * mat_B[440] +
//             mat_A[206] * mat_B[472] +
//             mat_A[207] * mat_B[504] +
//             mat_A[208] * mat_B[536] +
//             mat_A[209] * mat_B[568] +
//             mat_A[210] * mat_B[600] +
//             mat_A[211] * mat_B[632] +
//             mat_A[212] * mat_B[664] +
//             mat_A[213] * mat_B[696] +
//             mat_A[214] * mat_B[728] +
//             mat_A[215] * mat_B[760] +
//             mat_A[216] * mat_B[792] +
//             mat_A[217] * mat_B[824] +
//             mat_A[218] * mat_B[856] +
//             mat_A[219] * mat_B[888] +
//             mat_A[220] * mat_B[920] +
//             mat_A[221] * mat_B[952] +
//             mat_A[222] * mat_B[984] +
//             mat_A[223] * mat_B[1016];
//  mat_C[217] <= 
//             mat_A[192] * mat_B[25] +
//             mat_A[193] * mat_B[57] +
//             mat_A[194] * mat_B[89] +
//             mat_A[195] * mat_B[121] +
//             mat_A[196] * mat_B[153] +
//             mat_A[197] * mat_B[185] +
//             mat_A[198] * mat_B[217] +
//             mat_A[199] * mat_B[249] +
//             mat_A[200] * mat_B[281] +
//             mat_A[201] * mat_B[313] +
//             mat_A[202] * mat_B[345] +
//             mat_A[203] * mat_B[377] +
//             mat_A[204] * mat_B[409] +
//             mat_A[205] * mat_B[441] +
//             mat_A[206] * mat_B[473] +
//             mat_A[207] * mat_B[505] +
//             mat_A[208] * mat_B[537] +
//             mat_A[209] * mat_B[569] +
//             mat_A[210] * mat_B[601] +
//             mat_A[211] * mat_B[633] +
//             mat_A[212] * mat_B[665] +
//             mat_A[213] * mat_B[697] +
//             mat_A[214] * mat_B[729] +
//             mat_A[215] * mat_B[761] +
//             mat_A[216] * mat_B[793] +
//             mat_A[217] * mat_B[825] +
//             mat_A[218] * mat_B[857] +
//             mat_A[219] * mat_B[889] +
//             mat_A[220] * mat_B[921] +
//             mat_A[221] * mat_B[953] +
//             mat_A[222] * mat_B[985] +
//             mat_A[223] * mat_B[1017];
//  mat_C[218] <= 
//             mat_A[192] * mat_B[26] +
//             mat_A[193] * mat_B[58] +
//             mat_A[194] * mat_B[90] +
//             mat_A[195] * mat_B[122] +
//             mat_A[196] * mat_B[154] +
//             mat_A[197] * mat_B[186] +
//             mat_A[198] * mat_B[218] +
//             mat_A[199] * mat_B[250] +
//             mat_A[200] * mat_B[282] +
//             mat_A[201] * mat_B[314] +
//             mat_A[202] * mat_B[346] +
//             mat_A[203] * mat_B[378] +
//             mat_A[204] * mat_B[410] +
//             mat_A[205] * mat_B[442] +
//             mat_A[206] * mat_B[474] +
//             mat_A[207] * mat_B[506] +
//             mat_A[208] * mat_B[538] +
//             mat_A[209] * mat_B[570] +
//             mat_A[210] * mat_B[602] +
//             mat_A[211] * mat_B[634] +
//             mat_A[212] * mat_B[666] +
//             mat_A[213] * mat_B[698] +
//             mat_A[214] * mat_B[730] +
//             mat_A[215] * mat_B[762] +
//             mat_A[216] * mat_B[794] +
//             mat_A[217] * mat_B[826] +
//             mat_A[218] * mat_B[858] +
//             mat_A[219] * mat_B[890] +
//             mat_A[220] * mat_B[922] +
//             mat_A[221] * mat_B[954] +
//             mat_A[222] * mat_B[986] +
//             mat_A[223] * mat_B[1018];
//  mat_C[219] <= 
//             mat_A[192] * mat_B[27] +
//             mat_A[193] * mat_B[59] +
//             mat_A[194] * mat_B[91] +
//             mat_A[195] * mat_B[123] +
//             mat_A[196] * mat_B[155] +
//             mat_A[197] * mat_B[187] +
//             mat_A[198] * mat_B[219] +
//             mat_A[199] * mat_B[251] +
//             mat_A[200] * mat_B[283] +
//             mat_A[201] * mat_B[315] +
//             mat_A[202] * mat_B[347] +
//             mat_A[203] * mat_B[379] +
//             mat_A[204] * mat_B[411] +
//             mat_A[205] * mat_B[443] +
//             mat_A[206] * mat_B[475] +
//             mat_A[207] * mat_B[507] +
//             mat_A[208] * mat_B[539] +
//             mat_A[209] * mat_B[571] +
//             mat_A[210] * mat_B[603] +
//             mat_A[211] * mat_B[635] +
//             mat_A[212] * mat_B[667] +
//             mat_A[213] * mat_B[699] +
//             mat_A[214] * mat_B[731] +
//             mat_A[215] * mat_B[763] +
//             mat_A[216] * mat_B[795] +
//             mat_A[217] * mat_B[827] +
//             mat_A[218] * mat_B[859] +
//             mat_A[219] * mat_B[891] +
//             mat_A[220] * mat_B[923] +
//             mat_A[221] * mat_B[955] +
//             mat_A[222] * mat_B[987] +
//             mat_A[223] * mat_B[1019];
//  mat_C[220] <= 
//             mat_A[192] * mat_B[28] +
//             mat_A[193] * mat_B[60] +
//             mat_A[194] * mat_B[92] +
//             mat_A[195] * mat_B[124] +
//             mat_A[196] * mat_B[156] +
//             mat_A[197] * mat_B[188] +
//             mat_A[198] * mat_B[220] +
//             mat_A[199] * mat_B[252] +
//             mat_A[200] * mat_B[284] +
//             mat_A[201] * mat_B[316] +
//             mat_A[202] * mat_B[348] +
//             mat_A[203] * mat_B[380] +
//             mat_A[204] * mat_B[412] +
//             mat_A[205] * mat_B[444] +
//             mat_A[206] * mat_B[476] +
//             mat_A[207] * mat_B[508] +
//             mat_A[208] * mat_B[540] +
//             mat_A[209] * mat_B[572] +
//             mat_A[210] * mat_B[604] +
//             mat_A[211] * mat_B[636] +
//             mat_A[212] * mat_B[668] +
//             mat_A[213] * mat_B[700] +
//             mat_A[214] * mat_B[732] +
//             mat_A[215] * mat_B[764] +
//             mat_A[216] * mat_B[796] +
//             mat_A[217] * mat_B[828] +
//             mat_A[218] * mat_B[860] +
//             mat_A[219] * mat_B[892] +
//             mat_A[220] * mat_B[924] +
//             mat_A[221] * mat_B[956] +
//             mat_A[222] * mat_B[988] +
//             mat_A[223] * mat_B[1020];
//  mat_C[221] <= 
//             mat_A[192] * mat_B[29] +
//             mat_A[193] * mat_B[61] +
//             mat_A[194] * mat_B[93] +
//             mat_A[195] * mat_B[125] +
//             mat_A[196] * mat_B[157] +
//             mat_A[197] * mat_B[189] +
//             mat_A[198] * mat_B[221] +
//             mat_A[199] * mat_B[253] +
//             mat_A[200] * mat_B[285] +
//             mat_A[201] * mat_B[317] +
//             mat_A[202] * mat_B[349] +
//             mat_A[203] * mat_B[381] +
//             mat_A[204] * mat_B[413] +
//             mat_A[205] * mat_B[445] +
//             mat_A[206] * mat_B[477] +
//             mat_A[207] * mat_B[509] +
//             mat_A[208] * mat_B[541] +
//             mat_A[209] * mat_B[573] +
//             mat_A[210] * mat_B[605] +
//             mat_A[211] * mat_B[637] +
//             mat_A[212] * mat_B[669] +
//             mat_A[213] * mat_B[701] +
//             mat_A[214] * mat_B[733] +
//             mat_A[215] * mat_B[765] +
//             mat_A[216] * mat_B[797] +
//             mat_A[217] * mat_B[829] +
//             mat_A[218] * mat_B[861] +
//             mat_A[219] * mat_B[893] +
//             mat_A[220] * mat_B[925] +
//             mat_A[221] * mat_B[957] +
//             mat_A[222] * mat_B[989] +
//             mat_A[223] * mat_B[1021];
//  mat_C[222] <= 
//             mat_A[192] * mat_B[30] +
//             mat_A[193] * mat_B[62] +
//             mat_A[194] * mat_B[94] +
//             mat_A[195] * mat_B[126] +
//             mat_A[196] * mat_B[158] +
//             mat_A[197] * mat_B[190] +
//             mat_A[198] * mat_B[222] +
//             mat_A[199] * mat_B[254] +
//             mat_A[200] * mat_B[286] +
//             mat_A[201] * mat_B[318] +
//             mat_A[202] * mat_B[350] +
//             mat_A[203] * mat_B[382] +
//             mat_A[204] * mat_B[414] +
//             mat_A[205] * mat_B[446] +
//             mat_A[206] * mat_B[478] +
//             mat_A[207] * mat_B[510] +
//             mat_A[208] * mat_B[542] +
//             mat_A[209] * mat_B[574] +
//             mat_A[210] * mat_B[606] +
//             mat_A[211] * mat_B[638] +
//             mat_A[212] * mat_B[670] +
//             mat_A[213] * mat_B[702] +
//             mat_A[214] * mat_B[734] +
//             mat_A[215] * mat_B[766] +
//             mat_A[216] * mat_B[798] +
//             mat_A[217] * mat_B[830] +
//             mat_A[218] * mat_B[862] +
//             mat_A[219] * mat_B[894] +
//             mat_A[220] * mat_B[926] +
//             mat_A[221] * mat_B[958] +
//             mat_A[222] * mat_B[990] +
//             mat_A[223] * mat_B[1022];
//  mat_C[223] <= 
//             mat_A[192] * mat_B[31] +
//             mat_A[193] * mat_B[63] +
//             mat_A[194] * mat_B[95] +
//             mat_A[195] * mat_B[127] +
//             mat_A[196] * mat_B[159] +
//             mat_A[197] * mat_B[191] +
//             mat_A[198] * mat_B[223] +
//             mat_A[199] * mat_B[255] +
//             mat_A[200] * mat_B[287] +
//             mat_A[201] * mat_B[319] +
//             mat_A[202] * mat_B[351] +
//             mat_A[203] * mat_B[383] +
//             mat_A[204] * mat_B[415] +
//             mat_A[205] * mat_B[447] +
//             mat_A[206] * mat_B[479] +
//             mat_A[207] * mat_B[511] +
//             mat_A[208] * mat_B[543] +
//             mat_A[209] * mat_B[575] +
//             mat_A[210] * mat_B[607] +
//             mat_A[211] * mat_B[639] +
//             mat_A[212] * mat_B[671] +
//             mat_A[213] * mat_B[703] +
//             mat_A[214] * mat_B[735] +
//             mat_A[215] * mat_B[767] +
//             mat_A[216] * mat_B[799] +
//             mat_A[217] * mat_B[831] +
//             mat_A[218] * mat_B[863] +
//             mat_A[219] * mat_B[895] +
//             mat_A[220] * mat_B[927] +
//             mat_A[221] * mat_B[959] +
//             mat_A[222] * mat_B[991] +
//             mat_A[223] * mat_B[1023];
//  mat_C[224] <= 
//             mat_A[224] * mat_B[0] +
//             mat_A[225] * mat_B[32] +
//             mat_A[226] * mat_B[64] +
//             mat_A[227] * mat_B[96] +
//             mat_A[228] * mat_B[128] +
//             mat_A[229] * mat_B[160] +
//             mat_A[230] * mat_B[192] +
//             mat_A[231] * mat_B[224] +
//             mat_A[232] * mat_B[256] +
//             mat_A[233] * mat_B[288] +
//             mat_A[234] * mat_B[320] +
//             mat_A[235] * mat_B[352] +
//             mat_A[236] * mat_B[384] +
//             mat_A[237] * mat_B[416] +
//             mat_A[238] * mat_B[448] +
//             mat_A[239] * mat_B[480] +
//             mat_A[240] * mat_B[512] +
//             mat_A[241] * mat_B[544] +
//             mat_A[242] * mat_B[576] +
//             mat_A[243] * mat_B[608] +
//             mat_A[244] * mat_B[640] +
//             mat_A[245] * mat_B[672] +
//             mat_A[246] * mat_B[704] +
//             mat_A[247] * mat_B[736] +
//             mat_A[248] * mat_B[768] +
//             mat_A[249] * mat_B[800] +
//             mat_A[250] * mat_B[832] +
//             mat_A[251] * mat_B[864] +
//             mat_A[252] * mat_B[896] +
//             mat_A[253] * mat_B[928] +
//             mat_A[254] * mat_B[960] +
//             mat_A[255] * mat_B[992];
//  mat_C[225] <= 
//             mat_A[224] * mat_B[1] +
//             mat_A[225] * mat_B[33] +
//             mat_A[226] * mat_B[65] +
//             mat_A[227] * mat_B[97] +
//             mat_A[228] * mat_B[129] +
//             mat_A[229] * mat_B[161] +
//             mat_A[230] * mat_B[193] +
//             mat_A[231] * mat_B[225] +
//             mat_A[232] * mat_B[257] +
//             mat_A[233] * mat_B[289] +
//             mat_A[234] * mat_B[321] +
//             mat_A[235] * mat_B[353] +
//             mat_A[236] * mat_B[385] +
//             mat_A[237] * mat_B[417] +
//             mat_A[238] * mat_B[449] +
//             mat_A[239] * mat_B[481] +
//             mat_A[240] * mat_B[513] +
//             mat_A[241] * mat_B[545] +
//             mat_A[242] * mat_B[577] +
//             mat_A[243] * mat_B[609] +
//             mat_A[244] * mat_B[641] +
//             mat_A[245] * mat_B[673] +
//             mat_A[246] * mat_B[705] +
//             mat_A[247] * mat_B[737] +
//             mat_A[248] * mat_B[769] +
//             mat_A[249] * mat_B[801] +
//             mat_A[250] * mat_B[833] +
//             mat_A[251] * mat_B[865] +
//             mat_A[252] * mat_B[897] +
//             mat_A[253] * mat_B[929] +
//             mat_A[254] * mat_B[961] +
//             mat_A[255] * mat_B[993];
//  mat_C[226] <= 
//             mat_A[224] * mat_B[2] +
//             mat_A[225] * mat_B[34] +
//             mat_A[226] * mat_B[66] +
//             mat_A[227] * mat_B[98] +
//             mat_A[228] * mat_B[130] +
//             mat_A[229] * mat_B[162] +
//             mat_A[230] * mat_B[194] +
//             mat_A[231] * mat_B[226] +
//             mat_A[232] * mat_B[258] +
//             mat_A[233] * mat_B[290] +
//             mat_A[234] * mat_B[322] +
//             mat_A[235] * mat_B[354] +
//             mat_A[236] * mat_B[386] +
//             mat_A[237] * mat_B[418] +
//             mat_A[238] * mat_B[450] +
//             mat_A[239] * mat_B[482] +
//             mat_A[240] * mat_B[514] +
//             mat_A[241] * mat_B[546] +
//             mat_A[242] * mat_B[578] +
//             mat_A[243] * mat_B[610] +
//             mat_A[244] * mat_B[642] +
//             mat_A[245] * mat_B[674] +
//             mat_A[246] * mat_B[706] +
//             mat_A[247] * mat_B[738] +
//             mat_A[248] * mat_B[770] +
//             mat_A[249] * mat_B[802] +
//             mat_A[250] * mat_B[834] +
//             mat_A[251] * mat_B[866] +
//             mat_A[252] * mat_B[898] +
//             mat_A[253] * mat_B[930] +
//             mat_A[254] * mat_B[962] +
//             mat_A[255] * mat_B[994];
//  mat_C[227] <= 
//             mat_A[224] * mat_B[3] +
//             mat_A[225] * mat_B[35] +
//             mat_A[226] * mat_B[67] +
//             mat_A[227] * mat_B[99] +
//             mat_A[228] * mat_B[131] +
//             mat_A[229] * mat_B[163] +
//             mat_A[230] * mat_B[195] +
//             mat_A[231] * mat_B[227] +
//             mat_A[232] * mat_B[259] +
//             mat_A[233] * mat_B[291] +
//             mat_A[234] * mat_B[323] +
//             mat_A[235] * mat_B[355] +
//             mat_A[236] * mat_B[387] +
//             mat_A[237] * mat_B[419] +
//             mat_A[238] * mat_B[451] +
//             mat_A[239] * mat_B[483] +
//             mat_A[240] * mat_B[515] +
//             mat_A[241] * mat_B[547] +
//             mat_A[242] * mat_B[579] +
//             mat_A[243] * mat_B[611] +
//             mat_A[244] * mat_B[643] +
//             mat_A[245] * mat_B[675] +
//             mat_A[246] * mat_B[707] +
//             mat_A[247] * mat_B[739] +
//             mat_A[248] * mat_B[771] +
//             mat_A[249] * mat_B[803] +
//             mat_A[250] * mat_B[835] +
//             mat_A[251] * mat_B[867] +
//             mat_A[252] * mat_B[899] +
//             mat_A[253] * mat_B[931] +
//             mat_A[254] * mat_B[963] +
//             mat_A[255] * mat_B[995];
//  mat_C[228] <= 
//             mat_A[224] * mat_B[4] +
//             mat_A[225] * mat_B[36] +
//             mat_A[226] * mat_B[68] +
//             mat_A[227] * mat_B[100] +
//             mat_A[228] * mat_B[132] +
//             mat_A[229] * mat_B[164] +
//             mat_A[230] * mat_B[196] +
//             mat_A[231] * mat_B[228] +
//             mat_A[232] * mat_B[260] +
//             mat_A[233] * mat_B[292] +
//             mat_A[234] * mat_B[324] +
//             mat_A[235] * mat_B[356] +
//             mat_A[236] * mat_B[388] +
//             mat_A[237] * mat_B[420] +
//             mat_A[238] * mat_B[452] +
//             mat_A[239] * mat_B[484] +
//             mat_A[240] * mat_B[516] +
//             mat_A[241] * mat_B[548] +
//             mat_A[242] * mat_B[580] +
//             mat_A[243] * mat_B[612] +
//             mat_A[244] * mat_B[644] +
//             mat_A[245] * mat_B[676] +
//             mat_A[246] * mat_B[708] +
//             mat_A[247] * mat_B[740] +
//             mat_A[248] * mat_B[772] +
//             mat_A[249] * mat_B[804] +
//             mat_A[250] * mat_B[836] +
//             mat_A[251] * mat_B[868] +
//             mat_A[252] * mat_B[900] +
//             mat_A[253] * mat_B[932] +
//             mat_A[254] * mat_B[964] +
//             mat_A[255] * mat_B[996];
//  mat_C[229] <= 
//             mat_A[224] * mat_B[5] +
//             mat_A[225] * mat_B[37] +
//             mat_A[226] * mat_B[69] +
//             mat_A[227] * mat_B[101] +
//             mat_A[228] * mat_B[133] +
//             mat_A[229] * mat_B[165] +
//             mat_A[230] * mat_B[197] +
//             mat_A[231] * mat_B[229] +
//             mat_A[232] * mat_B[261] +
//             mat_A[233] * mat_B[293] +
//             mat_A[234] * mat_B[325] +
//             mat_A[235] * mat_B[357] +
//             mat_A[236] * mat_B[389] +
//             mat_A[237] * mat_B[421] +
//             mat_A[238] * mat_B[453] +
//             mat_A[239] * mat_B[485] +
//             mat_A[240] * mat_B[517] +
//             mat_A[241] * mat_B[549] +
//             mat_A[242] * mat_B[581] +
//             mat_A[243] * mat_B[613] +
//             mat_A[244] * mat_B[645] +
//             mat_A[245] * mat_B[677] +
//             mat_A[246] * mat_B[709] +
//             mat_A[247] * mat_B[741] +
//             mat_A[248] * mat_B[773] +
//             mat_A[249] * mat_B[805] +
//             mat_A[250] * mat_B[837] +
//             mat_A[251] * mat_B[869] +
//             mat_A[252] * mat_B[901] +
//             mat_A[253] * mat_B[933] +
//             mat_A[254] * mat_B[965] +
//             mat_A[255] * mat_B[997];
//  mat_C[230] <= 
//             mat_A[224] * mat_B[6] +
//             mat_A[225] * mat_B[38] +
//             mat_A[226] * mat_B[70] +
//             mat_A[227] * mat_B[102] +
//             mat_A[228] * mat_B[134] +
//             mat_A[229] * mat_B[166] +
//             mat_A[230] * mat_B[198] +
//             mat_A[231] * mat_B[230] +
//             mat_A[232] * mat_B[262] +
//             mat_A[233] * mat_B[294] +
//             mat_A[234] * mat_B[326] +
//             mat_A[235] * mat_B[358] +
//             mat_A[236] * mat_B[390] +
//             mat_A[237] * mat_B[422] +
//             mat_A[238] * mat_B[454] +
//             mat_A[239] * mat_B[486] +
//             mat_A[240] * mat_B[518] +
//             mat_A[241] * mat_B[550] +
//             mat_A[242] * mat_B[582] +
//             mat_A[243] * mat_B[614] +
//             mat_A[244] * mat_B[646] +
//             mat_A[245] * mat_B[678] +
//             mat_A[246] * mat_B[710] +
//             mat_A[247] * mat_B[742] +
//             mat_A[248] * mat_B[774] +
//             mat_A[249] * mat_B[806] +
//             mat_A[250] * mat_B[838] +
//             mat_A[251] * mat_B[870] +
//             mat_A[252] * mat_B[902] +
//             mat_A[253] * mat_B[934] +
//             mat_A[254] * mat_B[966] +
//             mat_A[255] * mat_B[998];
//  mat_C[231] <= 
//             mat_A[224] * mat_B[7] +
//             mat_A[225] * mat_B[39] +
//             mat_A[226] * mat_B[71] +
//             mat_A[227] * mat_B[103] +
//             mat_A[228] * mat_B[135] +
//             mat_A[229] * mat_B[167] +
//             mat_A[230] * mat_B[199] +
//             mat_A[231] * mat_B[231] +
//             mat_A[232] * mat_B[263] +
//             mat_A[233] * mat_B[295] +
//             mat_A[234] * mat_B[327] +
//             mat_A[235] * mat_B[359] +
//             mat_A[236] * mat_B[391] +
//             mat_A[237] * mat_B[423] +
//             mat_A[238] * mat_B[455] +
//             mat_A[239] * mat_B[487] +
//             mat_A[240] * mat_B[519] +
//             mat_A[241] * mat_B[551] +
//             mat_A[242] * mat_B[583] +
//             mat_A[243] * mat_B[615] +
//             mat_A[244] * mat_B[647] +
//             mat_A[245] * mat_B[679] +
//             mat_A[246] * mat_B[711] +
//             mat_A[247] * mat_B[743] +
//             mat_A[248] * mat_B[775] +
//             mat_A[249] * mat_B[807] +
//             mat_A[250] * mat_B[839] +
//             mat_A[251] * mat_B[871] +
//             mat_A[252] * mat_B[903] +
//             mat_A[253] * mat_B[935] +
//             mat_A[254] * mat_B[967] +
//             mat_A[255] * mat_B[999];
//  mat_C[232] <= 
//             mat_A[224] * mat_B[8] +
//             mat_A[225] * mat_B[40] +
//             mat_A[226] * mat_B[72] +
//             mat_A[227] * mat_B[104] +
//             mat_A[228] * mat_B[136] +
//             mat_A[229] * mat_B[168] +
//             mat_A[230] * mat_B[200] +
//             mat_A[231] * mat_B[232] +
//             mat_A[232] * mat_B[264] +
//             mat_A[233] * mat_B[296] +
//             mat_A[234] * mat_B[328] +
//             mat_A[235] * mat_B[360] +
//             mat_A[236] * mat_B[392] +
//             mat_A[237] * mat_B[424] +
//             mat_A[238] * mat_B[456] +
//             mat_A[239] * mat_B[488] +
//             mat_A[240] * mat_B[520] +
//             mat_A[241] * mat_B[552] +
//             mat_A[242] * mat_B[584] +
//             mat_A[243] * mat_B[616] +
//             mat_A[244] * mat_B[648] +
//             mat_A[245] * mat_B[680] +
//             mat_A[246] * mat_B[712] +
//             mat_A[247] * mat_B[744] +
//             mat_A[248] * mat_B[776] +
//             mat_A[249] * mat_B[808] +
//             mat_A[250] * mat_B[840] +
//             mat_A[251] * mat_B[872] +
//             mat_A[252] * mat_B[904] +
//             mat_A[253] * mat_B[936] +
//             mat_A[254] * mat_B[968] +
//             mat_A[255] * mat_B[1000];
//  mat_C[233] <= 
//             mat_A[224] * mat_B[9] +
//             mat_A[225] * mat_B[41] +
//             mat_A[226] * mat_B[73] +
//             mat_A[227] * mat_B[105] +
//             mat_A[228] * mat_B[137] +
//             mat_A[229] * mat_B[169] +
//             mat_A[230] * mat_B[201] +
//             mat_A[231] * mat_B[233] +
//             mat_A[232] * mat_B[265] +
//             mat_A[233] * mat_B[297] +
//             mat_A[234] * mat_B[329] +
//             mat_A[235] * mat_B[361] +
//             mat_A[236] * mat_B[393] +
//             mat_A[237] * mat_B[425] +
//             mat_A[238] * mat_B[457] +
//             mat_A[239] * mat_B[489] +
//             mat_A[240] * mat_B[521] +
//             mat_A[241] * mat_B[553] +
//             mat_A[242] * mat_B[585] +
//             mat_A[243] * mat_B[617] +
//             mat_A[244] * mat_B[649] +
//             mat_A[245] * mat_B[681] +
//             mat_A[246] * mat_B[713] +
//             mat_A[247] * mat_B[745] +
//             mat_A[248] * mat_B[777] +
//             mat_A[249] * mat_B[809] +
//             mat_A[250] * mat_B[841] +
//             mat_A[251] * mat_B[873] +
//             mat_A[252] * mat_B[905] +
//             mat_A[253] * mat_B[937] +
//             mat_A[254] * mat_B[969] +
//             mat_A[255] * mat_B[1001];
//  mat_C[234] <= 
//             mat_A[224] * mat_B[10] +
//             mat_A[225] * mat_B[42] +
//             mat_A[226] * mat_B[74] +
//             mat_A[227] * mat_B[106] +
//             mat_A[228] * mat_B[138] +
//             mat_A[229] * mat_B[170] +
//             mat_A[230] * mat_B[202] +
//             mat_A[231] * mat_B[234] +
//             mat_A[232] * mat_B[266] +
//             mat_A[233] * mat_B[298] +
//             mat_A[234] * mat_B[330] +
//             mat_A[235] * mat_B[362] +
//             mat_A[236] * mat_B[394] +
//             mat_A[237] * mat_B[426] +
//             mat_A[238] * mat_B[458] +
//             mat_A[239] * mat_B[490] +
//             mat_A[240] * mat_B[522] +
//             mat_A[241] * mat_B[554] +
//             mat_A[242] * mat_B[586] +
//             mat_A[243] * mat_B[618] +
//             mat_A[244] * mat_B[650] +
//             mat_A[245] * mat_B[682] +
//             mat_A[246] * mat_B[714] +
//             mat_A[247] * mat_B[746] +
//             mat_A[248] * mat_B[778] +
//             mat_A[249] * mat_B[810] +
//             mat_A[250] * mat_B[842] +
//             mat_A[251] * mat_B[874] +
//             mat_A[252] * mat_B[906] +
//             mat_A[253] * mat_B[938] +
//             mat_A[254] * mat_B[970] +
//             mat_A[255] * mat_B[1002];
//  mat_C[235] <= 
//             mat_A[224] * mat_B[11] +
//             mat_A[225] * mat_B[43] +
//             mat_A[226] * mat_B[75] +
//             mat_A[227] * mat_B[107] +
//             mat_A[228] * mat_B[139] +
//             mat_A[229] * mat_B[171] +
//             mat_A[230] * mat_B[203] +
//             mat_A[231] * mat_B[235] +
//             mat_A[232] * mat_B[267] +
//             mat_A[233] * mat_B[299] +
//             mat_A[234] * mat_B[331] +
//             mat_A[235] * mat_B[363] +
//             mat_A[236] * mat_B[395] +
//             mat_A[237] * mat_B[427] +
//             mat_A[238] * mat_B[459] +
//             mat_A[239] * mat_B[491] +
//             mat_A[240] * mat_B[523] +
//             mat_A[241] * mat_B[555] +
//             mat_A[242] * mat_B[587] +
//             mat_A[243] * mat_B[619] +
//             mat_A[244] * mat_B[651] +
//             mat_A[245] * mat_B[683] +
//             mat_A[246] * mat_B[715] +
//             mat_A[247] * mat_B[747] +
//             mat_A[248] * mat_B[779] +
//             mat_A[249] * mat_B[811] +
//             mat_A[250] * mat_B[843] +
//             mat_A[251] * mat_B[875] +
//             mat_A[252] * mat_B[907] +
//             mat_A[253] * mat_B[939] +
//             mat_A[254] * mat_B[971] +
//             mat_A[255] * mat_B[1003];
//  mat_C[236] <= 
//             mat_A[224] * mat_B[12] +
//             mat_A[225] * mat_B[44] +
//             mat_A[226] * mat_B[76] +
//             mat_A[227] * mat_B[108] +
//             mat_A[228] * mat_B[140] +
//             mat_A[229] * mat_B[172] +
//             mat_A[230] * mat_B[204] +
//             mat_A[231] * mat_B[236] +
//             mat_A[232] * mat_B[268] +
//             mat_A[233] * mat_B[300] +
//             mat_A[234] * mat_B[332] +
//             mat_A[235] * mat_B[364] +
//             mat_A[236] * mat_B[396] +
//             mat_A[237] * mat_B[428] +
//             mat_A[238] * mat_B[460] +
//             mat_A[239] * mat_B[492] +
//             mat_A[240] * mat_B[524] +
//             mat_A[241] * mat_B[556] +
//             mat_A[242] * mat_B[588] +
//             mat_A[243] * mat_B[620] +
//             mat_A[244] * mat_B[652] +
//             mat_A[245] * mat_B[684] +
//             mat_A[246] * mat_B[716] +
//             mat_A[247] * mat_B[748] +
//             mat_A[248] * mat_B[780] +
//             mat_A[249] * mat_B[812] +
//             mat_A[250] * mat_B[844] +
//             mat_A[251] * mat_B[876] +
//             mat_A[252] * mat_B[908] +
//             mat_A[253] * mat_B[940] +
//             mat_A[254] * mat_B[972] +
//             mat_A[255] * mat_B[1004];
//  mat_C[237] <= 
//             mat_A[224] * mat_B[13] +
//             mat_A[225] * mat_B[45] +
//             mat_A[226] * mat_B[77] +
//             mat_A[227] * mat_B[109] +
//             mat_A[228] * mat_B[141] +
//             mat_A[229] * mat_B[173] +
//             mat_A[230] * mat_B[205] +
//             mat_A[231] * mat_B[237] +
//             mat_A[232] * mat_B[269] +
//             mat_A[233] * mat_B[301] +
//             mat_A[234] * mat_B[333] +
//             mat_A[235] * mat_B[365] +
//             mat_A[236] * mat_B[397] +
//             mat_A[237] * mat_B[429] +
//             mat_A[238] * mat_B[461] +
//             mat_A[239] * mat_B[493] +
//             mat_A[240] * mat_B[525] +
//             mat_A[241] * mat_B[557] +
//             mat_A[242] * mat_B[589] +
//             mat_A[243] * mat_B[621] +
//             mat_A[244] * mat_B[653] +
//             mat_A[245] * mat_B[685] +
//             mat_A[246] * mat_B[717] +
//             mat_A[247] * mat_B[749] +
//             mat_A[248] * mat_B[781] +
//             mat_A[249] * mat_B[813] +
//             mat_A[250] * mat_B[845] +
//             mat_A[251] * mat_B[877] +
//             mat_A[252] * mat_B[909] +
//             mat_A[253] * mat_B[941] +
//             mat_A[254] * mat_B[973] +
//             mat_A[255] * mat_B[1005];
//  mat_C[238] <= 
//             mat_A[224] * mat_B[14] +
//             mat_A[225] * mat_B[46] +
//             mat_A[226] * mat_B[78] +
//             mat_A[227] * mat_B[110] +
//             mat_A[228] * mat_B[142] +
//             mat_A[229] * mat_B[174] +
//             mat_A[230] * mat_B[206] +
//             mat_A[231] * mat_B[238] +
//             mat_A[232] * mat_B[270] +
//             mat_A[233] * mat_B[302] +
//             mat_A[234] * mat_B[334] +
//             mat_A[235] * mat_B[366] +
//             mat_A[236] * mat_B[398] +
//             mat_A[237] * mat_B[430] +
//             mat_A[238] * mat_B[462] +
//             mat_A[239] * mat_B[494] +
//             mat_A[240] * mat_B[526] +
//             mat_A[241] * mat_B[558] +
//             mat_A[242] * mat_B[590] +
//             mat_A[243] * mat_B[622] +
//             mat_A[244] * mat_B[654] +
//             mat_A[245] * mat_B[686] +
//             mat_A[246] * mat_B[718] +
//             mat_A[247] * mat_B[750] +
//             mat_A[248] * mat_B[782] +
//             mat_A[249] * mat_B[814] +
//             mat_A[250] * mat_B[846] +
//             mat_A[251] * mat_B[878] +
//             mat_A[252] * mat_B[910] +
//             mat_A[253] * mat_B[942] +
//             mat_A[254] * mat_B[974] +
//             mat_A[255] * mat_B[1006];
//  mat_C[239] <= 
//             mat_A[224] * mat_B[15] +
//             mat_A[225] * mat_B[47] +
//             mat_A[226] * mat_B[79] +
//             mat_A[227] * mat_B[111] +
//             mat_A[228] * mat_B[143] +
//             mat_A[229] * mat_B[175] +
//             mat_A[230] * mat_B[207] +
//             mat_A[231] * mat_B[239] +
//             mat_A[232] * mat_B[271] +
//             mat_A[233] * mat_B[303] +
//             mat_A[234] * mat_B[335] +
//             mat_A[235] * mat_B[367] +
//             mat_A[236] * mat_B[399] +
//             mat_A[237] * mat_B[431] +
//             mat_A[238] * mat_B[463] +
//             mat_A[239] * mat_B[495] +
//             mat_A[240] * mat_B[527] +
//             mat_A[241] * mat_B[559] +
//             mat_A[242] * mat_B[591] +
//             mat_A[243] * mat_B[623] +
//             mat_A[244] * mat_B[655] +
//             mat_A[245] * mat_B[687] +
//             mat_A[246] * mat_B[719] +
//             mat_A[247] * mat_B[751] +
//             mat_A[248] * mat_B[783] +
//             mat_A[249] * mat_B[815] +
//             mat_A[250] * mat_B[847] +
//             mat_A[251] * mat_B[879] +
//             mat_A[252] * mat_B[911] +
//             mat_A[253] * mat_B[943] +
//             mat_A[254] * mat_B[975] +
//             mat_A[255] * mat_B[1007];
//  mat_C[240] <= 
//             mat_A[224] * mat_B[16] +
//             mat_A[225] * mat_B[48] +
//             mat_A[226] * mat_B[80] +
//             mat_A[227] * mat_B[112] +
//             mat_A[228] * mat_B[144] +
//             mat_A[229] * mat_B[176] +
//             mat_A[230] * mat_B[208] +
//             mat_A[231] * mat_B[240] +
//             mat_A[232] * mat_B[272] +
//             mat_A[233] * mat_B[304] +
//             mat_A[234] * mat_B[336] +
//             mat_A[235] * mat_B[368] +
//             mat_A[236] * mat_B[400] +
//             mat_A[237] * mat_B[432] +
//             mat_A[238] * mat_B[464] +
//             mat_A[239] * mat_B[496] +
//             mat_A[240] * mat_B[528] +
//             mat_A[241] * mat_B[560] +
//             mat_A[242] * mat_B[592] +
//             mat_A[243] * mat_B[624] +
//             mat_A[244] * mat_B[656] +
//             mat_A[245] * mat_B[688] +
//             mat_A[246] * mat_B[720] +
//             mat_A[247] * mat_B[752] +
//             mat_A[248] * mat_B[784] +
//             mat_A[249] * mat_B[816] +
//             mat_A[250] * mat_B[848] +
//             mat_A[251] * mat_B[880] +
//             mat_A[252] * mat_B[912] +
//             mat_A[253] * mat_B[944] +
//             mat_A[254] * mat_B[976] +
//             mat_A[255] * mat_B[1008];
//  mat_C[241] <= 
//             mat_A[224] * mat_B[17] +
//             mat_A[225] * mat_B[49] +
//             mat_A[226] * mat_B[81] +
//             mat_A[227] * mat_B[113] +
//             mat_A[228] * mat_B[145] +
//             mat_A[229] * mat_B[177] +
//             mat_A[230] * mat_B[209] +
//             mat_A[231] * mat_B[241] +
//             mat_A[232] * mat_B[273] +
//             mat_A[233] * mat_B[305] +
//             mat_A[234] * mat_B[337] +
//             mat_A[235] * mat_B[369] +
//             mat_A[236] * mat_B[401] +
//             mat_A[237] * mat_B[433] +
//             mat_A[238] * mat_B[465] +
//             mat_A[239] * mat_B[497] +
//             mat_A[240] * mat_B[529] +
//             mat_A[241] * mat_B[561] +
//             mat_A[242] * mat_B[593] +
//             mat_A[243] * mat_B[625] +
//             mat_A[244] * mat_B[657] +
//             mat_A[245] * mat_B[689] +
//             mat_A[246] * mat_B[721] +
//             mat_A[247] * mat_B[753] +
//             mat_A[248] * mat_B[785] +
//             mat_A[249] * mat_B[817] +
//             mat_A[250] * mat_B[849] +
//             mat_A[251] * mat_B[881] +
//             mat_A[252] * mat_B[913] +
//             mat_A[253] * mat_B[945] +
//             mat_A[254] * mat_B[977] +
//             mat_A[255] * mat_B[1009];
//  mat_C[242] <= 
//             mat_A[224] * mat_B[18] +
//             mat_A[225] * mat_B[50] +
//             mat_A[226] * mat_B[82] +
//             mat_A[227] * mat_B[114] +
//             mat_A[228] * mat_B[146] +
//             mat_A[229] * mat_B[178] +
//             mat_A[230] * mat_B[210] +
//             mat_A[231] * mat_B[242] +
//             mat_A[232] * mat_B[274] +
//             mat_A[233] * mat_B[306] +
//             mat_A[234] * mat_B[338] +
//             mat_A[235] * mat_B[370] +
//             mat_A[236] * mat_B[402] +
//             mat_A[237] * mat_B[434] +
//             mat_A[238] * mat_B[466] +
//             mat_A[239] * mat_B[498] +
//             mat_A[240] * mat_B[530] +
//             mat_A[241] * mat_B[562] +
//             mat_A[242] * mat_B[594] +
//             mat_A[243] * mat_B[626] +
//             mat_A[244] * mat_B[658] +
//             mat_A[245] * mat_B[690] +
//             mat_A[246] * mat_B[722] +
//             mat_A[247] * mat_B[754] +
//             mat_A[248] * mat_B[786] +
//             mat_A[249] * mat_B[818] +
//             mat_A[250] * mat_B[850] +
//             mat_A[251] * mat_B[882] +
//             mat_A[252] * mat_B[914] +
//             mat_A[253] * mat_B[946] +
//             mat_A[254] * mat_B[978] +
//             mat_A[255] * mat_B[1010];
//  mat_C[243] <= 
//             mat_A[224] * mat_B[19] +
//             mat_A[225] * mat_B[51] +
//             mat_A[226] * mat_B[83] +
//             mat_A[227] * mat_B[115] +
//             mat_A[228] * mat_B[147] +
//             mat_A[229] * mat_B[179] +
//             mat_A[230] * mat_B[211] +
//             mat_A[231] * mat_B[243] +
//             mat_A[232] * mat_B[275] +
//             mat_A[233] * mat_B[307] +
//             mat_A[234] * mat_B[339] +
//             mat_A[235] * mat_B[371] +
//             mat_A[236] * mat_B[403] +
//             mat_A[237] * mat_B[435] +
//             mat_A[238] * mat_B[467] +
//             mat_A[239] * mat_B[499] +
//             mat_A[240] * mat_B[531] +
//             mat_A[241] * mat_B[563] +
//             mat_A[242] * mat_B[595] +
//             mat_A[243] * mat_B[627] +
//             mat_A[244] * mat_B[659] +
//             mat_A[245] * mat_B[691] +
//             mat_A[246] * mat_B[723] +
//             mat_A[247] * mat_B[755] +
//             mat_A[248] * mat_B[787] +
//             mat_A[249] * mat_B[819] +
//             mat_A[250] * mat_B[851] +
//             mat_A[251] * mat_B[883] +
//             mat_A[252] * mat_B[915] +
//             mat_A[253] * mat_B[947] +
//             mat_A[254] * mat_B[979] +
//             mat_A[255] * mat_B[1011];
//  mat_C[244] <= 
//             mat_A[224] * mat_B[20] +
//             mat_A[225] * mat_B[52] +
//             mat_A[226] * mat_B[84] +
//             mat_A[227] * mat_B[116] +
//             mat_A[228] * mat_B[148] +
//             mat_A[229] * mat_B[180] +
//             mat_A[230] * mat_B[212] +
//             mat_A[231] * mat_B[244] +
//             mat_A[232] * mat_B[276] +
//             mat_A[233] * mat_B[308] +
//             mat_A[234] * mat_B[340] +
//             mat_A[235] * mat_B[372] +
//             mat_A[236] * mat_B[404] +
//             mat_A[237] * mat_B[436] +
//             mat_A[238] * mat_B[468] +
//             mat_A[239] * mat_B[500] +
//             mat_A[240] * mat_B[532] +
//             mat_A[241] * mat_B[564] +
//             mat_A[242] * mat_B[596] +
//             mat_A[243] * mat_B[628] +
//             mat_A[244] * mat_B[660] +
//             mat_A[245] * mat_B[692] +
//             mat_A[246] * mat_B[724] +
//             mat_A[247] * mat_B[756] +
//             mat_A[248] * mat_B[788] +
//             mat_A[249] * mat_B[820] +
//             mat_A[250] * mat_B[852] +
//             mat_A[251] * mat_B[884] +
//             mat_A[252] * mat_B[916] +
//             mat_A[253] * mat_B[948] +
//             mat_A[254] * mat_B[980] +
//             mat_A[255] * mat_B[1012];
//  mat_C[245] <= 
//             mat_A[224] * mat_B[21] +
//             mat_A[225] * mat_B[53] +
//             mat_A[226] * mat_B[85] +
//             mat_A[227] * mat_B[117] +
//             mat_A[228] * mat_B[149] +
//             mat_A[229] * mat_B[181] +
//             mat_A[230] * mat_B[213] +
//             mat_A[231] * mat_B[245] +
//             mat_A[232] * mat_B[277] +
//             mat_A[233] * mat_B[309] +
//             mat_A[234] * mat_B[341] +
//             mat_A[235] * mat_B[373] +
//             mat_A[236] * mat_B[405] +
//             mat_A[237] * mat_B[437] +
//             mat_A[238] * mat_B[469] +
//             mat_A[239] * mat_B[501] +
//             mat_A[240] * mat_B[533] +
//             mat_A[241] * mat_B[565] +
//             mat_A[242] * mat_B[597] +
//             mat_A[243] * mat_B[629] +
//             mat_A[244] * mat_B[661] +
//             mat_A[245] * mat_B[693] +
//             mat_A[246] * mat_B[725] +
//             mat_A[247] * mat_B[757] +
//             mat_A[248] * mat_B[789] +
//             mat_A[249] * mat_B[821] +
//             mat_A[250] * mat_B[853] +
//             mat_A[251] * mat_B[885] +
//             mat_A[252] * mat_B[917] +
//             mat_A[253] * mat_B[949] +
//             mat_A[254] * mat_B[981] +
//             mat_A[255] * mat_B[1013];
//  mat_C[246] <= 
//             mat_A[224] * mat_B[22] +
//             mat_A[225] * mat_B[54] +
//             mat_A[226] * mat_B[86] +
//             mat_A[227] * mat_B[118] +
//             mat_A[228] * mat_B[150] +
//             mat_A[229] * mat_B[182] +
//             mat_A[230] * mat_B[214] +
//             mat_A[231] * mat_B[246] +
//             mat_A[232] * mat_B[278] +
//             mat_A[233] * mat_B[310] +
//             mat_A[234] * mat_B[342] +
//             mat_A[235] * mat_B[374] +
//             mat_A[236] * mat_B[406] +
//             mat_A[237] * mat_B[438] +
//             mat_A[238] * mat_B[470] +
//             mat_A[239] * mat_B[502] +
//             mat_A[240] * mat_B[534] +
//             mat_A[241] * mat_B[566] +
//             mat_A[242] * mat_B[598] +
//             mat_A[243] * mat_B[630] +
//             mat_A[244] * mat_B[662] +
//             mat_A[245] * mat_B[694] +
//             mat_A[246] * mat_B[726] +
//             mat_A[247] * mat_B[758] +
//             mat_A[248] * mat_B[790] +
//             mat_A[249] * mat_B[822] +
//             mat_A[250] * mat_B[854] +
//             mat_A[251] * mat_B[886] +
//             mat_A[252] * mat_B[918] +
//             mat_A[253] * mat_B[950] +
//             mat_A[254] * mat_B[982] +
//             mat_A[255] * mat_B[1014];
//  mat_C[247] <= 
//             mat_A[224] * mat_B[23] +
//             mat_A[225] * mat_B[55] +
//             mat_A[226] * mat_B[87] +
//             mat_A[227] * mat_B[119] +
//             mat_A[228] * mat_B[151] +
//             mat_A[229] * mat_B[183] +
//             mat_A[230] * mat_B[215] +
//             mat_A[231] * mat_B[247] +
//             mat_A[232] * mat_B[279] +
//             mat_A[233] * mat_B[311] +
//             mat_A[234] * mat_B[343] +
//             mat_A[235] * mat_B[375] +
//             mat_A[236] * mat_B[407] +
//             mat_A[237] * mat_B[439] +
//             mat_A[238] * mat_B[471] +
//             mat_A[239] * mat_B[503] +
//             mat_A[240] * mat_B[535] +
//             mat_A[241] * mat_B[567] +
//             mat_A[242] * mat_B[599] +
//             mat_A[243] * mat_B[631] +
//             mat_A[244] * mat_B[663] +
//             mat_A[245] * mat_B[695] +
//             mat_A[246] * mat_B[727] +
//             mat_A[247] * mat_B[759] +
//             mat_A[248] * mat_B[791] +
//             mat_A[249] * mat_B[823] +
//             mat_A[250] * mat_B[855] +
//             mat_A[251] * mat_B[887] +
//             mat_A[252] * mat_B[919] +
//             mat_A[253] * mat_B[951] +
//             mat_A[254] * mat_B[983] +
//             mat_A[255] * mat_B[1015];
//  mat_C[248] <= 
//             mat_A[224] * mat_B[24] +
//             mat_A[225] * mat_B[56] +
//             mat_A[226] * mat_B[88] +
//             mat_A[227] * mat_B[120] +
//             mat_A[228] * mat_B[152] +
//             mat_A[229] * mat_B[184] +
//             mat_A[230] * mat_B[216] +
//             mat_A[231] * mat_B[248] +
//             mat_A[232] * mat_B[280] +
//             mat_A[233] * mat_B[312] +
//             mat_A[234] * mat_B[344] +
//             mat_A[235] * mat_B[376] +
//             mat_A[236] * mat_B[408] +
//             mat_A[237] * mat_B[440] +
//             mat_A[238] * mat_B[472] +
//             mat_A[239] * mat_B[504] +
//             mat_A[240] * mat_B[536] +
//             mat_A[241] * mat_B[568] +
//             mat_A[242] * mat_B[600] +
//             mat_A[243] * mat_B[632] +
//             mat_A[244] * mat_B[664] +
//             mat_A[245] * mat_B[696] +
//             mat_A[246] * mat_B[728] +
//             mat_A[247] * mat_B[760] +
//             mat_A[248] * mat_B[792] +
//             mat_A[249] * mat_B[824] +
//             mat_A[250] * mat_B[856] +
//             mat_A[251] * mat_B[888] +
//             mat_A[252] * mat_B[920] +
//             mat_A[253] * mat_B[952] +
//             mat_A[254] * mat_B[984] +
//             mat_A[255] * mat_B[1016];
//  mat_C[249] <= 
//             mat_A[224] * mat_B[25] +
//             mat_A[225] * mat_B[57] +
//             mat_A[226] * mat_B[89] +
//             mat_A[227] * mat_B[121] +
//             mat_A[228] * mat_B[153] +
//             mat_A[229] * mat_B[185] +
//             mat_A[230] * mat_B[217] +
//             mat_A[231] * mat_B[249] +
//             mat_A[232] * mat_B[281] +
//             mat_A[233] * mat_B[313] +
//             mat_A[234] * mat_B[345] +
//             mat_A[235] * mat_B[377] +
//             mat_A[236] * mat_B[409] +
//             mat_A[237] * mat_B[441] +
//             mat_A[238] * mat_B[473] +
//             mat_A[239] * mat_B[505] +
//             mat_A[240] * mat_B[537] +
//             mat_A[241] * mat_B[569] +
//             mat_A[242] * mat_B[601] +
//             mat_A[243] * mat_B[633] +
//             mat_A[244] * mat_B[665] +
//             mat_A[245] * mat_B[697] +
//             mat_A[246] * mat_B[729] +
//             mat_A[247] * mat_B[761] +
//             mat_A[248] * mat_B[793] +
//             mat_A[249] * mat_B[825] +
//             mat_A[250] * mat_B[857] +
//             mat_A[251] * mat_B[889] +
//             mat_A[252] * mat_B[921] +
//             mat_A[253] * mat_B[953] +
//             mat_A[254] * mat_B[985] +
//             mat_A[255] * mat_B[1017];
//  mat_C[250] <= 
//             mat_A[224] * mat_B[26] +
//             mat_A[225] * mat_B[58] +
//             mat_A[226] * mat_B[90] +
//             mat_A[227] * mat_B[122] +
//             mat_A[228] * mat_B[154] +
//             mat_A[229] * mat_B[186] +
//             mat_A[230] * mat_B[218] +
//             mat_A[231] * mat_B[250] +
//             mat_A[232] * mat_B[282] +
//             mat_A[233] * mat_B[314] +
//             mat_A[234] * mat_B[346] +
//             mat_A[235] * mat_B[378] +
//             mat_A[236] * mat_B[410] +
//             mat_A[237] * mat_B[442] +
//             mat_A[238] * mat_B[474] +
//             mat_A[239] * mat_B[506] +
//             mat_A[240] * mat_B[538] +
//             mat_A[241] * mat_B[570] +
//             mat_A[242] * mat_B[602] +
//             mat_A[243] * mat_B[634] +
//             mat_A[244] * mat_B[666] +
//             mat_A[245] * mat_B[698] +
//             mat_A[246] * mat_B[730] +
//             mat_A[247] * mat_B[762] +
//             mat_A[248] * mat_B[794] +
//             mat_A[249] * mat_B[826] +
//             mat_A[250] * mat_B[858] +
//             mat_A[251] * mat_B[890] +
//             mat_A[252] * mat_B[922] +
//             mat_A[253] * mat_B[954] +
//             mat_A[254] * mat_B[986] +
//             mat_A[255] * mat_B[1018];
//  mat_C[251] <= 
//             mat_A[224] * mat_B[27] +
//             mat_A[225] * mat_B[59] +
//             mat_A[226] * mat_B[91] +
//             mat_A[227] * mat_B[123] +
//             mat_A[228] * mat_B[155] +
//             mat_A[229] * mat_B[187] +
//             mat_A[230] * mat_B[219] +
//             mat_A[231] * mat_B[251] +
//             mat_A[232] * mat_B[283] +
//             mat_A[233] * mat_B[315] +
//             mat_A[234] * mat_B[347] +
//             mat_A[235] * mat_B[379] +
//             mat_A[236] * mat_B[411] +
//             mat_A[237] * mat_B[443] +
//             mat_A[238] * mat_B[475] +
//             mat_A[239] * mat_B[507] +
//             mat_A[240] * mat_B[539] +
//             mat_A[241] * mat_B[571] +
//             mat_A[242] * mat_B[603] +
//             mat_A[243] * mat_B[635] +
//             mat_A[244] * mat_B[667] +
//             mat_A[245] * mat_B[699] +
//             mat_A[246] * mat_B[731] +
//             mat_A[247] * mat_B[763] +
//             mat_A[248] * mat_B[795] +
//             mat_A[249] * mat_B[827] +
//             mat_A[250] * mat_B[859] +
//             mat_A[251] * mat_B[891] +
//             mat_A[252] * mat_B[923] +
//             mat_A[253] * mat_B[955] +
//             mat_A[254] * mat_B[987] +
//             mat_A[255] * mat_B[1019];
//  mat_C[252] <= 
//             mat_A[224] * mat_B[28] +
//             mat_A[225] * mat_B[60] +
//             mat_A[226] * mat_B[92] +
//             mat_A[227] * mat_B[124] +
//             mat_A[228] * mat_B[156] +
//             mat_A[229] * mat_B[188] +
//             mat_A[230] * mat_B[220] +
//             mat_A[231] * mat_B[252] +
//             mat_A[232] * mat_B[284] +
//             mat_A[233] * mat_B[316] +
//             mat_A[234] * mat_B[348] +
//             mat_A[235] * mat_B[380] +
//             mat_A[236] * mat_B[412] +
//             mat_A[237] * mat_B[444] +
//             mat_A[238] * mat_B[476] +
//             mat_A[239] * mat_B[508] +
//             mat_A[240] * mat_B[540] +
//             mat_A[241] * mat_B[572] +
//             mat_A[242] * mat_B[604] +
//             mat_A[243] * mat_B[636] +
//             mat_A[244] * mat_B[668] +
//             mat_A[245] * mat_B[700] +
//             mat_A[246] * mat_B[732] +
//             mat_A[247] * mat_B[764] +
//             mat_A[248] * mat_B[796] +
//             mat_A[249] * mat_B[828] +
//             mat_A[250] * mat_B[860] +
//             mat_A[251] * mat_B[892] +
//             mat_A[252] * mat_B[924] +
//             mat_A[253] * mat_B[956] +
//             mat_A[254] * mat_B[988] +
//             mat_A[255] * mat_B[1020];
//  mat_C[253] <= 
//             mat_A[224] * mat_B[29] +
//             mat_A[225] * mat_B[61] +
//             mat_A[226] * mat_B[93] +
//             mat_A[227] * mat_B[125] +
//             mat_A[228] * mat_B[157] +
//             mat_A[229] * mat_B[189] +
//             mat_A[230] * mat_B[221] +
//             mat_A[231] * mat_B[253] +
//             mat_A[232] * mat_B[285] +
//             mat_A[233] * mat_B[317] +
//             mat_A[234] * mat_B[349] +
//             mat_A[235] * mat_B[381] +
//             mat_A[236] * mat_B[413] +
//             mat_A[237] * mat_B[445] +
//             mat_A[238] * mat_B[477] +
//             mat_A[239] * mat_B[509] +
//             mat_A[240] * mat_B[541] +
//             mat_A[241] * mat_B[573] +
//             mat_A[242] * mat_B[605] +
//             mat_A[243] * mat_B[637] +
//             mat_A[244] * mat_B[669] +
//             mat_A[245] * mat_B[701] +
//             mat_A[246] * mat_B[733] +
//             mat_A[247] * mat_B[765] +
//             mat_A[248] * mat_B[797] +
//             mat_A[249] * mat_B[829] +
//             mat_A[250] * mat_B[861] +
//             mat_A[251] * mat_B[893] +
//             mat_A[252] * mat_B[925] +
//             mat_A[253] * mat_B[957] +
//             mat_A[254] * mat_B[989] +
//             mat_A[255] * mat_B[1021];
//  mat_C[254] <= 
//             mat_A[224] * mat_B[30] +
//             mat_A[225] * mat_B[62] +
//             mat_A[226] * mat_B[94] +
//             mat_A[227] * mat_B[126] +
//             mat_A[228] * mat_B[158] +
//             mat_A[229] * mat_B[190] +
//             mat_A[230] * mat_B[222] +
//             mat_A[231] * mat_B[254] +
//             mat_A[232] * mat_B[286] +
//             mat_A[233] * mat_B[318] +
//             mat_A[234] * mat_B[350] +
//             mat_A[235] * mat_B[382] +
//             mat_A[236] * mat_B[414] +
//             mat_A[237] * mat_B[446] +
//             mat_A[238] * mat_B[478] +
//             mat_A[239] * mat_B[510] +
//             mat_A[240] * mat_B[542] +
//             mat_A[241] * mat_B[574] +
//             mat_A[242] * mat_B[606] +
//             mat_A[243] * mat_B[638] +
//             mat_A[244] * mat_B[670] +
//             mat_A[245] * mat_B[702] +
//             mat_A[246] * mat_B[734] +
//             mat_A[247] * mat_B[766] +
//             mat_A[248] * mat_B[798] +
//             mat_A[249] * mat_B[830] +
//             mat_A[250] * mat_B[862] +
//             mat_A[251] * mat_B[894] +
//             mat_A[252] * mat_B[926] +
//             mat_A[253] * mat_B[958] +
//             mat_A[254] * mat_B[990] +
//             mat_A[255] * mat_B[1022];
//  mat_C[255] <= 
//             mat_A[224] * mat_B[31] +
//             mat_A[225] * mat_B[63] +
//             mat_A[226] * mat_B[95] +
//             mat_A[227] * mat_B[127] +
//             mat_A[228] * mat_B[159] +
//             mat_A[229] * mat_B[191] +
//             mat_A[230] * mat_B[223] +
//             mat_A[231] * mat_B[255] +
//             mat_A[232] * mat_B[287] +
//             mat_A[233] * mat_B[319] +
//             mat_A[234] * mat_B[351] +
//             mat_A[235] * mat_B[383] +
//             mat_A[236] * mat_B[415] +
//             mat_A[237] * mat_B[447] +
//             mat_A[238] * mat_B[479] +
//             mat_A[239] * mat_B[511] +
//             mat_A[240] * mat_B[543] +
//             mat_A[241] * mat_B[575] +
//             mat_A[242] * mat_B[607] +
//             mat_A[243] * mat_B[639] +
//             mat_A[244] * mat_B[671] +
//             mat_A[245] * mat_B[703] +
//             mat_A[246] * mat_B[735] +
//             mat_A[247] * mat_B[767] +
//             mat_A[248] * mat_B[799] +
//             mat_A[249] * mat_B[831] +
//             mat_A[250] * mat_B[863] +
//             mat_A[251] * mat_B[895] +
//             mat_A[252] * mat_B[927] +
//             mat_A[253] * mat_B[959] +
//             mat_A[254] * mat_B[991] +
//             mat_A[255] * mat_B[1023];
//  mat_C[256] <= 
//             mat_A[256] * mat_B[0] +
//             mat_A[257] * mat_B[32] +
//             mat_A[258] * mat_B[64] +
//             mat_A[259] * mat_B[96] +
//             mat_A[260] * mat_B[128] +
//             mat_A[261] * mat_B[160] +
//             mat_A[262] * mat_B[192] +
//             mat_A[263] * mat_B[224] +
//             mat_A[264] * mat_B[256] +
//             mat_A[265] * mat_B[288] +
//             mat_A[266] * mat_B[320] +
//             mat_A[267] * mat_B[352] +
//             mat_A[268] * mat_B[384] +
//             mat_A[269] * mat_B[416] +
//             mat_A[270] * mat_B[448] +
//             mat_A[271] * mat_B[480] +
//             mat_A[272] * mat_B[512] +
//             mat_A[273] * mat_B[544] +
//             mat_A[274] * mat_B[576] +
//             mat_A[275] * mat_B[608] +
//             mat_A[276] * mat_B[640] +
//             mat_A[277] * mat_B[672] +
//             mat_A[278] * mat_B[704] +
//             mat_A[279] * mat_B[736] +
//             mat_A[280] * mat_B[768] +
//             mat_A[281] * mat_B[800] +
//             mat_A[282] * mat_B[832] +
//             mat_A[283] * mat_B[864] +
//             mat_A[284] * mat_B[896] +
//             mat_A[285] * mat_B[928] +
//             mat_A[286] * mat_B[960] +
//             mat_A[287] * mat_B[992];
//  mat_C[257] <= 
//             mat_A[256] * mat_B[1] +
//             mat_A[257] * mat_B[33] +
//             mat_A[258] * mat_B[65] +
//             mat_A[259] * mat_B[97] +
//             mat_A[260] * mat_B[129] +
//             mat_A[261] * mat_B[161] +
//             mat_A[262] * mat_B[193] +
//             mat_A[263] * mat_B[225] +
//             mat_A[264] * mat_B[257] +
//             mat_A[265] * mat_B[289] +
//             mat_A[266] * mat_B[321] +
//             mat_A[267] * mat_B[353] +
//             mat_A[268] * mat_B[385] +
//             mat_A[269] * mat_B[417] +
//             mat_A[270] * mat_B[449] +
//             mat_A[271] * mat_B[481] +
//             mat_A[272] * mat_B[513] +
//             mat_A[273] * mat_B[545] +
//             mat_A[274] * mat_B[577] +
//             mat_A[275] * mat_B[609] +
//             mat_A[276] * mat_B[641] +
//             mat_A[277] * mat_B[673] +
//             mat_A[278] * mat_B[705] +
//             mat_A[279] * mat_B[737] +
//             mat_A[280] * mat_B[769] +
//             mat_A[281] * mat_B[801] +
//             mat_A[282] * mat_B[833] +
//             mat_A[283] * mat_B[865] +
//             mat_A[284] * mat_B[897] +
//             mat_A[285] * mat_B[929] +
//             mat_A[286] * mat_B[961] +
//             mat_A[287] * mat_B[993];
//  mat_C[258] <= 
//             mat_A[256] * mat_B[2] +
//             mat_A[257] * mat_B[34] +
//             mat_A[258] * mat_B[66] +
//             mat_A[259] * mat_B[98] +
//             mat_A[260] * mat_B[130] +
//             mat_A[261] * mat_B[162] +
//             mat_A[262] * mat_B[194] +
//             mat_A[263] * mat_B[226] +
//             mat_A[264] * mat_B[258] +
//             mat_A[265] * mat_B[290] +
//             mat_A[266] * mat_B[322] +
//             mat_A[267] * mat_B[354] +
//             mat_A[268] * mat_B[386] +
//             mat_A[269] * mat_B[418] +
//             mat_A[270] * mat_B[450] +
//             mat_A[271] * mat_B[482] +
//             mat_A[272] * mat_B[514] +
//             mat_A[273] * mat_B[546] +
//             mat_A[274] * mat_B[578] +
//             mat_A[275] * mat_B[610] +
//             mat_A[276] * mat_B[642] +
//             mat_A[277] * mat_B[674] +
//             mat_A[278] * mat_B[706] +
//             mat_A[279] * mat_B[738] +
//             mat_A[280] * mat_B[770] +
//             mat_A[281] * mat_B[802] +
//             mat_A[282] * mat_B[834] +
//             mat_A[283] * mat_B[866] +
//             mat_A[284] * mat_B[898] +
//             mat_A[285] * mat_B[930] +
//             mat_A[286] * mat_B[962] +
//             mat_A[287] * mat_B[994];
//  mat_C[259] <= 
//             mat_A[256] * mat_B[3] +
//             mat_A[257] * mat_B[35] +
//             mat_A[258] * mat_B[67] +
//             mat_A[259] * mat_B[99] +
//             mat_A[260] * mat_B[131] +
//             mat_A[261] * mat_B[163] +
//             mat_A[262] * mat_B[195] +
//             mat_A[263] * mat_B[227] +
//             mat_A[264] * mat_B[259] +
//             mat_A[265] * mat_B[291] +
//             mat_A[266] * mat_B[323] +
//             mat_A[267] * mat_B[355] +
//             mat_A[268] * mat_B[387] +
//             mat_A[269] * mat_B[419] +
//             mat_A[270] * mat_B[451] +
//             mat_A[271] * mat_B[483] +
//             mat_A[272] * mat_B[515] +
//             mat_A[273] * mat_B[547] +
//             mat_A[274] * mat_B[579] +
//             mat_A[275] * mat_B[611] +
//             mat_A[276] * mat_B[643] +
//             mat_A[277] * mat_B[675] +
//             mat_A[278] * mat_B[707] +
//             mat_A[279] * mat_B[739] +
//             mat_A[280] * mat_B[771] +
//             mat_A[281] * mat_B[803] +
//             mat_A[282] * mat_B[835] +
//             mat_A[283] * mat_B[867] +
//             mat_A[284] * mat_B[899] +
//             mat_A[285] * mat_B[931] +
//             mat_A[286] * mat_B[963] +
//             mat_A[287] * mat_B[995];
//  mat_C[260] <= 
//             mat_A[256] * mat_B[4] +
//             mat_A[257] * mat_B[36] +
//             mat_A[258] * mat_B[68] +
//             mat_A[259] * mat_B[100] +
//             mat_A[260] * mat_B[132] +
//             mat_A[261] * mat_B[164] +
//             mat_A[262] * mat_B[196] +
//             mat_A[263] * mat_B[228] +
//             mat_A[264] * mat_B[260] +
//             mat_A[265] * mat_B[292] +
//             mat_A[266] * mat_B[324] +
//             mat_A[267] * mat_B[356] +
//             mat_A[268] * mat_B[388] +
//             mat_A[269] * mat_B[420] +
//             mat_A[270] * mat_B[452] +
//             mat_A[271] * mat_B[484] +
//             mat_A[272] * mat_B[516] +
//             mat_A[273] * mat_B[548] +
//             mat_A[274] * mat_B[580] +
//             mat_A[275] * mat_B[612] +
//             mat_A[276] * mat_B[644] +
//             mat_A[277] * mat_B[676] +
//             mat_A[278] * mat_B[708] +
//             mat_A[279] * mat_B[740] +
//             mat_A[280] * mat_B[772] +
//             mat_A[281] * mat_B[804] +
//             mat_A[282] * mat_B[836] +
//             mat_A[283] * mat_B[868] +
//             mat_A[284] * mat_B[900] +
//             mat_A[285] * mat_B[932] +
//             mat_A[286] * mat_B[964] +
//             mat_A[287] * mat_B[996];
//  mat_C[261] <= 
//             mat_A[256] * mat_B[5] +
//             mat_A[257] * mat_B[37] +
//             mat_A[258] * mat_B[69] +
//             mat_A[259] * mat_B[101] +
//             mat_A[260] * mat_B[133] +
//             mat_A[261] * mat_B[165] +
//             mat_A[262] * mat_B[197] +
//             mat_A[263] * mat_B[229] +
//             mat_A[264] * mat_B[261] +
//             mat_A[265] * mat_B[293] +
//             mat_A[266] * mat_B[325] +
//             mat_A[267] * mat_B[357] +
//             mat_A[268] * mat_B[389] +
//             mat_A[269] * mat_B[421] +
//             mat_A[270] * mat_B[453] +
//             mat_A[271] * mat_B[485] +
//             mat_A[272] * mat_B[517] +
//             mat_A[273] * mat_B[549] +
//             mat_A[274] * mat_B[581] +
//             mat_A[275] * mat_B[613] +
//             mat_A[276] * mat_B[645] +
//             mat_A[277] * mat_B[677] +
//             mat_A[278] * mat_B[709] +
//             mat_A[279] * mat_B[741] +
//             mat_A[280] * mat_B[773] +
//             mat_A[281] * mat_B[805] +
//             mat_A[282] * mat_B[837] +
//             mat_A[283] * mat_B[869] +
//             mat_A[284] * mat_B[901] +
//             mat_A[285] * mat_B[933] +
//             mat_A[286] * mat_B[965] +
//             mat_A[287] * mat_B[997];
//  mat_C[262] <= 
//             mat_A[256] * mat_B[6] +
//             mat_A[257] * mat_B[38] +
//             mat_A[258] * mat_B[70] +
//             mat_A[259] * mat_B[102] +
//             mat_A[260] * mat_B[134] +
//             mat_A[261] * mat_B[166] +
//             mat_A[262] * mat_B[198] +
//             mat_A[263] * mat_B[230] +
//             mat_A[264] * mat_B[262] +
//             mat_A[265] * mat_B[294] +
//             mat_A[266] * mat_B[326] +
//             mat_A[267] * mat_B[358] +
//             mat_A[268] * mat_B[390] +
//             mat_A[269] * mat_B[422] +
//             mat_A[270] * mat_B[454] +
//             mat_A[271] * mat_B[486] +
//             mat_A[272] * mat_B[518] +
//             mat_A[273] * mat_B[550] +
//             mat_A[274] * mat_B[582] +
//             mat_A[275] * mat_B[614] +
//             mat_A[276] * mat_B[646] +
//             mat_A[277] * mat_B[678] +
//             mat_A[278] * mat_B[710] +
//             mat_A[279] * mat_B[742] +
//             mat_A[280] * mat_B[774] +
//             mat_A[281] * mat_B[806] +
//             mat_A[282] * mat_B[838] +
//             mat_A[283] * mat_B[870] +
//             mat_A[284] * mat_B[902] +
//             mat_A[285] * mat_B[934] +
//             mat_A[286] * mat_B[966] +
//             mat_A[287] * mat_B[998];
//  mat_C[263] <= 
//             mat_A[256] * mat_B[7] +
//             mat_A[257] * mat_B[39] +
//             mat_A[258] * mat_B[71] +
//             mat_A[259] * mat_B[103] +
//             mat_A[260] * mat_B[135] +
//             mat_A[261] * mat_B[167] +
//             mat_A[262] * mat_B[199] +
//             mat_A[263] * mat_B[231] +
//             mat_A[264] * mat_B[263] +
//             mat_A[265] * mat_B[295] +
//             mat_A[266] * mat_B[327] +
//             mat_A[267] * mat_B[359] +
//             mat_A[268] * mat_B[391] +
//             mat_A[269] * mat_B[423] +
//             mat_A[270] * mat_B[455] +
//             mat_A[271] * mat_B[487] +
//             mat_A[272] * mat_B[519] +
//             mat_A[273] * mat_B[551] +
//             mat_A[274] * mat_B[583] +
//             mat_A[275] * mat_B[615] +
//             mat_A[276] * mat_B[647] +
//             mat_A[277] * mat_B[679] +
//             mat_A[278] * mat_B[711] +
//             mat_A[279] * mat_B[743] +
//             mat_A[280] * mat_B[775] +
//             mat_A[281] * mat_B[807] +
//             mat_A[282] * mat_B[839] +
//             mat_A[283] * mat_B[871] +
//             mat_A[284] * mat_B[903] +
//             mat_A[285] * mat_B[935] +
//             mat_A[286] * mat_B[967] +
//             mat_A[287] * mat_B[999];
//  mat_C[264] <= 
//             mat_A[256] * mat_B[8] +
//             mat_A[257] * mat_B[40] +
//             mat_A[258] * mat_B[72] +
//             mat_A[259] * mat_B[104] +
//             mat_A[260] * mat_B[136] +
//             mat_A[261] * mat_B[168] +
//             mat_A[262] * mat_B[200] +
//             mat_A[263] * mat_B[232] +
//             mat_A[264] * mat_B[264] +
//             mat_A[265] * mat_B[296] +
//             mat_A[266] * mat_B[328] +
//             mat_A[267] * mat_B[360] +
//             mat_A[268] * mat_B[392] +
//             mat_A[269] * mat_B[424] +
//             mat_A[270] * mat_B[456] +
//             mat_A[271] * mat_B[488] +
//             mat_A[272] * mat_B[520] +
//             mat_A[273] * mat_B[552] +
//             mat_A[274] * mat_B[584] +
//             mat_A[275] * mat_B[616] +
//             mat_A[276] * mat_B[648] +
//             mat_A[277] * mat_B[680] +
//             mat_A[278] * mat_B[712] +
//             mat_A[279] * mat_B[744] +
//             mat_A[280] * mat_B[776] +
//             mat_A[281] * mat_B[808] +
//             mat_A[282] * mat_B[840] +
//             mat_A[283] * mat_B[872] +
//             mat_A[284] * mat_B[904] +
//             mat_A[285] * mat_B[936] +
//             mat_A[286] * mat_B[968] +
//             mat_A[287] * mat_B[1000];
//  mat_C[265] <= 
//             mat_A[256] * mat_B[9] +
//             mat_A[257] * mat_B[41] +
//             mat_A[258] * mat_B[73] +
//             mat_A[259] * mat_B[105] +
//             mat_A[260] * mat_B[137] +
//             mat_A[261] * mat_B[169] +
//             mat_A[262] * mat_B[201] +
//             mat_A[263] * mat_B[233] +
//             mat_A[264] * mat_B[265] +
//             mat_A[265] * mat_B[297] +
//             mat_A[266] * mat_B[329] +
//             mat_A[267] * mat_B[361] +
//             mat_A[268] * mat_B[393] +
//             mat_A[269] * mat_B[425] +
//             mat_A[270] * mat_B[457] +
//             mat_A[271] * mat_B[489] +
//             mat_A[272] * mat_B[521] +
//             mat_A[273] * mat_B[553] +
//             mat_A[274] * mat_B[585] +
//             mat_A[275] * mat_B[617] +
//             mat_A[276] * mat_B[649] +
//             mat_A[277] * mat_B[681] +
//             mat_A[278] * mat_B[713] +
//             mat_A[279] * mat_B[745] +
//             mat_A[280] * mat_B[777] +
//             mat_A[281] * mat_B[809] +
//             mat_A[282] * mat_B[841] +
//             mat_A[283] * mat_B[873] +
//             mat_A[284] * mat_B[905] +
//             mat_A[285] * mat_B[937] +
//             mat_A[286] * mat_B[969] +
//             mat_A[287] * mat_B[1001];
//  mat_C[266] <= 
//             mat_A[256] * mat_B[10] +
//             mat_A[257] * mat_B[42] +
//             mat_A[258] * mat_B[74] +
//             mat_A[259] * mat_B[106] +
//             mat_A[260] * mat_B[138] +
//             mat_A[261] * mat_B[170] +
//             mat_A[262] * mat_B[202] +
//             mat_A[263] * mat_B[234] +
//             mat_A[264] * mat_B[266] +
//             mat_A[265] * mat_B[298] +
//             mat_A[266] * mat_B[330] +
//             mat_A[267] * mat_B[362] +
//             mat_A[268] * mat_B[394] +
//             mat_A[269] * mat_B[426] +
//             mat_A[270] * mat_B[458] +
//             mat_A[271] * mat_B[490] +
//             mat_A[272] * mat_B[522] +
//             mat_A[273] * mat_B[554] +
//             mat_A[274] * mat_B[586] +
//             mat_A[275] * mat_B[618] +
//             mat_A[276] * mat_B[650] +
//             mat_A[277] * mat_B[682] +
//             mat_A[278] * mat_B[714] +
//             mat_A[279] * mat_B[746] +
//             mat_A[280] * mat_B[778] +
//             mat_A[281] * mat_B[810] +
//             mat_A[282] * mat_B[842] +
//             mat_A[283] * mat_B[874] +
//             mat_A[284] * mat_B[906] +
//             mat_A[285] * mat_B[938] +
//             mat_A[286] * mat_B[970] +
//             mat_A[287] * mat_B[1002];
//  mat_C[267] <= 
//             mat_A[256] * mat_B[11] +
//             mat_A[257] * mat_B[43] +
//             mat_A[258] * mat_B[75] +
//             mat_A[259] * mat_B[107] +
//             mat_A[260] * mat_B[139] +
//             mat_A[261] * mat_B[171] +
//             mat_A[262] * mat_B[203] +
//             mat_A[263] * mat_B[235] +
//             mat_A[264] * mat_B[267] +
//             mat_A[265] * mat_B[299] +
//             mat_A[266] * mat_B[331] +
//             mat_A[267] * mat_B[363] +
//             mat_A[268] * mat_B[395] +
//             mat_A[269] * mat_B[427] +
//             mat_A[270] * mat_B[459] +
//             mat_A[271] * mat_B[491] +
//             mat_A[272] * mat_B[523] +
//             mat_A[273] * mat_B[555] +
//             mat_A[274] * mat_B[587] +
//             mat_A[275] * mat_B[619] +
//             mat_A[276] * mat_B[651] +
//             mat_A[277] * mat_B[683] +
//             mat_A[278] * mat_B[715] +
//             mat_A[279] * mat_B[747] +
//             mat_A[280] * mat_B[779] +
//             mat_A[281] * mat_B[811] +
//             mat_A[282] * mat_B[843] +
//             mat_A[283] * mat_B[875] +
//             mat_A[284] * mat_B[907] +
//             mat_A[285] * mat_B[939] +
//             mat_A[286] * mat_B[971] +
//             mat_A[287] * mat_B[1003];
//  mat_C[268] <= 
//             mat_A[256] * mat_B[12] +
//             mat_A[257] * mat_B[44] +
//             mat_A[258] * mat_B[76] +
//             mat_A[259] * mat_B[108] +
//             mat_A[260] * mat_B[140] +
//             mat_A[261] * mat_B[172] +
//             mat_A[262] * mat_B[204] +
//             mat_A[263] * mat_B[236] +
//             mat_A[264] * mat_B[268] +
//             mat_A[265] * mat_B[300] +
//             mat_A[266] * mat_B[332] +
//             mat_A[267] * mat_B[364] +
//             mat_A[268] * mat_B[396] +
//             mat_A[269] * mat_B[428] +
//             mat_A[270] * mat_B[460] +
//             mat_A[271] * mat_B[492] +
//             mat_A[272] * mat_B[524] +
//             mat_A[273] * mat_B[556] +
//             mat_A[274] * mat_B[588] +
//             mat_A[275] * mat_B[620] +
//             mat_A[276] * mat_B[652] +
//             mat_A[277] * mat_B[684] +
//             mat_A[278] * mat_B[716] +
//             mat_A[279] * mat_B[748] +
//             mat_A[280] * mat_B[780] +
//             mat_A[281] * mat_B[812] +
//             mat_A[282] * mat_B[844] +
//             mat_A[283] * mat_B[876] +
//             mat_A[284] * mat_B[908] +
//             mat_A[285] * mat_B[940] +
//             mat_A[286] * mat_B[972] +
//             mat_A[287] * mat_B[1004];
//  mat_C[269] <= 
//             mat_A[256] * mat_B[13] +
//             mat_A[257] * mat_B[45] +
//             mat_A[258] * mat_B[77] +
//             mat_A[259] * mat_B[109] +
//             mat_A[260] * mat_B[141] +
//             mat_A[261] * mat_B[173] +
//             mat_A[262] * mat_B[205] +
//             mat_A[263] * mat_B[237] +
//             mat_A[264] * mat_B[269] +
//             mat_A[265] * mat_B[301] +
//             mat_A[266] * mat_B[333] +
//             mat_A[267] * mat_B[365] +
//             mat_A[268] * mat_B[397] +
//             mat_A[269] * mat_B[429] +
//             mat_A[270] * mat_B[461] +
//             mat_A[271] * mat_B[493] +
//             mat_A[272] * mat_B[525] +
//             mat_A[273] * mat_B[557] +
//             mat_A[274] * mat_B[589] +
//             mat_A[275] * mat_B[621] +
//             mat_A[276] * mat_B[653] +
//             mat_A[277] * mat_B[685] +
//             mat_A[278] * mat_B[717] +
//             mat_A[279] * mat_B[749] +
//             mat_A[280] * mat_B[781] +
//             mat_A[281] * mat_B[813] +
//             mat_A[282] * mat_B[845] +
//             mat_A[283] * mat_B[877] +
//             mat_A[284] * mat_B[909] +
//             mat_A[285] * mat_B[941] +
//             mat_A[286] * mat_B[973] +
//             mat_A[287] * mat_B[1005];
//  mat_C[270] <= 
//             mat_A[256] * mat_B[14] +
//             mat_A[257] * mat_B[46] +
//             mat_A[258] * mat_B[78] +
//             mat_A[259] * mat_B[110] +
//             mat_A[260] * mat_B[142] +
//             mat_A[261] * mat_B[174] +
//             mat_A[262] * mat_B[206] +
//             mat_A[263] * mat_B[238] +
//             mat_A[264] * mat_B[270] +
//             mat_A[265] * mat_B[302] +
//             mat_A[266] * mat_B[334] +
//             mat_A[267] * mat_B[366] +
//             mat_A[268] * mat_B[398] +
//             mat_A[269] * mat_B[430] +
//             mat_A[270] * mat_B[462] +
//             mat_A[271] * mat_B[494] +
//             mat_A[272] * mat_B[526] +
//             mat_A[273] * mat_B[558] +
//             mat_A[274] * mat_B[590] +
//             mat_A[275] * mat_B[622] +
//             mat_A[276] * mat_B[654] +
//             mat_A[277] * mat_B[686] +
//             mat_A[278] * mat_B[718] +
//             mat_A[279] * mat_B[750] +
//             mat_A[280] * mat_B[782] +
//             mat_A[281] * mat_B[814] +
//             mat_A[282] * mat_B[846] +
//             mat_A[283] * mat_B[878] +
//             mat_A[284] * mat_B[910] +
//             mat_A[285] * mat_B[942] +
//             mat_A[286] * mat_B[974] +
//             mat_A[287] * mat_B[1006];
//  mat_C[271] <= 
//             mat_A[256] * mat_B[15] +
//             mat_A[257] * mat_B[47] +
//             mat_A[258] * mat_B[79] +
//             mat_A[259] * mat_B[111] +
//             mat_A[260] * mat_B[143] +
//             mat_A[261] * mat_B[175] +
//             mat_A[262] * mat_B[207] +
//             mat_A[263] * mat_B[239] +
//             mat_A[264] * mat_B[271] +
//             mat_A[265] * mat_B[303] +
//             mat_A[266] * mat_B[335] +
//             mat_A[267] * mat_B[367] +
//             mat_A[268] * mat_B[399] +
//             mat_A[269] * mat_B[431] +
//             mat_A[270] * mat_B[463] +
//             mat_A[271] * mat_B[495] +
//             mat_A[272] * mat_B[527] +
//             mat_A[273] * mat_B[559] +
//             mat_A[274] * mat_B[591] +
//             mat_A[275] * mat_B[623] +
//             mat_A[276] * mat_B[655] +
//             mat_A[277] * mat_B[687] +
//             mat_A[278] * mat_B[719] +
//             mat_A[279] * mat_B[751] +
//             mat_A[280] * mat_B[783] +
//             mat_A[281] * mat_B[815] +
//             mat_A[282] * mat_B[847] +
//             mat_A[283] * mat_B[879] +
//             mat_A[284] * mat_B[911] +
//             mat_A[285] * mat_B[943] +
//             mat_A[286] * mat_B[975] +
//             mat_A[287] * mat_B[1007];
//  mat_C[272] <= 
//             mat_A[256] * mat_B[16] +
//             mat_A[257] * mat_B[48] +
//             mat_A[258] * mat_B[80] +
//             mat_A[259] * mat_B[112] +
//             mat_A[260] * mat_B[144] +
//             mat_A[261] * mat_B[176] +
//             mat_A[262] * mat_B[208] +
//             mat_A[263] * mat_B[240] +
//             mat_A[264] * mat_B[272] +
//             mat_A[265] * mat_B[304] +
//             mat_A[266] * mat_B[336] +
//             mat_A[267] * mat_B[368] +
//             mat_A[268] * mat_B[400] +
//             mat_A[269] * mat_B[432] +
//             mat_A[270] * mat_B[464] +
//             mat_A[271] * mat_B[496] +
//             mat_A[272] * mat_B[528] +
//             mat_A[273] * mat_B[560] +
//             mat_A[274] * mat_B[592] +
//             mat_A[275] * mat_B[624] +
//             mat_A[276] * mat_B[656] +
//             mat_A[277] * mat_B[688] +
//             mat_A[278] * mat_B[720] +
//             mat_A[279] * mat_B[752] +
//             mat_A[280] * mat_B[784] +
//             mat_A[281] * mat_B[816] +
//             mat_A[282] * mat_B[848] +
//             mat_A[283] * mat_B[880] +
//             mat_A[284] * mat_B[912] +
//             mat_A[285] * mat_B[944] +
//             mat_A[286] * mat_B[976] +
//             mat_A[287] * mat_B[1008];
//  mat_C[273] <= 
//             mat_A[256] * mat_B[17] +
//             mat_A[257] * mat_B[49] +
//             mat_A[258] * mat_B[81] +
//             mat_A[259] * mat_B[113] +
//             mat_A[260] * mat_B[145] +
//             mat_A[261] * mat_B[177] +
//             mat_A[262] * mat_B[209] +
//             mat_A[263] * mat_B[241] +
//             mat_A[264] * mat_B[273] +
//             mat_A[265] * mat_B[305] +
//             mat_A[266] * mat_B[337] +
//             mat_A[267] * mat_B[369] +
//             mat_A[268] * mat_B[401] +
//             mat_A[269] * mat_B[433] +
//             mat_A[270] * mat_B[465] +
//             mat_A[271] * mat_B[497] +
//             mat_A[272] * mat_B[529] +
//             mat_A[273] * mat_B[561] +
//             mat_A[274] * mat_B[593] +
//             mat_A[275] * mat_B[625] +
//             mat_A[276] * mat_B[657] +
//             mat_A[277] * mat_B[689] +
//             mat_A[278] * mat_B[721] +
//             mat_A[279] * mat_B[753] +
//             mat_A[280] * mat_B[785] +
//             mat_A[281] * mat_B[817] +
//             mat_A[282] * mat_B[849] +
//             mat_A[283] * mat_B[881] +
//             mat_A[284] * mat_B[913] +
//             mat_A[285] * mat_B[945] +
//             mat_A[286] * mat_B[977] +
//             mat_A[287] * mat_B[1009];
//  mat_C[274] <= 
//             mat_A[256] * mat_B[18] +
//             mat_A[257] * mat_B[50] +
//             mat_A[258] * mat_B[82] +
//             mat_A[259] * mat_B[114] +
//             mat_A[260] * mat_B[146] +
//             mat_A[261] * mat_B[178] +
//             mat_A[262] * mat_B[210] +
//             mat_A[263] * mat_B[242] +
//             mat_A[264] * mat_B[274] +
//             mat_A[265] * mat_B[306] +
//             mat_A[266] * mat_B[338] +
//             mat_A[267] * mat_B[370] +
//             mat_A[268] * mat_B[402] +
//             mat_A[269] * mat_B[434] +
//             mat_A[270] * mat_B[466] +
//             mat_A[271] * mat_B[498] +
//             mat_A[272] * mat_B[530] +
//             mat_A[273] * mat_B[562] +
//             mat_A[274] * mat_B[594] +
//             mat_A[275] * mat_B[626] +
//             mat_A[276] * mat_B[658] +
//             mat_A[277] * mat_B[690] +
//             mat_A[278] * mat_B[722] +
//             mat_A[279] * mat_B[754] +
//             mat_A[280] * mat_B[786] +
//             mat_A[281] * mat_B[818] +
//             mat_A[282] * mat_B[850] +
//             mat_A[283] * mat_B[882] +
//             mat_A[284] * mat_B[914] +
//             mat_A[285] * mat_B[946] +
//             mat_A[286] * mat_B[978] +
//             mat_A[287] * mat_B[1010];
//  mat_C[275] <= 
//             mat_A[256] * mat_B[19] +
//             mat_A[257] * mat_B[51] +
//             mat_A[258] * mat_B[83] +
//             mat_A[259] * mat_B[115] +
//             mat_A[260] * mat_B[147] +
//             mat_A[261] * mat_B[179] +
//             mat_A[262] * mat_B[211] +
//             mat_A[263] * mat_B[243] +
//             mat_A[264] * mat_B[275] +
//             mat_A[265] * mat_B[307] +
//             mat_A[266] * mat_B[339] +
//             mat_A[267] * mat_B[371] +
//             mat_A[268] * mat_B[403] +
//             mat_A[269] * mat_B[435] +
//             mat_A[270] * mat_B[467] +
//             mat_A[271] * mat_B[499] +
//             mat_A[272] * mat_B[531] +
//             mat_A[273] * mat_B[563] +
//             mat_A[274] * mat_B[595] +
//             mat_A[275] * mat_B[627] +
//             mat_A[276] * mat_B[659] +
//             mat_A[277] * mat_B[691] +
//             mat_A[278] * mat_B[723] +
//             mat_A[279] * mat_B[755] +
//             mat_A[280] * mat_B[787] +
//             mat_A[281] * mat_B[819] +
//             mat_A[282] * mat_B[851] +
//             mat_A[283] * mat_B[883] +
//             mat_A[284] * mat_B[915] +
//             mat_A[285] * mat_B[947] +
//             mat_A[286] * mat_B[979] +
//             mat_A[287] * mat_B[1011];
//  mat_C[276] <= 
//             mat_A[256] * mat_B[20] +
//             mat_A[257] * mat_B[52] +
//             mat_A[258] * mat_B[84] +
//             mat_A[259] * mat_B[116] +
//             mat_A[260] * mat_B[148] +
//             mat_A[261] * mat_B[180] +
//             mat_A[262] * mat_B[212] +
//             mat_A[263] * mat_B[244] +
//             mat_A[264] * mat_B[276] +
//             mat_A[265] * mat_B[308] +
//             mat_A[266] * mat_B[340] +
//             mat_A[267] * mat_B[372] +
//             mat_A[268] * mat_B[404] +
//             mat_A[269] * mat_B[436] +
//             mat_A[270] * mat_B[468] +
//             mat_A[271] * mat_B[500] +
//             mat_A[272] * mat_B[532] +
//             mat_A[273] * mat_B[564] +
//             mat_A[274] * mat_B[596] +
//             mat_A[275] * mat_B[628] +
//             mat_A[276] * mat_B[660] +
//             mat_A[277] * mat_B[692] +
//             mat_A[278] * mat_B[724] +
//             mat_A[279] * mat_B[756] +
//             mat_A[280] * mat_B[788] +
//             mat_A[281] * mat_B[820] +
//             mat_A[282] * mat_B[852] +
//             mat_A[283] * mat_B[884] +
//             mat_A[284] * mat_B[916] +
//             mat_A[285] * mat_B[948] +
//             mat_A[286] * mat_B[980] +
//             mat_A[287] * mat_B[1012];
//  mat_C[277] <= 
//             mat_A[256] * mat_B[21] +
//             mat_A[257] * mat_B[53] +
//             mat_A[258] * mat_B[85] +
//             mat_A[259] * mat_B[117] +
//             mat_A[260] * mat_B[149] +
//             mat_A[261] * mat_B[181] +
//             mat_A[262] * mat_B[213] +
//             mat_A[263] * mat_B[245] +
//             mat_A[264] * mat_B[277] +
//             mat_A[265] * mat_B[309] +
//             mat_A[266] * mat_B[341] +
//             mat_A[267] * mat_B[373] +
//             mat_A[268] * mat_B[405] +
//             mat_A[269] * mat_B[437] +
//             mat_A[270] * mat_B[469] +
//             mat_A[271] * mat_B[501] +
//             mat_A[272] * mat_B[533] +
//             mat_A[273] * mat_B[565] +
//             mat_A[274] * mat_B[597] +
//             mat_A[275] * mat_B[629] +
//             mat_A[276] * mat_B[661] +
//             mat_A[277] * mat_B[693] +
//             mat_A[278] * mat_B[725] +
//             mat_A[279] * mat_B[757] +
//             mat_A[280] * mat_B[789] +
//             mat_A[281] * mat_B[821] +
//             mat_A[282] * mat_B[853] +
//             mat_A[283] * mat_B[885] +
//             mat_A[284] * mat_B[917] +
//             mat_A[285] * mat_B[949] +
//             mat_A[286] * mat_B[981] +
//             mat_A[287] * mat_B[1013];
//  mat_C[278] <= 
//             mat_A[256] * mat_B[22] +
//             mat_A[257] * mat_B[54] +
//             mat_A[258] * mat_B[86] +
//             mat_A[259] * mat_B[118] +
//             mat_A[260] * mat_B[150] +
//             mat_A[261] * mat_B[182] +
//             mat_A[262] * mat_B[214] +
//             mat_A[263] * mat_B[246] +
//             mat_A[264] * mat_B[278] +
//             mat_A[265] * mat_B[310] +
//             mat_A[266] * mat_B[342] +
//             mat_A[267] * mat_B[374] +
//             mat_A[268] * mat_B[406] +
//             mat_A[269] * mat_B[438] +
//             mat_A[270] * mat_B[470] +
//             mat_A[271] * mat_B[502] +
//             mat_A[272] * mat_B[534] +
//             mat_A[273] * mat_B[566] +
//             mat_A[274] * mat_B[598] +
//             mat_A[275] * mat_B[630] +
//             mat_A[276] * mat_B[662] +
//             mat_A[277] * mat_B[694] +
//             mat_A[278] * mat_B[726] +
//             mat_A[279] * mat_B[758] +
//             mat_A[280] * mat_B[790] +
//             mat_A[281] * mat_B[822] +
//             mat_A[282] * mat_B[854] +
//             mat_A[283] * mat_B[886] +
//             mat_A[284] * mat_B[918] +
//             mat_A[285] * mat_B[950] +
//             mat_A[286] * mat_B[982] +
//             mat_A[287] * mat_B[1014];
//  mat_C[279] <= 
//             mat_A[256] * mat_B[23] +
//             mat_A[257] * mat_B[55] +
//             mat_A[258] * mat_B[87] +
//             mat_A[259] * mat_B[119] +
//             mat_A[260] * mat_B[151] +
//             mat_A[261] * mat_B[183] +
//             mat_A[262] * mat_B[215] +
//             mat_A[263] * mat_B[247] +
//             mat_A[264] * mat_B[279] +
//             mat_A[265] * mat_B[311] +
//             mat_A[266] * mat_B[343] +
//             mat_A[267] * mat_B[375] +
//             mat_A[268] * mat_B[407] +
//             mat_A[269] * mat_B[439] +
//             mat_A[270] * mat_B[471] +
//             mat_A[271] * mat_B[503] +
//             mat_A[272] * mat_B[535] +
//             mat_A[273] * mat_B[567] +
//             mat_A[274] * mat_B[599] +
//             mat_A[275] * mat_B[631] +
//             mat_A[276] * mat_B[663] +
//             mat_A[277] * mat_B[695] +
//             mat_A[278] * mat_B[727] +
//             mat_A[279] * mat_B[759] +
//             mat_A[280] * mat_B[791] +
//             mat_A[281] * mat_B[823] +
//             mat_A[282] * mat_B[855] +
//             mat_A[283] * mat_B[887] +
//             mat_A[284] * mat_B[919] +
//             mat_A[285] * mat_B[951] +
//             mat_A[286] * mat_B[983] +
//             mat_A[287] * mat_B[1015];
//  mat_C[280] <= 
//             mat_A[256] * mat_B[24] +
//             mat_A[257] * mat_B[56] +
//             mat_A[258] * mat_B[88] +
//             mat_A[259] * mat_B[120] +
//             mat_A[260] * mat_B[152] +
//             mat_A[261] * mat_B[184] +
//             mat_A[262] * mat_B[216] +
//             mat_A[263] * mat_B[248] +
//             mat_A[264] * mat_B[280] +
//             mat_A[265] * mat_B[312] +
//             mat_A[266] * mat_B[344] +
//             mat_A[267] * mat_B[376] +
//             mat_A[268] * mat_B[408] +
//             mat_A[269] * mat_B[440] +
//             mat_A[270] * mat_B[472] +
//             mat_A[271] * mat_B[504] +
//             mat_A[272] * mat_B[536] +
//             mat_A[273] * mat_B[568] +
//             mat_A[274] * mat_B[600] +
//             mat_A[275] * mat_B[632] +
//             mat_A[276] * mat_B[664] +
//             mat_A[277] * mat_B[696] +
//             mat_A[278] * mat_B[728] +
//             mat_A[279] * mat_B[760] +
//             mat_A[280] * mat_B[792] +
//             mat_A[281] * mat_B[824] +
//             mat_A[282] * mat_B[856] +
//             mat_A[283] * mat_B[888] +
//             mat_A[284] * mat_B[920] +
//             mat_A[285] * mat_B[952] +
//             mat_A[286] * mat_B[984] +
//             mat_A[287] * mat_B[1016];
//  mat_C[281] <= 
//             mat_A[256] * mat_B[25] +
//             mat_A[257] * mat_B[57] +
//             mat_A[258] * mat_B[89] +
//             mat_A[259] * mat_B[121] +
//             mat_A[260] * mat_B[153] +
//             mat_A[261] * mat_B[185] +
//             mat_A[262] * mat_B[217] +
//             mat_A[263] * mat_B[249] +
//             mat_A[264] * mat_B[281] +
//             mat_A[265] * mat_B[313] +
//             mat_A[266] * mat_B[345] +
//             mat_A[267] * mat_B[377] +
//             mat_A[268] * mat_B[409] +
//             mat_A[269] * mat_B[441] +
//             mat_A[270] * mat_B[473] +
//             mat_A[271] * mat_B[505] +
//             mat_A[272] * mat_B[537] +
//             mat_A[273] * mat_B[569] +
//             mat_A[274] * mat_B[601] +
//             mat_A[275] * mat_B[633] +
//             mat_A[276] * mat_B[665] +
//             mat_A[277] * mat_B[697] +
//             mat_A[278] * mat_B[729] +
//             mat_A[279] * mat_B[761] +
//             mat_A[280] * mat_B[793] +
//             mat_A[281] * mat_B[825] +
//             mat_A[282] * mat_B[857] +
//             mat_A[283] * mat_B[889] +
//             mat_A[284] * mat_B[921] +
//             mat_A[285] * mat_B[953] +
//             mat_A[286] * mat_B[985] +
//             mat_A[287] * mat_B[1017];
//  mat_C[282] <= 
//             mat_A[256] * mat_B[26] +
//             mat_A[257] * mat_B[58] +
//             mat_A[258] * mat_B[90] +
//             mat_A[259] * mat_B[122] +
//             mat_A[260] * mat_B[154] +
//             mat_A[261] * mat_B[186] +
//             mat_A[262] * mat_B[218] +
//             mat_A[263] * mat_B[250] +
//             mat_A[264] * mat_B[282] +
//             mat_A[265] * mat_B[314] +
//             mat_A[266] * mat_B[346] +
//             mat_A[267] * mat_B[378] +
//             mat_A[268] * mat_B[410] +
//             mat_A[269] * mat_B[442] +
//             mat_A[270] * mat_B[474] +
//             mat_A[271] * mat_B[506] +
//             mat_A[272] * mat_B[538] +
//             mat_A[273] * mat_B[570] +
//             mat_A[274] * mat_B[602] +
//             mat_A[275] * mat_B[634] +
//             mat_A[276] * mat_B[666] +
//             mat_A[277] * mat_B[698] +
//             mat_A[278] * mat_B[730] +
//             mat_A[279] * mat_B[762] +
//             mat_A[280] * mat_B[794] +
//             mat_A[281] * mat_B[826] +
//             mat_A[282] * mat_B[858] +
//             mat_A[283] * mat_B[890] +
//             mat_A[284] * mat_B[922] +
//             mat_A[285] * mat_B[954] +
//             mat_A[286] * mat_B[986] +
//             mat_A[287] * mat_B[1018];
//  mat_C[283] <= 
//             mat_A[256] * mat_B[27] +
//             mat_A[257] * mat_B[59] +
//             mat_A[258] * mat_B[91] +
//             mat_A[259] * mat_B[123] +
//             mat_A[260] * mat_B[155] +
//             mat_A[261] * mat_B[187] +
//             mat_A[262] * mat_B[219] +
//             mat_A[263] * mat_B[251] +
//             mat_A[264] * mat_B[283] +
//             mat_A[265] * mat_B[315] +
//             mat_A[266] * mat_B[347] +
//             mat_A[267] * mat_B[379] +
//             mat_A[268] * mat_B[411] +
//             mat_A[269] * mat_B[443] +
//             mat_A[270] * mat_B[475] +
//             mat_A[271] * mat_B[507] +
//             mat_A[272] * mat_B[539] +
//             mat_A[273] * mat_B[571] +
//             mat_A[274] * mat_B[603] +
//             mat_A[275] * mat_B[635] +
//             mat_A[276] * mat_B[667] +
//             mat_A[277] * mat_B[699] +
//             mat_A[278] * mat_B[731] +
//             mat_A[279] * mat_B[763] +
//             mat_A[280] * mat_B[795] +
//             mat_A[281] * mat_B[827] +
//             mat_A[282] * mat_B[859] +
//             mat_A[283] * mat_B[891] +
//             mat_A[284] * mat_B[923] +
//             mat_A[285] * mat_B[955] +
//             mat_A[286] * mat_B[987] +
//             mat_A[287] * mat_B[1019];
//  mat_C[284] <= 
//             mat_A[256] * mat_B[28] +
//             mat_A[257] * mat_B[60] +
//             mat_A[258] * mat_B[92] +
//             mat_A[259] * mat_B[124] +
//             mat_A[260] * mat_B[156] +
//             mat_A[261] * mat_B[188] +
//             mat_A[262] * mat_B[220] +
//             mat_A[263] * mat_B[252] +
//             mat_A[264] * mat_B[284] +
//             mat_A[265] * mat_B[316] +
//             mat_A[266] * mat_B[348] +
//             mat_A[267] * mat_B[380] +
//             mat_A[268] * mat_B[412] +
//             mat_A[269] * mat_B[444] +
//             mat_A[270] * mat_B[476] +
//             mat_A[271] * mat_B[508] +
//             mat_A[272] * mat_B[540] +
//             mat_A[273] * mat_B[572] +
//             mat_A[274] * mat_B[604] +
//             mat_A[275] * mat_B[636] +
//             mat_A[276] * mat_B[668] +
//             mat_A[277] * mat_B[700] +
//             mat_A[278] * mat_B[732] +
//             mat_A[279] * mat_B[764] +
//             mat_A[280] * mat_B[796] +
//             mat_A[281] * mat_B[828] +
//             mat_A[282] * mat_B[860] +
//             mat_A[283] * mat_B[892] +
//             mat_A[284] * mat_B[924] +
//             mat_A[285] * mat_B[956] +
//             mat_A[286] * mat_B[988] +
//             mat_A[287] * mat_B[1020];
//  mat_C[285] <= 
//             mat_A[256] * mat_B[29] +
//             mat_A[257] * mat_B[61] +
//             mat_A[258] * mat_B[93] +
//             mat_A[259] * mat_B[125] +
//             mat_A[260] * mat_B[157] +
//             mat_A[261] * mat_B[189] +
//             mat_A[262] * mat_B[221] +
//             mat_A[263] * mat_B[253] +
//             mat_A[264] * mat_B[285] +
//             mat_A[265] * mat_B[317] +
//             mat_A[266] * mat_B[349] +
//             mat_A[267] * mat_B[381] +
//             mat_A[268] * mat_B[413] +
//             mat_A[269] * mat_B[445] +
//             mat_A[270] * mat_B[477] +
//             mat_A[271] * mat_B[509] +
//             mat_A[272] * mat_B[541] +
//             mat_A[273] * mat_B[573] +
//             mat_A[274] * mat_B[605] +
//             mat_A[275] * mat_B[637] +
//             mat_A[276] * mat_B[669] +
//             mat_A[277] * mat_B[701] +
//             mat_A[278] * mat_B[733] +
//             mat_A[279] * mat_B[765] +
//             mat_A[280] * mat_B[797] +
//             mat_A[281] * mat_B[829] +
//             mat_A[282] * mat_B[861] +
//             mat_A[283] * mat_B[893] +
//             mat_A[284] * mat_B[925] +
//             mat_A[285] * mat_B[957] +
//             mat_A[286] * mat_B[989] +
//             mat_A[287] * mat_B[1021];
//  mat_C[286] <= 
//             mat_A[256] * mat_B[30] +
//             mat_A[257] * mat_B[62] +
//             mat_A[258] * mat_B[94] +
//             mat_A[259] * mat_B[126] +
//             mat_A[260] * mat_B[158] +
//             mat_A[261] * mat_B[190] +
//             mat_A[262] * mat_B[222] +
//             mat_A[263] * mat_B[254] +
//             mat_A[264] * mat_B[286] +
//             mat_A[265] * mat_B[318] +
//             mat_A[266] * mat_B[350] +
//             mat_A[267] * mat_B[382] +
//             mat_A[268] * mat_B[414] +
//             mat_A[269] * mat_B[446] +
//             mat_A[270] * mat_B[478] +
//             mat_A[271] * mat_B[510] +
//             mat_A[272] * mat_B[542] +
//             mat_A[273] * mat_B[574] +
//             mat_A[274] * mat_B[606] +
//             mat_A[275] * mat_B[638] +
//             mat_A[276] * mat_B[670] +
//             mat_A[277] * mat_B[702] +
//             mat_A[278] * mat_B[734] +
//             mat_A[279] * mat_B[766] +
//             mat_A[280] * mat_B[798] +
//             mat_A[281] * mat_B[830] +
//             mat_A[282] * mat_B[862] +
//             mat_A[283] * mat_B[894] +
//             mat_A[284] * mat_B[926] +
//             mat_A[285] * mat_B[958] +
//             mat_A[286] * mat_B[990] +
//             mat_A[287] * mat_B[1022];
//  mat_C[287] <= 
//             mat_A[256] * mat_B[31] +
//             mat_A[257] * mat_B[63] +
//             mat_A[258] * mat_B[95] +
//             mat_A[259] * mat_B[127] +
//             mat_A[260] * mat_B[159] +
//             mat_A[261] * mat_B[191] +
//             mat_A[262] * mat_B[223] +
//             mat_A[263] * mat_B[255] +
//             mat_A[264] * mat_B[287] +
//             mat_A[265] * mat_B[319] +
//             mat_A[266] * mat_B[351] +
//             mat_A[267] * mat_B[383] +
//             mat_A[268] * mat_B[415] +
//             mat_A[269] * mat_B[447] +
//             mat_A[270] * mat_B[479] +
//             mat_A[271] * mat_B[511] +
//             mat_A[272] * mat_B[543] +
//             mat_A[273] * mat_B[575] +
//             mat_A[274] * mat_B[607] +
//             mat_A[275] * mat_B[639] +
//             mat_A[276] * mat_B[671] +
//             mat_A[277] * mat_B[703] +
//             mat_A[278] * mat_B[735] +
//             mat_A[279] * mat_B[767] +
//             mat_A[280] * mat_B[799] +
//             mat_A[281] * mat_B[831] +
//             mat_A[282] * mat_B[863] +
//             mat_A[283] * mat_B[895] +
//             mat_A[284] * mat_B[927] +
//             mat_A[285] * mat_B[959] +
//             mat_A[286] * mat_B[991] +
//             mat_A[287] * mat_B[1023];
//  mat_C[288] <= 
//             mat_A[288] * mat_B[0] +
//             mat_A[289] * mat_B[32] +
//             mat_A[290] * mat_B[64] +
//             mat_A[291] * mat_B[96] +
//             mat_A[292] * mat_B[128] +
//             mat_A[293] * mat_B[160] +
//             mat_A[294] * mat_B[192] +
//             mat_A[295] * mat_B[224] +
//             mat_A[296] * mat_B[256] +
//             mat_A[297] * mat_B[288] +
//             mat_A[298] * mat_B[320] +
//             mat_A[299] * mat_B[352] +
//             mat_A[300] * mat_B[384] +
//             mat_A[301] * mat_B[416] +
//             mat_A[302] * mat_B[448] +
//             mat_A[303] * mat_B[480] +
//             mat_A[304] * mat_B[512] +
//             mat_A[305] * mat_B[544] +
//             mat_A[306] * mat_B[576] +
//             mat_A[307] * mat_B[608] +
//             mat_A[308] * mat_B[640] +
//             mat_A[309] * mat_B[672] +
//             mat_A[310] * mat_B[704] +
//             mat_A[311] * mat_B[736] +
//             mat_A[312] * mat_B[768] +
//             mat_A[313] * mat_B[800] +
//             mat_A[314] * mat_B[832] +
//             mat_A[315] * mat_B[864] +
//             mat_A[316] * mat_B[896] +
//             mat_A[317] * mat_B[928] +
//             mat_A[318] * mat_B[960] +
//             mat_A[319] * mat_B[992];
//  mat_C[289] <= 
//             mat_A[288] * mat_B[1] +
//             mat_A[289] * mat_B[33] +
//             mat_A[290] * mat_B[65] +
//             mat_A[291] * mat_B[97] +
//             mat_A[292] * mat_B[129] +
//             mat_A[293] * mat_B[161] +
//             mat_A[294] * mat_B[193] +
//             mat_A[295] * mat_B[225] +
//             mat_A[296] * mat_B[257] +
//             mat_A[297] * mat_B[289] +
//             mat_A[298] * mat_B[321] +
//             mat_A[299] * mat_B[353] +
//             mat_A[300] * mat_B[385] +
//             mat_A[301] * mat_B[417] +
//             mat_A[302] * mat_B[449] +
//             mat_A[303] * mat_B[481] +
//             mat_A[304] * mat_B[513] +
//             mat_A[305] * mat_B[545] +
//             mat_A[306] * mat_B[577] +
//             mat_A[307] * mat_B[609] +
//             mat_A[308] * mat_B[641] +
//             mat_A[309] * mat_B[673] +
//             mat_A[310] * mat_B[705] +
//             mat_A[311] * mat_B[737] +
//             mat_A[312] * mat_B[769] +
//             mat_A[313] * mat_B[801] +
//             mat_A[314] * mat_B[833] +
//             mat_A[315] * mat_B[865] +
//             mat_A[316] * mat_B[897] +
//             mat_A[317] * mat_B[929] +
//             mat_A[318] * mat_B[961] +
//             mat_A[319] * mat_B[993];
//  mat_C[290] <= 
//             mat_A[288] * mat_B[2] +
//             mat_A[289] * mat_B[34] +
//             mat_A[290] * mat_B[66] +
//             mat_A[291] * mat_B[98] +
//             mat_A[292] * mat_B[130] +
//             mat_A[293] * mat_B[162] +
//             mat_A[294] * mat_B[194] +
//             mat_A[295] * mat_B[226] +
//             mat_A[296] * mat_B[258] +
//             mat_A[297] * mat_B[290] +
//             mat_A[298] * mat_B[322] +
//             mat_A[299] * mat_B[354] +
//             mat_A[300] * mat_B[386] +
//             mat_A[301] * mat_B[418] +
//             mat_A[302] * mat_B[450] +
//             mat_A[303] * mat_B[482] +
//             mat_A[304] * mat_B[514] +
//             mat_A[305] * mat_B[546] +
//             mat_A[306] * mat_B[578] +
//             mat_A[307] * mat_B[610] +
//             mat_A[308] * mat_B[642] +
//             mat_A[309] * mat_B[674] +
//             mat_A[310] * mat_B[706] +
//             mat_A[311] * mat_B[738] +
//             mat_A[312] * mat_B[770] +
//             mat_A[313] * mat_B[802] +
//             mat_A[314] * mat_B[834] +
//             mat_A[315] * mat_B[866] +
//             mat_A[316] * mat_B[898] +
//             mat_A[317] * mat_B[930] +
//             mat_A[318] * mat_B[962] +
//             mat_A[319] * mat_B[994];
//  mat_C[291] <= 
//             mat_A[288] * mat_B[3] +
//             mat_A[289] * mat_B[35] +
//             mat_A[290] * mat_B[67] +
//             mat_A[291] * mat_B[99] +
//             mat_A[292] * mat_B[131] +
//             mat_A[293] * mat_B[163] +
//             mat_A[294] * mat_B[195] +
//             mat_A[295] * mat_B[227] +
//             mat_A[296] * mat_B[259] +
//             mat_A[297] * mat_B[291] +
//             mat_A[298] * mat_B[323] +
//             mat_A[299] * mat_B[355] +
//             mat_A[300] * mat_B[387] +
//             mat_A[301] * mat_B[419] +
//             mat_A[302] * mat_B[451] +
//             mat_A[303] * mat_B[483] +
//             mat_A[304] * mat_B[515] +
//             mat_A[305] * mat_B[547] +
//             mat_A[306] * mat_B[579] +
//             mat_A[307] * mat_B[611] +
//             mat_A[308] * mat_B[643] +
//             mat_A[309] * mat_B[675] +
//             mat_A[310] * mat_B[707] +
//             mat_A[311] * mat_B[739] +
//             mat_A[312] * mat_B[771] +
//             mat_A[313] * mat_B[803] +
//             mat_A[314] * mat_B[835] +
//             mat_A[315] * mat_B[867] +
//             mat_A[316] * mat_B[899] +
//             mat_A[317] * mat_B[931] +
//             mat_A[318] * mat_B[963] +
//             mat_A[319] * mat_B[995];
//  mat_C[292] <= 
//             mat_A[288] * mat_B[4] +
//             mat_A[289] * mat_B[36] +
//             mat_A[290] * mat_B[68] +
//             mat_A[291] * mat_B[100] +
//             mat_A[292] * mat_B[132] +
//             mat_A[293] * mat_B[164] +
//             mat_A[294] * mat_B[196] +
//             mat_A[295] * mat_B[228] +
//             mat_A[296] * mat_B[260] +
//             mat_A[297] * mat_B[292] +
//             mat_A[298] * mat_B[324] +
//             mat_A[299] * mat_B[356] +
//             mat_A[300] * mat_B[388] +
//             mat_A[301] * mat_B[420] +
//             mat_A[302] * mat_B[452] +
//             mat_A[303] * mat_B[484] +
//             mat_A[304] * mat_B[516] +
//             mat_A[305] * mat_B[548] +
//             mat_A[306] * mat_B[580] +
//             mat_A[307] * mat_B[612] +
//             mat_A[308] * mat_B[644] +
//             mat_A[309] * mat_B[676] +
//             mat_A[310] * mat_B[708] +
//             mat_A[311] * mat_B[740] +
//             mat_A[312] * mat_B[772] +
//             mat_A[313] * mat_B[804] +
//             mat_A[314] * mat_B[836] +
//             mat_A[315] * mat_B[868] +
//             mat_A[316] * mat_B[900] +
//             mat_A[317] * mat_B[932] +
//             mat_A[318] * mat_B[964] +
//             mat_A[319] * mat_B[996];
//  mat_C[293] <= 
//             mat_A[288] * mat_B[5] +
//             mat_A[289] * mat_B[37] +
//             mat_A[290] * mat_B[69] +
//             mat_A[291] * mat_B[101] +
//             mat_A[292] * mat_B[133] +
//             mat_A[293] * mat_B[165] +
//             mat_A[294] * mat_B[197] +
//             mat_A[295] * mat_B[229] +
//             mat_A[296] * mat_B[261] +
//             mat_A[297] * mat_B[293] +
//             mat_A[298] * mat_B[325] +
//             mat_A[299] * mat_B[357] +
//             mat_A[300] * mat_B[389] +
//             mat_A[301] * mat_B[421] +
//             mat_A[302] * mat_B[453] +
//             mat_A[303] * mat_B[485] +
//             mat_A[304] * mat_B[517] +
//             mat_A[305] * mat_B[549] +
//             mat_A[306] * mat_B[581] +
//             mat_A[307] * mat_B[613] +
//             mat_A[308] * mat_B[645] +
//             mat_A[309] * mat_B[677] +
//             mat_A[310] * mat_B[709] +
//             mat_A[311] * mat_B[741] +
//             mat_A[312] * mat_B[773] +
//             mat_A[313] * mat_B[805] +
//             mat_A[314] * mat_B[837] +
//             mat_A[315] * mat_B[869] +
//             mat_A[316] * mat_B[901] +
//             mat_A[317] * mat_B[933] +
//             mat_A[318] * mat_B[965] +
//             mat_A[319] * mat_B[997];
//  mat_C[294] <= 
//             mat_A[288] * mat_B[6] +
//             mat_A[289] * mat_B[38] +
//             mat_A[290] * mat_B[70] +
//             mat_A[291] * mat_B[102] +
//             mat_A[292] * mat_B[134] +
//             mat_A[293] * mat_B[166] +
//             mat_A[294] * mat_B[198] +
//             mat_A[295] * mat_B[230] +
//             mat_A[296] * mat_B[262] +
//             mat_A[297] * mat_B[294] +
//             mat_A[298] * mat_B[326] +
//             mat_A[299] * mat_B[358] +
//             mat_A[300] * mat_B[390] +
//             mat_A[301] * mat_B[422] +
//             mat_A[302] * mat_B[454] +
//             mat_A[303] * mat_B[486] +
//             mat_A[304] * mat_B[518] +
//             mat_A[305] * mat_B[550] +
//             mat_A[306] * mat_B[582] +
//             mat_A[307] * mat_B[614] +
//             mat_A[308] * mat_B[646] +
//             mat_A[309] * mat_B[678] +
//             mat_A[310] * mat_B[710] +
//             mat_A[311] * mat_B[742] +
//             mat_A[312] * mat_B[774] +
//             mat_A[313] * mat_B[806] +
//             mat_A[314] * mat_B[838] +
//             mat_A[315] * mat_B[870] +
//             mat_A[316] * mat_B[902] +
//             mat_A[317] * mat_B[934] +
//             mat_A[318] * mat_B[966] +
//             mat_A[319] * mat_B[998];
//  mat_C[295] <= 
//             mat_A[288] * mat_B[7] +
//             mat_A[289] * mat_B[39] +
//             mat_A[290] * mat_B[71] +
//             mat_A[291] * mat_B[103] +
//             mat_A[292] * mat_B[135] +
//             mat_A[293] * mat_B[167] +
//             mat_A[294] * mat_B[199] +
//             mat_A[295] * mat_B[231] +
//             mat_A[296] * mat_B[263] +
//             mat_A[297] * mat_B[295] +
//             mat_A[298] * mat_B[327] +
//             mat_A[299] * mat_B[359] +
//             mat_A[300] * mat_B[391] +
//             mat_A[301] * mat_B[423] +
//             mat_A[302] * mat_B[455] +
//             mat_A[303] * mat_B[487] +
//             mat_A[304] * mat_B[519] +
//             mat_A[305] * mat_B[551] +
//             mat_A[306] * mat_B[583] +
//             mat_A[307] * mat_B[615] +
//             mat_A[308] * mat_B[647] +
//             mat_A[309] * mat_B[679] +
//             mat_A[310] * mat_B[711] +
//             mat_A[311] * mat_B[743] +
//             mat_A[312] * mat_B[775] +
//             mat_A[313] * mat_B[807] +
//             mat_A[314] * mat_B[839] +
//             mat_A[315] * mat_B[871] +
//             mat_A[316] * mat_B[903] +
//             mat_A[317] * mat_B[935] +
//             mat_A[318] * mat_B[967] +
//             mat_A[319] * mat_B[999];
//  mat_C[296] <= 
//             mat_A[288] * mat_B[8] +
//             mat_A[289] * mat_B[40] +
//             mat_A[290] * mat_B[72] +
//             mat_A[291] * mat_B[104] +
//             mat_A[292] * mat_B[136] +
//             mat_A[293] * mat_B[168] +
//             mat_A[294] * mat_B[200] +
//             mat_A[295] * mat_B[232] +
//             mat_A[296] * mat_B[264] +
//             mat_A[297] * mat_B[296] +
//             mat_A[298] * mat_B[328] +
//             mat_A[299] * mat_B[360] +
//             mat_A[300] * mat_B[392] +
//             mat_A[301] * mat_B[424] +
//             mat_A[302] * mat_B[456] +
//             mat_A[303] * mat_B[488] +
//             mat_A[304] * mat_B[520] +
//             mat_A[305] * mat_B[552] +
//             mat_A[306] * mat_B[584] +
//             mat_A[307] * mat_B[616] +
//             mat_A[308] * mat_B[648] +
//             mat_A[309] * mat_B[680] +
//             mat_A[310] * mat_B[712] +
//             mat_A[311] * mat_B[744] +
//             mat_A[312] * mat_B[776] +
//             mat_A[313] * mat_B[808] +
//             mat_A[314] * mat_B[840] +
//             mat_A[315] * mat_B[872] +
//             mat_A[316] * mat_B[904] +
//             mat_A[317] * mat_B[936] +
//             mat_A[318] * mat_B[968] +
//             mat_A[319] * mat_B[1000];
//  mat_C[297] <= 
//             mat_A[288] * mat_B[9] +
//             mat_A[289] * mat_B[41] +
//             mat_A[290] * mat_B[73] +
//             mat_A[291] * mat_B[105] +
//             mat_A[292] * mat_B[137] +
//             mat_A[293] * mat_B[169] +
//             mat_A[294] * mat_B[201] +
//             mat_A[295] * mat_B[233] +
//             mat_A[296] * mat_B[265] +
//             mat_A[297] * mat_B[297] +
//             mat_A[298] * mat_B[329] +
//             mat_A[299] * mat_B[361] +
//             mat_A[300] * mat_B[393] +
//             mat_A[301] * mat_B[425] +
//             mat_A[302] * mat_B[457] +
//             mat_A[303] * mat_B[489] +
//             mat_A[304] * mat_B[521] +
//             mat_A[305] * mat_B[553] +
//             mat_A[306] * mat_B[585] +
//             mat_A[307] * mat_B[617] +
//             mat_A[308] * mat_B[649] +
//             mat_A[309] * mat_B[681] +
//             mat_A[310] * mat_B[713] +
//             mat_A[311] * mat_B[745] +
//             mat_A[312] * mat_B[777] +
//             mat_A[313] * mat_B[809] +
//             mat_A[314] * mat_B[841] +
//             mat_A[315] * mat_B[873] +
//             mat_A[316] * mat_B[905] +
//             mat_A[317] * mat_B[937] +
//             mat_A[318] * mat_B[969] +
//             mat_A[319] * mat_B[1001];
//  mat_C[298] <= 
//             mat_A[288] * mat_B[10] +
//             mat_A[289] * mat_B[42] +
//             mat_A[290] * mat_B[74] +
//             mat_A[291] * mat_B[106] +
//             mat_A[292] * mat_B[138] +
//             mat_A[293] * mat_B[170] +
//             mat_A[294] * mat_B[202] +
//             mat_A[295] * mat_B[234] +
//             mat_A[296] * mat_B[266] +
//             mat_A[297] * mat_B[298] +
//             mat_A[298] * mat_B[330] +
//             mat_A[299] * mat_B[362] +
//             mat_A[300] * mat_B[394] +
//             mat_A[301] * mat_B[426] +
//             mat_A[302] * mat_B[458] +
//             mat_A[303] * mat_B[490] +
//             mat_A[304] * mat_B[522] +
//             mat_A[305] * mat_B[554] +
//             mat_A[306] * mat_B[586] +
//             mat_A[307] * mat_B[618] +
//             mat_A[308] * mat_B[650] +
//             mat_A[309] * mat_B[682] +
//             mat_A[310] * mat_B[714] +
//             mat_A[311] * mat_B[746] +
//             mat_A[312] * mat_B[778] +
//             mat_A[313] * mat_B[810] +
//             mat_A[314] * mat_B[842] +
//             mat_A[315] * mat_B[874] +
//             mat_A[316] * mat_B[906] +
//             mat_A[317] * mat_B[938] +
//             mat_A[318] * mat_B[970] +
//             mat_A[319] * mat_B[1002];
//  mat_C[299] <= 
//             mat_A[288] * mat_B[11] +
//             mat_A[289] * mat_B[43] +
//             mat_A[290] * mat_B[75] +
//             mat_A[291] * mat_B[107] +
//             mat_A[292] * mat_B[139] +
//             mat_A[293] * mat_B[171] +
//             mat_A[294] * mat_B[203] +
//             mat_A[295] * mat_B[235] +
//             mat_A[296] * mat_B[267] +
//             mat_A[297] * mat_B[299] +
//             mat_A[298] * mat_B[331] +
//             mat_A[299] * mat_B[363] +
//             mat_A[300] * mat_B[395] +
//             mat_A[301] * mat_B[427] +
//             mat_A[302] * mat_B[459] +
//             mat_A[303] * mat_B[491] +
//             mat_A[304] * mat_B[523] +
//             mat_A[305] * mat_B[555] +
//             mat_A[306] * mat_B[587] +
//             mat_A[307] * mat_B[619] +
//             mat_A[308] * mat_B[651] +
//             mat_A[309] * mat_B[683] +
//             mat_A[310] * mat_B[715] +
//             mat_A[311] * mat_B[747] +
//             mat_A[312] * mat_B[779] +
//             mat_A[313] * mat_B[811] +
//             mat_A[314] * mat_B[843] +
//             mat_A[315] * mat_B[875] +
//             mat_A[316] * mat_B[907] +
//             mat_A[317] * mat_B[939] +
//             mat_A[318] * mat_B[971] +
//             mat_A[319] * mat_B[1003];
//  mat_C[300] <= 
//             mat_A[288] * mat_B[12] +
//             mat_A[289] * mat_B[44] +
//             mat_A[290] * mat_B[76] +
//             mat_A[291] * mat_B[108] +
//             mat_A[292] * mat_B[140] +
//             mat_A[293] * mat_B[172] +
//             mat_A[294] * mat_B[204] +
//             mat_A[295] * mat_B[236] +
//             mat_A[296] * mat_B[268] +
//             mat_A[297] * mat_B[300] +
//             mat_A[298] * mat_B[332] +
//             mat_A[299] * mat_B[364] +
//             mat_A[300] * mat_B[396] +
//             mat_A[301] * mat_B[428] +
//             mat_A[302] * mat_B[460] +
//             mat_A[303] * mat_B[492] +
//             mat_A[304] * mat_B[524] +
//             mat_A[305] * mat_B[556] +
//             mat_A[306] * mat_B[588] +
//             mat_A[307] * mat_B[620] +
//             mat_A[308] * mat_B[652] +
//             mat_A[309] * mat_B[684] +
//             mat_A[310] * mat_B[716] +
//             mat_A[311] * mat_B[748] +
//             mat_A[312] * mat_B[780] +
//             mat_A[313] * mat_B[812] +
//             mat_A[314] * mat_B[844] +
//             mat_A[315] * mat_B[876] +
//             mat_A[316] * mat_B[908] +
//             mat_A[317] * mat_B[940] +
//             mat_A[318] * mat_B[972] +
//             mat_A[319] * mat_B[1004];
//  mat_C[301] <= 
//             mat_A[288] * mat_B[13] +
//             mat_A[289] * mat_B[45] +
//             mat_A[290] * mat_B[77] +
//             mat_A[291] * mat_B[109] +
//             mat_A[292] * mat_B[141] +
//             mat_A[293] * mat_B[173] +
//             mat_A[294] * mat_B[205] +
//             mat_A[295] * mat_B[237] +
//             mat_A[296] * mat_B[269] +
//             mat_A[297] * mat_B[301] +
//             mat_A[298] * mat_B[333] +
//             mat_A[299] * mat_B[365] +
//             mat_A[300] * mat_B[397] +
//             mat_A[301] * mat_B[429] +
//             mat_A[302] * mat_B[461] +
//             mat_A[303] * mat_B[493] +
//             mat_A[304] * mat_B[525] +
//             mat_A[305] * mat_B[557] +
//             mat_A[306] * mat_B[589] +
//             mat_A[307] * mat_B[621] +
//             mat_A[308] * mat_B[653] +
//             mat_A[309] * mat_B[685] +
//             mat_A[310] * mat_B[717] +
//             mat_A[311] * mat_B[749] +
//             mat_A[312] * mat_B[781] +
//             mat_A[313] * mat_B[813] +
//             mat_A[314] * mat_B[845] +
//             mat_A[315] * mat_B[877] +
//             mat_A[316] * mat_B[909] +
//             mat_A[317] * mat_B[941] +
//             mat_A[318] * mat_B[973] +
//             mat_A[319] * mat_B[1005];
//  mat_C[302] <= 
//             mat_A[288] * mat_B[14] +
//             mat_A[289] * mat_B[46] +
//             mat_A[290] * mat_B[78] +
//             mat_A[291] * mat_B[110] +
//             mat_A[292] * mat_B[142] +
//             mat_A[293] * mat_B[174] +
//             mat_A[294] * mat_B[206] +
//             mat_A[295] * mat_B[238] +
//             mat_A[296] * mat_B[270] +
//             mat_A[297] * mat_B[302] +
//             mat_A[298] * mat_B[334] +
//             mat_A[299] * mat_B[366] +
//             mat_A[300] * mat_B[398] +
//             mat_A[301] * mat_B[430] +
//             mat_A[302] * mat_B[462] +
//             mat_A[303] * mat_B[494] +
//             mat_A[304] * mat_B[526] +
//             mat_A[305] * mat_B[558] +
//             mat_A[306] * mat_B[590] +
//             mat_A[307] * mat_B[622] +
//             mat_A[308] * mat_B[654] +
//             mat_A[309] * mat_B[686] +
//             mat_A[310] * mat_B[718] +
//             mat_A[311] * mat_B[750] +
//             mat_A[312] * mat_B[782] +
//             mat_A[313] * mat_B[814] +
//             mat_A[314] * mat_B[846] +
//             mat_A[315] * mat_B[878] +
//             mat_A[316] * mat_B[910] +
//             mat_A[317] * mat_B[942] +
//             mat_A[318] * mat_B[974] +
//             mat_A[319] * mat_B[1006];
//  mat_C[303] <= 
//             mat_A[288] * mat_B[15] +
//             mat_A[289] * mat_B[47] +
//             mat_A[290] * mat_B[79] +
//             mat_A[291] * mat_B[111] +
//             mat_A[292] * mat_B[143] +
//             mat_A[293] * mat_B[175] +
//             mat_A[294] * mat_B[207] +
//             mat_A[295] * mat_B[239] +
//             mat_A[296] * mat_B[271] +
//             mat_A[297] * mat_B[303] +
//             mat_A[298] * mat_B[335] +
//             mat_A[299] * mat_B[367] +
//             mat_A[300] * mat_B[399] +
//             mat_A[301] * mat_B[431] +
//             mat_A[302] * mat_B[463] +
//             mat_A[303] * mat_B[495] +
//             mat_A[304] * mat_B[527] +
//             mat_A[305] * mat_B[559] +
//             mat_A[306] * mat_B[591] +
//             mat_A[307] * mat_B[623] +
//             mat_A[308] * mat_B[655] +
//             mat_A[309] * mat_B[687] +
//             mat_A[310] * mat_B[719] +
//             mat_A[311] * mat_B[751] +
//             mat_A[312] * mat_B[783] +
//             mat_A[313] * mat_B[815] +
//             mat_A[314] * mat_B[847] +
//             mat_A[315] * mat_B[879] +
//             mat_A[316] * mat_B[911] +
//             mat_A[317] * mat_B[943] +
//             mat_A[318] * mat_B[975] +
//             mat_A[319] * mat_B[1007];
//  mat_C[304] <= 
//             mat_A[288] * mat_B[16] +
//             mat_A[289] * mat_B[48] +
//             mat_A[290] * mat_B[80] +
//             mat_A[291] * mat_B[112] +
//             mat_A[292] * mat_B[144] +
//             mat_A[293] * mat_B[176] +
//             mat_A[294] * mat_B[208] +
//             mat_A[295] * mat_B[240] +
//             mat_A[296] * mat_B[272] +
//             mat_A[297] * mat_B[304] +
//             mat_A[298] * mat_B[336] +
//             mat_A[299] * mat_B[368] +
//             mat_A[300] * mat_B[400] +
//             mat_A[301] * mat_B[432] +
//             mat_A[302] * mat_B[464] +
//             mat_A[303] * mat_B[496] +
//             mat_A[304] * mat_B[528] +
//             mat_A[305] * mat_B[560] +
//             mat_A[306] * mat_B[592] +
//             mat_A[307] * mat_B[624] +
//             mat_A[308] * mat_B[656] +
//             mat_A[309] * mat_B[688] +
//             mat_A[310] * mat_B[720] +
//             mat_A[311] * mat_B[752] +
//             mat_A[312] * mat_B[784] +
//             mat_A[313] * mat_B[816] +
//             mat_A[314] * mat_B[848] +
//             mat_A[315] * mat_B[880] +
//             mat_A[316] * mat_B[912] +
//             mat_A[317] * mat_B[944] +
//             mat_A[318] * mat_B[976] +
//             mat_A[319] * mat_B[1008];
//  mat_C[305] <= 
//             mat_A[288] * mat_B[17] +
//             mat_A[289] * mat_B[49] +
//             mat_A[290] * mat_B[81] +
//             mat_A[291] * mat_B[113] +
//             mat_A[292] * mat_B[145] +
//             mat_A[293] * mat_B[177] +
//             mat_A[294] * mat_B[209] +
//             mat_A[295] * mat_B[241] +
//             mat_A[296] * mat_B[273] +
//             mat_A[297] * mat_B[305] +
//             mat_A[298] * mat_B[337] +
//             mat_A[299] * mat_B[369] +
//             mat_A[300] * mat_B[401] +
//             mat_A[301] * mat_B[433] +
//             mat_A[302] * mat_B[465] +
//             mat_A[303] * mat_B[497] +
//             mat_A[304] * mat_B[529] +
//             mat_A[305] * mat_B[561] +
//             mat_A[306] * mat_B[593] +
//             mat_A[307] * mat_B[625] +
//             mat_A[308] * mat_B[657] +
//             mat_A[309] * mat_B[689] +
//             mat_A[310] * mat_B[721] +
//             mat_A[311] * mat_B[753] +
//             mat_A[312] * mat_B[785] +
//             mat_A[313] * mat_B[817] +
//             mat_A[314] * mat_B[849] +
//             mat_A[315] * mat_B[881] +
//             mat_A[316] * mat_B[913] +
//             mat_A[317] * mat_B[945] +
//             mat_A[318] * mat_B[977] +
//             mat_A[319] * mat_B[1009];
//  mat_C[306] <= 
//             mat_A[288] * mat_B[18] +
//             mat_A[289] * mat_B[50] +
//             mat_A[290] * mat_B[82] +
//             mat_A[291] * mat_B[114] +
//             mat_A[292] * mat_B[146] +
//             mat_A[293] * mat_B[178] +
//             mat_A[294] * mat_B[210] +
//             mat_A[295] * mat_B[242] +
//             mat_A[296] * mat_B[274] +
//             mat_A[297] * mat_B[306] +
//             mat_A[298] * mat_B[338] +
//             mat_A[299] * mat_B[370] +
//             mat_A[300] * mat_B[402] +
//             mat_A[301] * mat_B[434] +
//             mat_A[302] * mat_B[466] +
//             mat_A[303] * mat_B[498] +
//             mat_A[304] * mat_B[530] +
//             mat_A[305] * mat_B[562] +
//             mat_A[306] * mat_B[594] +
//             mat_A[307] * mat_B[626] +
//             mat_A[308] * mat_B[658] +
//             mat_A[309] * mat_B[690] +
//             mat_A[310] * mat_B[722] +
//             mat_A[311] * mat_B[754] +
//             mat_A[312] * mat_B[786] +
//             mat_A[313] * mat_B[818] +
//             mat_A[314] * mat_B[850] +
//             mat_A[315] * mat_B[882] +
//             mat_A[316] * mat_B[914] +
//             mat_A[317] * mat_B[946] +
//             mat_A[318] * mat_B[978] +
//             mat_A[319] * mat_B[1010];
//  mat_C[307] <= 
//             mat_A[288] * mat_B[19] +
//             mat_A[289] * mat_B[51] +
//             mat_A[290] * mat_B[83] +
//             mat_A[291] * mat_B[115] +
//             mat_A[292] * mat_B[147] +
//             mat_A[293] * mat_B[179] +
//             mat_A[294] * mat_B[211] +
//             mat_A[295] * mat_B[243] +
//             mat_A[296] * mat_B[275] +
//             mat_A[297] * mat_B[307] +
//             mat_A[298] * mat_B[339] +
//             mat_A[299] * mat_B[371] +
//             mat_A[300] * mat_B[403] +
//             mat_A[301] * mat_B[435] +
//             mat_A[302] * mat_B[467] +
//             mat_A[303] * mat_B[499] +
//             mat_A[304] * mat_B[531] +
//             mat_A[305] * mat_B[563] +
//             mat_A[306] * mat_B[595] +
//             mat_A[307] * mat_B[627] +
//             mat_A[308] * mat_B[659] +
//             mat_A[309] * mat_B[691] +
//             mat_A[310] * mat_B[723] +
//             mat_A[311] * mat_B[755] +
//             mat_A[312] * mat_B[787] +
//             mat_A[313] * mat_B[819] +
//             mat_A[314] * mat_B[851] +
//             mat_A[315] * mat_B[883] +
//             mat_A[316] * mat_B[915] +
//             mat_A[317] * mat_B[947] +
//             mat_A[318] * mat_B[979] +
//             mat_A[319] * mat_B[1011];
//  mat_C[308] <= 
//             mat_A[288] * mat_B[20] +
//             mat_A[289] * mat_B[52] +
//             mat_A[290] * mat_B[84] +
//             mat_A[291] * mat_B[116] +
//             mat_A[292] * mat_B[148] +
//             mat_A[293] * mat_B[180] +
//             mat_A[294] * mat_B[212] +
//             mat_A[295] * mat_B[244] +
//             mat_A[296] * mat_B[276] +
//             mat_A[297] * mat_B[308] +
//             mat_A[298] * mat_B[340] +
//             mat_A[299] * mat_B[372] +
//             mat_A[300] * mat_B[404] +
//             mat_A[301] * mat_B[436] +
//             mat_A[302] * mat_B[468] +
//             mat_A[303] * mat_B[500] +
//             mat_A[304] * mat_B[532] +
//             mat_A[305] * mat_B[564] +
//             mat_A[306] * mat_B[596] +
//             mat_A[307] * mat_B[628] +
//             mat_A[308] * mat_B[660] +
//             mat_A[309] * mat_B[692] +
//             mat_A[310] * mat_B[724] +
//             mat_A[311] * mat_B[756] +
//             mat_A[312] * mat_B[788] +
//             mat_A[313] * mat_B[820] +
//             mat_A[314] * mat_B[852] +
//             mat_A[315] * mat_B[884] +
//             mat_A[316] * mat_B[916] +
//             mat_A[317] * mat_B[948] +
//             mat_A[318] * mat_B[980] +
//             mat_A[319] * mat_B[1012];
//  mat_C[309] <= 
//             mat_A[288] * mat_B[21] +
//             mat_A[289] * mat_B[53] +
//             mat_A[290] * mat_B[85] +
//             mat_A[291] * mat_B[117] +
//             mat_A[292] * mat_B[149] +
//             mat_A[293] * mat_B[181] +
//             mat_A[294] * mat_B[213] +
//             mat_A[295] * mat_B[245] +
//             mat_A[296] * mat_B[277] +
//             mat_A[297] * mat_B[309] +
//             mat_A[298] * mat_B[341] +
//             mat_A[299] * mat_B[373] +
//             mat_A[300] * mat_B[405] +
//             mat_A[301] * mat_B[437] +
//             mat_A[302] * mat_B[469] +
//             mat_A[303] * mat_B[501] +
//             mat_A[304] * mat_B[533] +
//             mat_A[305] * mat_B[565] +
//             mat_A[306] * mat_B[597] +
//             mat_A[307] * mat_B[629] +
//             mat_A[308] * mat_B[661] +
//             mat_A[309] * mat_B[693] +
//             mat_A[310] * mat_B[725] +
//             mat_A[311] * mat_B[757] +
//             mat_A[312] * mat_B[789] +
//             mat_A[313] * mat_B[821] +
//             mat_A[314] * mat_B[853] +
//             mat_A[315] * mat_B[885] +
//             mat_A[316] * mat_B[917] +
//             mat_A[317] * mat_B[949] +
//             mat_A[318] * mat_B[981] +
//             mat_A[319] * mat_B[1013];
//  mat_C[310] <= 
//             mat_A[288] * mat_B[22] +
//             mat_A[289] * mat_B[54] +
//             mat_A[290] * mat_B[86] +
//             mat_A[291] * mat_B[118] +
//             mat_A[292] * mat_B[150] +
//             mat_A[293] * mat_B[182] +
//             mat_A[294] * mat_B[214] +
//             mat_A[295] * mat_B[246] +
//             mat_A[296] * mat_B[278] +
//             mat_A[297] * mat_B[310] +
//             mat_A[298] * mat_B[342] +
//             mat_A[299] * mat_B[374] +
//             mat_A[300] * mat_B[406] +
//             mat_A[301] * mat_B[438] +
//             mat_A[302] * mat_B[470] +
//             mat_A[303] * mat_B[502] +
//             mat_A[304] * mat_B[534] +
//             mat_A[305] * mat_B[566] +
//             mat_A[306] * mat_B[598] +
//             mat_A[307] * mat_B[630] +
//             mat_A[308] * mat_B[662] +
//             mat_A[309] * mat_B[694] +
//             mat_A[310] * mat_B[726] +
//             mat_A[311] * mat_B[758] +
//             mat_A[312] * mat_B[790] +
//             mat_A[313] * mat_B[822] +
//             mat_A[314] * mat_B[854] +
//             mat_A[315] * mat_B[886] +
//             mat_A[316] * mat_B[918] +
//             mat_A[317] * mat_B[950] +
//             mat_A[318] * mat_B[982] +
//             mat_A[319] * mat_B[1014];
//  mat_C[311] <= 
//             mat_A[288] * mat_B[23] +
//             mat_A[289] * mat_B[55] +
//             mat_A[290] * mat_B[87] +
//             mat_A[291] * mat_B[119] +
//             mat_A[292] * mat_B[151] +
//             mat_A[293] * mat_B[183] +
//             mat_A[294] * mat_B[215] +
//             mat_A[295] * mat_B[247] +
//             mat_A[296] * mat_B[279] +
//             mat_A[297] * mat_B[311] +
//             mat_A[298] * mat_B[343] +
//             mat_A[299] * mat_B[375] +
//             mat_A[300] * mat_B[407] +
//             mat_A[301] * mat_B[439] +
//             mat_A[302] * mat_B[471] +
//             mat_A[303] * mat_B[503] +
//             mat_A[304] * mat_B[535] +
//             mat_A[305] * mat_B[567] +
//             mat_A[306] * mat_B[599] +
//             mat_A[307] * mat_B[631] +
//             mat_A[308] * mat_B[663] +
//             mat_A[309] * mat_B[695] +
//             mat_A[310] * mat_B[727] +
//             mat_A[311] * mat_B[759] +
//             mat_A[312] * mat_B[791] +
//             mat_A[313] * mat_B[823] +
//             mat_A[314] * mat_B[855] +
//             mat_A[315] * mat_B[887] +
//             mat_A[316] * mat_B[919] +
//             mat_A[317] * mat_B[951] +
//             mat_A[318] * mat_B[983] +
//             mat_A[319] * mat_B[1015];
//  mat_C[312] <= 
//             mat_A[288] * mat_B[24] +
//             mat_A[289] * mat_B[56] +
//             mat_A[290] * mat_B[88] +
//             mat_A[291] * mat_B[120] +
//             mat_A[292] * mat_B[152] +
//             mat_A[293] * mat_B[184] +
//             mat_A[294] * mat_B[216] +
//             mat_A[295] * mat_B[248] +
//             mat_A[296] * mat_B[280] +
//             mat_A[297] * mat_B[312] +
//             mat_A[298] * mat_B[344] +
//             mat_A[299] * mat_B[376] +
//             mat_A[300] * mat_B[408] +
//             mat_A[301] * mat_B[440] +
//             mat_A[302] * mat_B[472] +
//             mat_A[303] * mat_B[504] +
//             mat_A[304] * mat_B[536] +
//             mat_A[305] * mat_B[568] +
//             mat_A[306] * mat_B[600] +
//             mat_A[307] * mat_B[632] +
//             mat_A[308] * mat_B[664] +
//             mat_A[309] * mat_B[696] +
//             mat_A[310] * mat_B[728] +
//             mat_A[311] * mat_B[760] +
//             mat_A[312] * mat_B[792] +
//             mat_A[313] * mat_B[824] +
//             mat_A[314] * mat_B[856] +
//             mat_A[315] * mat_B[888] +
//             mat_A[316] * mat_B[920] +
//             mat_A[317] * mat_B[952] +
//             mat_A[318] * mat_B[984] +
//             mat_A[319] * mat_B[1016];
//  mat_C[313] <= 
//             mat_A[288] * mat_B[25] +
//             mat_A[289] * mat_B[57] +
//             mat_A[290] * mat_B[89] +
//             mat_A[291] * mat_B[121] +
//             mat_A[292] * mat_B[153] +
//             mat_A[293] * mat_B[185] +
//             mat_A[294] * mat_B[217] +
//             mat_A[295] * mat_B[249] +
//             mat_A[296] * mat_B[281] +
//             mat_A[297] * mat_B[313] +
//             mat_A[298] * mat_B[345] +
//             mat_A[299] * mat_B[377] +
//             mat_A[300] * mat_B[409] +
//             mat_A[301] * mat_B[441] +
//             mat_A[302] * mat_B[473] +
//             mat_A[303] * mat_B[505] +
//             mat_A[304] * mat_B[537] +
//             mat_A[305] * mat_B[569] +
//             mat_A[306] * mat_B[601] +
//             mat_A[307] * mat_B[633] +
//             mat_A[308] * mat_B[665] +
//             mat_A[309] * mat_B[697] +
//             mat_A[310] * mat_B[729] +
//             mat_A[311] * mat_B[761] +
//             mat_A[312] * mat_B[793] +
//             mat_A[313] * mat_B[825] +
//             mat_A[314] * mat_B[857] +
//             mat_A[315] * mat_B[889] +
//             mat_A[316] * mat_B[921] +
//             mat_A[317] * mat_B[953] +
//             mat_A[318] * mat_B[985] +
//             mat_A[319] * mat_B[1017];
//  mat_C[314] <= 
//             mat_A[288] * mat_B[26] +
//             mat_A[289] * mat_B[58] +
//             mat_A[290] * mat_B[90] +
//             mat_A[291] * mat_B[122] +
//             mat_A[292] * mat_B[154] +
//             mat_A[293] * mat_B[186] +
//             mat_A[294] * mat_B[218] +
//             mat_A[295] * mat_B[250] +
//             mat_A[296] * mat_B[282] +
//             mat_A[297] * mat_B[314] +
//             mat_A[298] * mat_B[346] +
//             mat_A[299] * mat_B[378] +
//             mat_A[300] * mat_B[410] +
//             mat_A[301] * mat_B[442] +
//             mat_A[302] * mat_B[474] +
//             mat_A[303] * mat_B[506] +
//             mat_A[304] * mat_B[538] +
//             mat_A[305] * mat_B[570] +
//             mat_A[306] * mat_B[602] +
//             mat_A[307] * mat_B[634] +
//             mat_A[308] * mat_B[666] +
//             mat_A[309] * mat_B[698] +
//             mat_A[310] * mat_B[730] +
//             mat_A[311] * mat_B[762] +
//             mat_A[312] * mat_B[794] +
//             mat_A[313] * mat_B[826] +
//             mat_A[314] * mat_B[858] +
//             mat_A[315] * mat_B[890] +
//             mat_A[316] * mat_B[922] +
//             mat_A[317] * mat_B[954] +
//             mat_A[318] * mat_B[986] +
//             mat_A[319] * mat_B[1018];
//  mat_C[315] <= 
//             mat_A[288] * mat_B[27] +
//             mat_A[289] * mat_B[59] +
//             mat_A[290] * mat_B[91] +
//             mat_A[291] * mat_B[123] +
//             mat_A[292] * mat_B[155] +
//             mat_A[293] * mat_B[187] +
//             mat_A[294] * mat_B[219] +
//             mat_A[295] * mat_B[251] +
//             mat_A[296] * mat_B[283] +
//             mat_A[297] * mat_B[315] +
//             mat_A[298] * mat_B[347] +
//             mat_A[299] * mat_B[379] +
//             mat_A[300] * mat_B[411] +
//             mat_A[301] * mat_B[443] +
//             mat_A[302] * mat_B[475] +
//             mat_A[303] * mat_B[507] +
//             mat_A[304] * mat_B[539] +
//             mat_A[305] * mat_B[571] +
//             mat_A[306] * mat_B[603] +
//             mat_A[307] * mat_B[635] +
//             mat_A[308] * mat_B[667] +
//             mat_A[309] * mat_B[699] +
//             mat_A[310] * mat_B[731] +
//             mat_A[311] * mat_B[763] +
//             mat_A[312] * mat_B[795] +
//             mat_A[313] * mat_B[827] +
//             mat_A[314] * mat_B[859] +
//             mat_A[315] * mat_B[891] +
//             mat_A[316] * mat_B[923] +
//             mat_A[317] * mat_B[955] +
//             mat_A[318] * mat_B[987] +
//             mat_A[319] * mat_B[1019];
//  mat_C[316] <= 
//             mat_A[288] * mat_B[28] +
//             mat_A[289] * mat_B[60] +
//             mat_A[290] * mat_B[92] +
//             mat_A[291] * mat_B[124] +
//             mat_A[292] * mat_B[156] +
//             mat_A[293] * mat_B[188] +
//             mat_A[294] * mat_B[220] +
//             mat_A[295] * mat_B[252] +
//             mat_A[296] * mat_B[284] +
//             mat_A[297] * mat_B[316] +
//             mat_A[298] * mat_B[348] +
//             mat_A[299] * mat_B[380] +
//             mat_A[300] * mat_B[412] +
//             mat_A[301] * mat_B[444] +
//             mat_A[302] * mat_B[476] +
//             mat_A[303] * mat_B[508] +
//             mat_A[304] * mat_B[540] +
//             mat_A[305] * mat_B[572] +
//             mat_A[306] * mat_B[604] +
//             mat_A[307] * mat_B[636] +
//             mat_A[308] * mat_B[668] +
//             mat_A[309] * mat_B[700] +
//             mat_A[310] * mat_B[732] +
//             mat_A[311] * mat_B[764] +
//             mat_A[312] * mat_B[796] +
//             mat_A[313] * mat_B[828] +
//             mat_A[314] * mat_B[860] +
//             mat_A[315] * mat_B[892] +
//             mat_A[316] * mat_B[924] +
//             mat_A[317] * mat_B[956] +
//             mat_A[318] * mat_B[988] +
//             mat_A[319] * mat_B[1020];
//  mat_C[317] <= 
//             mat_A[288] * mat_B[29] +
//             mat_A[289] * mat_B[61] +
//             mat_A[290] * mat_B[93] +
//             mat_A[291] * mat_B[125] +
//             mat_A[292] * mat_B[157] +
//             mat_A[293] * mat_B[189] +
//             mat_A[294] * mat_B[221] +
//             mat_A[295] * mat_B[253] +
//             mat_A[296] * mat_B[285] +
//             mat_A[297] * mat_B[317] +
//             mat_A[298] * mat_B[349] +
//             mat_A[299] * mat_B[381] +
//             mat_A[300] * mat_B[413] +
//             mat_A[301] * mat_B[445] +
//             mat_A[302] * mat_B[477] +
//             mat_A[303] * mat_B[509] +
//             mat_A[304] * mat_B[541] +
//             mat_A[305] * mat_B[573] +
//             mat_A[306] * mat_B[605] +
//             mat_A[307] * mat_B[637] +
//             mat_A[308] * mat_B[669] +
//             mat_A[309] * mat_B[701] +
//             mat_A[310] * mat_B[733] +
//             mat_A[311] * mat_B[765] +
//             mat_A[312] * mat_B[797] +
//             mat_A[313] * mat_B[829] +
//             mat_A[314] * mat_B[861] +
//             mat_A[315] * mat_B[893] +
//             mat_A[316] * mat_B[925] +
//             mat_A[317] * mat_B[957] +
//             mat_A[318] * mat_B[989] +
//             mat_A[319] * mat_B[1021];
//  mat_C[318] <= 
//             mat_A[288] * mat_B[30] +
//             mat_A[289] * mat_B[62] +
//             mat_A[290] * mat_B[94] +
//             mat_A[291] * mat_B[126] +
//             mat_A[292] * mat_B[158] +
//             mat_A[293] * mat_B[190] +
//             mat_A[294] * mat_B[222] +
//             mat_A[295] * mat_B[254] +
//             mat_A[296] * mat_B[286] +
//             mat_A[297] * mat_B[318] +
//             mat_A[298] * mat_B[350] +
//             mat_A[299] * mat_B[382] +
//             mat_A[300] * mat_B[414] +
//             mat_A[301] * mat_B[446] +
//             mat_A[302] * mat_B[478] +
//             mat_A[303] * mat_B[510] +
//             mat_A[304] * mat_B[542] +
//             mat_A[305] * mat_B[574] +
//             mat_A[306] * mat_B[606] +
//             mat_A[307] * mat_B[638] +
//             mat_A[308] * mat_B[670] +
//             mat_A[309] * mat_B[702] +
//             mat_A[310] * mat_B[734] +
//             mat_A[311] * mat_B[766] +
//             mat_A[312] * mat_B[798] +
//             mat_A[313] * mat_B[830] +
//             mat_A[314] * mat_B[862] +
//             mat_A[315] * mat_B[894] +
//             mat_A[316] * mat_B[926] +
//             mat_A[317] * mat_B[958] +
//             mat_A[318] * mat_B[990] +
//             mat_A[319] * mat_B[1022];
//  mat_C[319] <= 
//             mat_A[288] * mat_B[31] +
//             mat_A[289] * mat_B[63] +
//             mat_A[290] * mat_B[95] +
//             mat_A[291] * mat_B[127] +
//             mat_A[292] * mat_B[159] +
//             mat_A[293] * mat_B[191] +
//             mat_A[294] * mat_B[223] +
//             mat_A[295] * mat_B[255] +
//             mat_A[296] * mat_B[287] +
//             mat_A[297] * mat_B[319] +
//             mat_A[298] * mat_B[351] +
//             mat_A[299] * mat_B[383] +
//             mat_A[300] * mat_B[415] +
//             mat_A[301] * mat_B[447] +
//             mat_A[302] * mat_B[479] +
//             mat_A[303] * mat_B[511] +
//             mat_A[304] * mat_B[543] +
//             mat_A[305] * mat_B[575] +
//             mat_A[306] * mat_B[607] +
//             mat_A[307] * mat_B[639] +
//             mat_A[308] * mat_B[671] +
//             mat_A[309] * mat_B[703] +
//             mat_A[310] * mat_B[735] +
//             mat_A[311] * mat_B[767] +
//             mat_A[312] * mat_B[799] +
//             mat_A[313] * mat_B[831] +
//             mat_A[314] * mat_B[863] +
//             mat_A[315] * mat_B[895] +
//             mat_A[316] * mat_B[927] +
//             mat_A[317] * mat_B[959] +
//             mat_A[318] * mat_B[991] +
//             mat_A[319] * mat_B[1023];
//  mat_C[320] <= 
//             mat_A[320] * mat_B[0] +
//             mat_A[321] * mat_B[32] +
//             mat_A[322] * mat_B[64] +
//             mat_A[323] * mat_B[96] +
//             mat_A[324] * mat_B[128] +
//             mat_A[325] * mat_B[160] +
//             mat_A[326] * mat_B[192] +
//             mat_A[327] * mat_B[224] +
//             mat_A[328] * mat_B[256] +
//             mat_A[329] * mat_B[288] +
//             mat_A[330] * mat_B[320] +
//             mat_A[331] * mat_B[352] +
//             mat_A[332] * mat_B[384] +
//             mat_A[333] * mat_B[416] +
//             mat_A[334] * mat_B[448] +
//             mat_A[335] * mat_B[480] +
//             mat_A[336] * mat_B[512] +
//             mat_A[337] * mat_B[544] +
//             mat_A[338] * mat_B[576] +
//             mat_A[339] * mat_B[608] +
//             mat_A[340] * mat_B[640] +
//             mat_A[341] * mat_B[672] +
//             mat_A[342] * mat_B[704] +
//             mat_A[343] * mat_B[736] +
//             mat_A[344] * mat_B[768] +
//             mat_A[345] * mat_B[800] +
//             mat_A[346] * mat_B[832] +
//             mat_A[347] * mat_B[864] +
//             mat_A[348] * mat_B[896] +
//             mat_A[349] * mat_B[928] +
//             mat_A[350] * mat_B[960] +
//             mat_A[351] * mat_B[992];
//  mat_C[321] <= 
//             mat_A[320] * mat_B[1] +
//             mat_A[321] * mat_B[33] +
//             mat_A[322] * mat_B[65] +
//             mat_A[323] * mat_B[97] +
//             mat_A[324] * mat_B[129] +
//             mat_A[325] * mat_B[161] +
//             mat_A[326] * mat_B[193] +
//             mat_A[327] * mat_B[225] +
//             mat_A[328] * mat_B[257] +
//             mat_A[329] * mat_B[289] +
//             mat_A[330] * mat_B[321] +
//             mat_A[331] * mat_B[353] +
//             mat_A[332] * mat_B[385] +
//             mat_A[333] * mat_B[417] +
//             mat_A[334] * mat_B[449] +
//             mat_A[335] * mat_B[481] +
//             mat_A[336] * mat_B[513] +
//             mat_A[337] * mat_B[545] +
//             mat_A[338] * mat_B[577] +
//             mat_A[339] * mat_B[609] +
//             mat_A[340] * mat_B[641] +
//             mat_A[341] * mat_B[673] +
//             mat_A[342] * mat_B[705] +
//             mat_A[343] * mat_B[737] +
//             mat_A[344] * mat_B[769] +
//             mat_A[345] * mat_B[801] +
//             mat_A[346] * mat_B[833] +
//             mat_A[347] * mat_B[865] +
//             mat_A[348] * mat_B[897] +
//             mat_A[349] * mat_B[929] +
//             mat_A[350] * mat_B[961] +
//             mat_A[351] * mat_B[993];
//  mat_C[322] <= 
//             mat_A[320] * mat_B[2] +
//             mat_A[321] * mat_B[34] +
//             mat_A[322] * mat_B[66] +
//             mat_A[323] * mat_B[98] +
//             mat_A[324] * mat_B[130] +
//             mat_A[325] * mat_B[162] +
//             mat_A[326] * mat_B[194] +
//             mat_A[327] * mat_B[226] +
//             mat_A[328] * mat_B[258] +
//             mat_A[329] * mat_B[290] +
//             mat_A[330] * mat_B[322] +
//             mat_A[331] * mat_B[354] +
//             mat_A[332] * mat_B[386] +
//             mat_A[333] * mat_B[418] +
//             mat_A[334] * mat_B[450] +
//             mat_A[335] * mat_B[482] +
//             mat_A[336] * mat_B[514] +
//             mat_A[337] * mat_B[546] +
//             mat_A[338] * mat_B[578] +
//             mat_A[339] * mat_B[610] +
//             mat_A[340] * mat_B[642] +
//             mat_A[341] * mat_B[674] +
//             mat_A[342] * mat_B[706] +
//             mat_A[343] * mat_B[738] +
//             mat_A[344] * mat_B[770] +
//             mat_A[345] * mat_B[802] +
//             mat_A[346] * mat_B[834] +
//             mat_A[347] * mat_B[866] +
//             mat_A[348] * mat_B[898] +
//             mat_A[349] * mat_B[930] +
//             mat_A[350] * mat_B[962] +
//             mat_A[351] * mat_B[994];
//  mat_C[323] <= 
//             mat_A[320] * mat_B[3] +
//             mat_A[321] * mat_B[35] +
//             mat_A[322] * mat_B[67] +
//             mat_A[323] * mat_B[99] +
//             mat_A[324] * mat_B[131] +
//             mat_A[325] * mat_B[163] +
//             mat_A[326] * mat_B[195] +
//             mat_A[327] * mat_B[227] +
//             mat_A[328] * mat_B[259] +
//             mat_A[329] * mat_B[291] +
//             mat_A[330] * mat_B[323] +
//             mat_A[331] * mat_B[355] +
//             mat_A[332] * mat_B[387] +
//             mat_A[333] * mat_B[419] +
//             mat_A[334] * mat_B[451] +
//             mat_A[335] * mat_B[483] +
//             mat_A[336] * mat_B[515] +
//             mat_A[337] * mat_B[547] +
//             mat_A[338] * mat_B[579] +
//             mat_A[339] * mat_B[611] +
//             mat_A[340] * mat_B[643] +
//             mat_A[341] * mat_B[675] +
//             mat_A[342] * mat_B[707] +
//             mat_A[343] * mat_B[739] +
//             mat_A[344] * mat_B[771] +
//             mat_A[345] * mat_B[803] +
//             mat_A[346] * mat_B[835] +
//             mat_A[347] * mat_B[867] +
//             mat_A[348] * mat_B[899] +
//             mat_A[349] * mat_B[931] +
//             mat_A[350] * mat_B[963] +
//             mat_A[351] * mat_B[995];
//  mat_C[324] <= 
//             mat_A[320] * mat_B[4] +
//             mat_A[321] * mat_B[36] +
//             mat_A[322] * mat_B[68] +
//             mat_A[323] * mat_B[100] +
//             mat_A[324] * mat_B[132] +
//             mat_A[325] * mat_B[164] +
//             mat_A[326] * mat_B[196] +
//             mat_A[327] * mat_B[228] +
//             mat_A[328] * mat_B[260] +
//             mat_A[329] * mat_B[292] +
//             mat_A[330] * mat_B[324] +
//             mat_A[331] * mat_B[356] +
//             mat_A[332] * mat_B[388] +
//             mat_A[333] * mat_B[420] +
//             mat_A[334] * mat_B[452] +
//             mat_A[335] * mat_B[484] +
//             mat_A[336] * mat_B[516] +
//             mat_A[337] * mat_B[548] +
//             mat_A[338] * mat_B[580] +
//             mat_A[339] * mat_B[612] +
//             mat_A[340] * mat_B[644] +
//             mat_A[341] * mat_B[676] +
//             mat_A[342] * mat_B[708] +
//             mat_A[343] * mat_B[740] +
//             mat_A[344] * mat_B[772] +
//             mat_A[345] * mat_B[804] +
//             mat_A[346] * mat_B[836] +
//             mat_A[347] * mat_B[868] +
//             mat_A[348] * mat_B[900] +
//             mat_A[349] * mat_B[932] +
//             mat_A[350] * mat_B[964] +
//             mat_A[351] * mat_B[996];
//  mat_C[325] <= 
//             mat_A[320] * mat_B[5] +
//             mat_A[321] * mat_B[37] +
//             mat_A[322] * mat_B[69] +
//             mat_A[323] * mat_B[101] +
//             mat_A[324] * mat_B[133] +
//             mat_A[325] * mat_B[165] +
//             mat_A[326] * mat_B[197] +
//             mat_A[327] * mat_B[229] +
//             mat_A[328] * mat_B[261] +
//             mat_A[329] * mat_B[293] +
//             mat_A[330] * mat_B[325] +
//             mat_A[331] * mat_B[357] +
//             mat_A[332] * mat_B[389] +
//             mat_A[333] * mat_B[421] +
//             mat_A[334] * mat_B[453] +
//             mat_A[335] * mat_B[485] +
//             mat_A[336] * mat_B[517] +
//             mat_A[337] * mat_B[549] +
//             mat_A[338] * mat_B[581] +
//             mat_A[339] * mat_B[613] +
//             mat_A[340] * mat_B[645] +
//             mat_A[341] * mat_B[677] +
//             mat_A[342] * mat_B[709] +
//             mat_A[343] * mat_B[741] +
//             mat_A[344] * mat_B[773] +
//             mat_A[345] * mat_B[805] +
//             mat_A[346] * mat_B[837] +
//             mat_A[347] * mat_B[869] +
//             mat_A[348] * mat_B[901] +
//             mat_A[349] * mat_B[933] +
//             mat_A[350] * mat_B[965] +
//             mat_A[351] * mat_B[997];
//  mat_C[326] <= 
//             mat_A[320] * mat_B[6] +
//             mat_A[321] * mat_B[38] +
//             mat_A[322] * mat_B[70] +
//             mat_A[323] * mat_B[102] +
//             mat_A[324] * mat_B[134] +
//             mat_A[325] * mat_B[166] +
//             mat_A[326] * mat_B[198] +
//             mat_A[327] * mat_B[230] +
//             mat_A[328] * mat_B[262] +
//             mat_A[329] * mat_B[294] +
//             mat_A[330] * mat_B[326] +
//             mat_A[331] * mat_B[358] +
//             mat_A[332] * mat_B[390] +
//             mat_A[333] * mat_B[422] +
//             mat_A[334] * mat_B[454] +
//             mat_A[335] * mat_B[486] +
//             mat_A[336] * mat_B[518] +
//             mat_A[337] * mat_B[550] +
//             mat_A[338] * mat_B[582] +
//             mat_A[339] * mat_B[614] +
//             mat_A[340] * mat_B[646] +
//             mat_A[341] * mat_B[678] +
//             mat_A[342] * mat_B[710] +
//             mat_A[343] * mat_B[742] +
//             mat_A[344] * mat_B[774] +
//             mat_A[345] * mat_B[806] +
//             mat_A[346] * mat_B[838] +
//             mat_A[347] * mat_B[870] +
//             mat_A[348] * mat_B[902] +
//             mat_A[349] * mat_B[934] +
//             mat_A[350] * mat_B[966] +
//             mat_A[351] * mat_B[998];
//  mat_C[327] <= 
//             mat_A[320] * mat_B[7] +
//             mat_A[321] * mat_B[39] +
//             mat_A[322] * mat_B[71] +
//             mat_A[323] * mat_B[103] +
//             mat_A[324] * mat_B[135] +
//             mat_A[325] * mat_B[167] +
//             mat_A[326] * mat_B[199] +
//             mat_A[327] * mat_B[231] +
//             mat_A[328] * mat_B[263] +
//             mat_A[329] * mat_B[295] +
//             mat_A[330] * mat_B[327] +
//             mat_A[331] * mat_B[359] +
//             mat_A[332] * mat_B[391] +
//             mat_A[333] * mat_B[423] +
//             mat_A[334] * mat_B[455] +
//             mat_A[335] * mat_B[487] +
//             mat_A[336] * mat_B[519] +
//             mat_A[337] * mat_B[551] +
//             mat_A[338] * mat_B[583] +
//             mat_A[339] * mat_B[615] +
//             mat_A[340] * mat_B[647] +
//             mat_A[341] * mat_B[679] +
//             mat_A[342] * mat_B[711] +
//             mat_A[343] * mat_B[743] +
//             mat_A[344] * mat_B[775] +
//             mat_A[345] * mat_B[807] +
//             mat_A[346] * mat_B[839] +
//             mat_A[347] * mat_B[871] +
//             mat_A[348] * mat_B[903] +
//             mat_A[349] * mat_B[935] +
//             mat_A[350] * mat_B[967] +
//             mat_A[351] * mat_B[999];
//  mat_C[328] <= 
//             mat_A[320] * mat_B[8] +
//             mat_A[321] * mat_B[40] +
//             mat_A[322] * mat_B[72] +
//             mat_A[323] * mat_B[104] +
//             mat_A[324] * mat_B[136] +
//             mat_A[325] * mat_B[168] +
//             mat_A[326] * mat_B[200] +
//             mat_A[327] * mat_B[232] +
//             mat_A[328] * mat_B[264] +
//             mat_A[329] * mat_B[296] +
//             mat_A[330] * mat_B[328] +
//             mat_A[331] * mat_B[360] +
//             mat_A[332] * mat_B[392] +
//             mat_A[333] * mat_B[424] +
//             mat_A[334] * mat_B[456] +
//             mat_A[335] * mat_B[488] +
//             mat_A[336] * mat_B[520] +
//             mat_A[337] * mat_B[552] +
//             mat_A[338] * mat_B[584] +
//             mat_A[339] * mat_B[616] +
//             mat_A[340] * mat_B[648] +
//             mat_A[341] * mat_B[680] +
//             mat_A[342] * mat_B[712] +
//             mat_A[343] * mat_B[744] +
//             mat_A[344] * mat_B[776] +
//             mat_A[345] * mat_B[808] +
//             mat_A[346] * mat_B[840] +
//             mat_A[347] * mat_B[872] +
//             mat_A[348] * mat_B[904] +
//             mat_A[349] * mat_B[936] +
//             mat_A[350] * mat_B[968] +
//             mat_A[351] * mat_B[1000];
//  mat_C[329] <= 
//             mat_A[320] * mat_B[9] +
//             mat_A[321] * mat_B[41] +
//             mat_A[322] * mat_B[73] +
//             mat_A[323] * mat_B[105] +
//             mat_A[324] * mat_B[137] +
//             mat_A[325] * mat_B[169] +
//             mat_A[326] * mat_B[201] +
//             mat_A[327] * mat_B[233] +
//             mat_A[328] * mat_B[265] +
//             mat_A[329] * mat_B[297] +
//             mat_A[330] * mat_B[329] +
//             mat_A[331] * mat_B[361] +
//             mat_A[332] * mat_B[393] +
//             mat_A[333] * mat_B[425] +
//             mat_A[334] * mat_B[457] +
//             mat_A[335] * mat_B[489] +
//             mat_A[336] * mat_B[521] +
//             mat_A[337] * mat_B[553] +
//             mat_A[338] * mat_B[585] +
//             mat_A[339] * mat_B[617] +
//             mat_A[340] * mat_B[649] +
//             mat_A[341] * mat_B[681] +
//             mat_A[342] * mat_B[713] +
//             mat_A[343] * mat_B[745] +
//             mat_A[344] * mat_B[777] +
//             mat_A[345] * mat_B[809] +
//             mat_A[346] * mat_B[841] +
//             mat_A[347] * mat_B[873] +
//             mat_A[348] * mat_B[905] +
//             mat_A[349] * mat_B[937] +
//             mat_A[350] * mat_B[969] +
//             mat_A[351] * mat_B[1001];
//  mat_C[330] <= 
//             mat_A[320] * mat_B[10] +
//             mat_A[321] * mat_B[42] +
//             mat_A[322] * mat_B[74] +
//             mat_A[323] * mat_B[106] +
//             mat_A[324] * mat_B[138] +
//             mat_A[325] * mat_B[170] +
//             mat_A[326] * mat_B[202] +
//             mat_A[327] * mat_B[234] +
//             mat_A[328] * mat_B[266] +
//             mat_A[329] * mat_B[298] +
//             mat_A[330] * mat_B[330] +
//             mat_A[331] * mat_B[362] +
//             mat_A[332] * mat_B[394] +
//             mat_A[333] * mat_B[426] +
//             mat_A[334] * mat_B[458] +
//             mat_A[335] * mat_B[490] +
//             mat_A[336] * mat_B[522] +
//             mat_A[337] * mat_B[554] +
//             mat_A[338] * mat_B[586] +
//             mat_A[339] * mat_B[618] +
//             mat_A[340] * mat_B[650] +
//             mat_A[341] * mat_B[682] +
//             mat_A[342] * mat_B[714] +
//             mat_A[343] * mat_B[746] +
//             mat_A[344] * mat_B[778] +
//             mat_A[345] * mat_B[810] +
//             mat_A[346] * mat_B[842] +
//             mat_A[347] * mat_B[874] +
//             mat_A[348] * mat_B[906] +
//             mat_A[349] * mat_B[938] +
//             mat_A[350] * mat_B[970] +
//             mat_A[351] * mat_B[1002];
//  mat_C[331] <= 
//             mat_A[320] * mat_B[11] +
//             mat_A[321] * mat_B[43] +
//             mat_A[322] * mat_B[75] +
//             mat_A[323] * mat_B[107] +
//             mat_A[324] * mat_B[139] +
//             mat_A[325] * mat_B[171] +
//             mat_A[326] * mat_B[203] +
//             mat_A[327] * mat_B[235] +
//             mat_A[328] * mat_B[267] +
//             mat_A[329] * mat_B[299] +
//             mat_A[330] * mat_B[331] +
//             mat_A[331] * mat_B[363] +
//             mat_A[332] * mat_B[395] +
//             mat_A[333] * mat_B[427] +
//             mat_A[334] * mat_B[459] +
//             mat_A[335] * mat_B[491] +
//             mat_A[336] * mat_B[523] +
//             mat_A[337] * mat_B[555] +
//             mat_A[338] * mat_B[587] +
//             mat_A[339] * mat_B[619] +
//             mat_A[340] * mat_B[651] +
//             mat_A[341] * mat_B[683] +
//             mat_A[342] * mat_B[715] +
//             mat_A[343] * mat_B[747] +
//             mat_A[344] * mat_B[779] +
//             mat_A[345] * mat_B[811] +
//             mat_A[346] * mat_B[843] +
//             mat_A[347] * mat_B[875] +
//             mat_A[348] * mat_B[907] +
//             mat_A[349] * mat_B[939] +
//             mat_A[350] * mat_B[971] +
//             mat_A[351] * mat_B[1003];
//  mat_C[332] <= 
//             mat_A[320] * mat_B[12] +
//             mat_A[321] * mat_B[44] +
//             mat_A[322] * mat_B[76] +
//             mat_A[323] * mat_B[108] +
//             mat_A[324] * mat_B[140] +
//             mat_A[325] * mat_B[172] +
//             mat_A[326] * mat_B[204] +
//             mat_A[327] * mat_B[236] +
//             mat_A[328] * mat_B[268] +
//             mat_A[329] * mat_B[300] +
//             mat_A[330] * mat_B[332] +
//             mat_A[331] * mat_B[364] +
//             mat_A[332] * mat_B[396] +
//             mat_A[333] * mat_B[428] +
//             mat_A[334] * mat_B[460] +
//             mat_A[335] * mat_B[492] +
//             mat_A[336] * mat_B[524] +
//             mat_A[337] * mat_B[556] +
//             mat_A[338] * mat_B[588] +
//             mat_A[339] * mat_B[620] +
//             mat_A[340] * mat_B[652] +
//             mat_A[341] * mat_B[684] +
//             mat_A[342] * mat_B[716] +
//             mat_A[343] * mat_B[748] +
//             mat_A[344] * mat_B[780] +
//             mat_A[345] * mat_B[812] +
//             mat_A[346] * mat_B[844] +
//             mat_A[347] * mat_B[876] +
//             mat_A[348] * mat_B[908] +
//             mat_A[349] * mat_B[940] +
//             mat_A[350] * mat_B[972] +
//             mat_A[351] * mat_B[1004];
//  mat_C[333] <= 
//             mat_A[320] * mat_B[13] +
//             mat_A[321] * mat_B[45] +
//             mat_A[322] * mat_B[77] +
//             mat_A[323] * mat_B[109] +
//             mat_A[324] * mat_B[141] +
//             mat_A[325] * mat_B[173] +
//             mat_A[326] * mat_B[205] +
//             mat_A[327] * mat_B[237] +
//             mat_A[328] * mat_B[269] +
//             mat_A[329] * mat_B[301] +
//             mat_A[330] * mat_B[333] +
//             mat_A[331] * mat_B[365] +
//             mat_A[332] * mat_B[397] +
//             mat_A[333] * mat_B[429] +
//             mat_A[334] * mat_B[461] +
//             mat_A[335] * mat_B[493] +
//             mat_A[336] * mat_B[525] +
//             mat_A[337] * mat_B[557] +
//             mat_A[338] * mat_B[589] +
//             mat_A[339] * mat_B[621] +
//             mat_A[340] * mat_B[653] +
//             mat_A[341] * mat_B[685] +
//             mat_A[342] * mat_B[717] +
//             mat_A[343] * mat_B[749] +
//             mat_A[344] * mat_B[781] +
//             mat_A[345] * mat_B[813] +
//             mat_A[346] * mat_B[845] +
//             mat_A[347] * mat_B[877] +
//             mat_A[348] * mat_B[909] +
//             mat_A[349] * mat_B[941] +
//             mat_A[350] * mat_B[973] +
//             mat_A[351] * mat_B[1005];
//  mat_C[334] <= 
//             mat_A[320] * mat_B[14] +
//             mat_A[321] * mat_B[46] +
//             mat_A[322] * mat_B[78] +
//             mat_A[323] * mat_B[110] +
//             mat_A[324] * mat_B[142] +
//             mat_A[325] * mat_B[174] +
//             mat_A[326] * mat_B[206] +
//             mat_A[327] * mat_B[238] +
//             mat_A[328] * mat_B[270] +
//             mat_A[329] * mat_B[302] +
//             mat_A[330] * mat_B[334] +
//             mat_A[331] * mat_B[366] +
//             mat_A[332] * mat_B[398] +
//             mat_A[333] * mat_B[430] +
//             mat_A[334] * mat_B[462] +
//             mat_A[335] * mat_B[494] +
//             mat_A[336] * mat_B[526] +
//             mat_A[337] * mat_B[558] +
//             mat_A[338] * mat_B[590] +
//             mat_A[339] * mat_B[622] +
//             mat_A[340] * mat_B[654] +
//             mat_A[341] * mat_B[686] +
//             mat_A[342] * mat_B[718] +
//             mat_A[343] * mat_B[750] +
//             mat_A[344] * mat_B[782] +
//             mat_A[345] * mat_B[814] +
//             mat_A[346] * mat_B[846] +
//             mat_A[347] * mat_B[878] +
//             mat_A[348] * mat_B[910] +
//             mat_A[349] * mat_B[942] +
//             mat_A[350] * mat_B[974] +
//             mat_A[351] * mat_B[1006];
//  mat_C[335] <= 
//             mat_A[320] * mat_B[15] +
//             mat_A[321] * mat_B[47] +
//             mat_A[322] * mat_B[79] +
//             mat_A[323] * mat_B[111] +
//             mat_A[324] * mat_B[143] +
//             mat_A[325] * mat_B[175] +
//             mat_A[326] * mat_B[207] +
//             mat_A[327] * mat_B[239] +
//             mat_A[328] * mat_B[271] +
//             mat_A[329] * mat_B[303] +
//             mat_A[330] * mat_B[335] +
//             mat_A[331] * mat_B[367] +
//             mat_A[332] * mat_B[399] +
//             mat_A[333] * mat_B[431] +
//             mat_A[334] * mat_B[463] +
//             mat_A[335] * mat_B[495] +
//             mat_A[336] * mat_B[527] +
//             mat_A[337] * mat_B[559] +
//             mat_A[338] * mat_B[591] +
//             mat_A[339] * mat_B[623] +
//             mat_A[340] * mat_B[655] +
//             mat_A[341] * mat_B[687] +
//             mat_A[342] * mat_B[719] +
//             mat_A[343] * mat_B[751] +
//             mat_A[344] * mat_B[783] +
//             mat_A[345] * mat_B[815] +
//             mat_A[346] * mat_B[847] +
//             mat_A[347] * mat_B[879] +
//             mat_A[348] * mat_B[911] +
//             mat_A[349] * mat_B[943] +
//             mat_A[350] * mat_B[975] +
//             mat_A[351] * mat_B[1007];
//  mat_C[336] <= 
//             mat_A[320] * mat_B[16] +
//             mat_A[321] * mat_B[48] +
//             mat_A[322] * mat_B[80] +
//             mat_A[323] * mat_B[112] +
//             mat_A[324] * mat_B[144] +
//             mat_A[325] * mat_B[176] +
//             mat_A[326] * mat_B[208] +
//             mat_A[327] * mat_B[240] +
//             mat_A[328] * mat_B[272] +
//             mat_A[329] * mat_B[304] +
//             mat_A[330] * mat_B[336] +
//             mat_A[331] * mat_B[368] +
//             mat_A[332] * mat_B[400] +
//             mat_A[333] * mat_B[432] +
//             mat_A[334] * mat_B[464] +
//             mat_A[335] * mat_B[496] +
//             mat_A[336] * mat_B[528] +
//             mat_A[337] * mat_B[560] +
//             mat_A[338] * mat_B[592] +
//             mat_A[339] * mat_B[624] +
//             mat_A[340] * mat_B[656] +
//             mat_A[341] * mat_B[688] +
//             mat_A[342] * mat_B[720] +
//             mat_A[343] * mat_B[752] +
//             mat_A[344] * mat_B[784] +
//             mat_A[345] * mat_B[816] +
//             mat_A[346] * mat_B[848] +
//             mat_A[347] * mat_B[880] +
//             mat_A[348] * mat_B[912] +
//             mat_A[349] * mat_B[944] +
//             mat_A[350] * mat_B[976] +
//             mat_A[351] * mat_B[1008];
//  mat_C[337] <= 
//             mat_A[320] * mat_B[17] +
//             mat_A[321] * mat_B[49] +
//             mat_A[322] * mat_B[81] +
//             mat_A[323] * mat_B[113] +
//             mat_A[324] * mat_B[145] +
//             mat_A[325] * mat_B[177] +
//             mat_A[326] * mat_B[209] +
//             mat_A[327] * mat_B[241] +
//             mat_A[328] * mat_B[273] +
//             mat_A[329] * mat_B[305] +
//             mat_A[330] * mat_B[337] +
//             mat_A[331] * mat_B[369] +
//             mat_A[332] * mat_B[401] +
//             mat_A[333] * mat_B[433] +
//             mat_A[334] * mat_B[465] +
//             mat_A[335] * mat_B[497] +
//             mat_A[336] * mat_B[529] +
//             mat_A[337] * mat_B[561] +
//             mat_A[338] * mat_B[593] +
//             mat_A[339] * mat_B[625] +
//             mat_A[340] * mat_B[657] +
//             mat_A[341] * mat_B[689] +
//             mat_A[342] * mat_B[721] +
//             mat_A[343] * mat_B[753] +
//             mat_A[344] * mat_B[785] +
//             mat_A[345] * mat_B[817] +
//             mat_A[346] * mat_B[849] +
//             mat_A[347] * mat_B[881] +
//             mat_A[348] * mat_B[913] +
//             mat_A[349] * mat_B[945] +
//             mat_A[350] * mat_B[977] +
//             mat_A[351] * mat_B[1009];
//  mat_C[338] <= 
//             mat_A[320] * mat_B[18] +
//             mat_A[321] * mat_B[50] +
//             mat_A[322] * mat_B[82] +
//             mat_A[323] * mat_B[114] +
//             mat_A[324] * mat_B[146] +
//             mat_A[325] * mat_B[178] +
//             mat_A[326] * mat_B[210] +
//             mat_A[327] * mat_B[242] +
//             mat_A[328] * mat_B[274] +
//             mat_A[329] * mat_B[306] +
//             mat_A[330] * mat_B[338] +
//             mat_A[331] * mat_B[370] +
//             mat_A[332] * mat_B[402] +
//             mat_A[333] * mat_B[434] +
//             mat_A[334] * mat_B[466] +
//             mat_A[335] * mat_B[498] +
//             mat_A[336] * mat_B[530] +
//             mat_A[337] * mat_B[562] +
//             mat_A[338] * mat_B[594] +
//             mat_A[339] * mat_B[626] +
//             mat_A[340] * mat_B[658] +
//             mat_A[341] * mat_B[690] +
//             mat_A[342] * mat_B[722] +
//             mat_A[343] * mat_B[754] +
//             mat_A[344] * mat_B[786] +
//             mat_A[345] * mat_B[818] +
//             mat_A[346] * mat_B[850] +
//             mat_A[347] * mat_B[882] +
//             mat_A[348] * mat_B[914] +
//             mat_A[349] * mat_B[946] +
//             mat_A[350] * mat_B[978] +
//             mat_A[351] * mat_B[1010];
//  mat_C[339] <= 
//             mat_A[320] * mat_B[19] +
//             mat_A[321] * mat_B[51] +
//             mat_A[322] * mat_B[83] +
//             mat_A[323] * mat_B[115] +
//             mat_A[324] * mat_B[147] +
//             mat_A[325] * mat_B[179] +
//             mat_A[326] * mat_B[211] +
//             mat_A[327] * mat_B[243] +
//             mat_A[328] * mat_B[275] +
//             mat_A[329] * mat_B[307] +
//             mat_A[330] * mat_B[339] +
//             mat_A[331] * mat_B[371] +
//             mat_A[332] * mat_B[403] +
//             mat_A[333] * mat_B[435] +
//             mat_A[334] * mat_B[467] +
//             mat_A[335] * mat_B[499] +
//             mat_A[336] * mat_B[531] +
//             mat_A[337] * mat_B[563] +
//             mat_A[338] * mat_B[595] +
//             mat_A[339] * mat_B[627] +
//             mat_A[340] * mat_B[659] +
//             mat_A[341] * mat_B[691] +
//             mat_A[342] * mat_B[723] +
//             mat_A[343] * mat_B[755] +
//             mat_A[344] * mat_B[787] +
//             mat_A[345] * mat_B[819] +
//             mat_A[346] * mat_B[851] +
//             mat_A[347] * mat_B[883] +
//             mat_A[348] * mat_B[915] +
//             mat_A[349] * mat_B[947] +
//             mat_A[350] * mat_B[979] +
//             mat_A[351] * mat_B[1011];
//  mat_C[340] <= 
//             mat_A[320] * mat_B[20] +
//             mat_A[321] * mat_B[52] +
//             mat_A[322] * mat_B[84] +
//             mat_A[323] * mat_B[116] +
//             mat_A[324] * mat_B[148] +
//             mat_A[325] * mat_B[180] +
//             mat_A[326] * mat_B[212] +
//             mat_A[327] * mat_B[244] +
//             mat_A[328] * mat_B[276] +
//             mat_A[329] * mat_B[308] +
//             mat_A[330] * mat_B[340] +
//             mat_A[331] * mat_B[372] +
//             mat_A[332] * mat_B[404] +
//             mat_A[333] * mat_B[436] +
//             mat_A[334] * mat_B[468] +
//             mat_A[335] * mat_B[500] +
//             mat_A[336] * mat_B[532] +
//             mat_A[337] * mat_B[564] +
//             mat_A[338] * mat_B[596] +
//             mat_A[339] * mat_B[628] +
//             mat_A[340] * mat_B[660] +
//             mat_A[341] * mat_B[692] +
//             mat_A[342] * mat_B[724] +
//             mat_A[343] * mat_B[756] +
//             mat_A[344] * mat_B[788] +
//             mat_A[345] * mat_B[820] +
//             mat_A[346] * mat_B[852] +
//             mat_A[347] * mat_B[884] +
//             mat_A[348] * mat_B[916] +
//             mat_A[349] * mat_B[948] +
//             mat_A[350] * mat_B[980] +
//             mat_A[351] * mat_B[1012];
//  mat_C[341] <= 
//             mat_A[320] * mat_B[21] +
//             mat_A[321] * mat_B[53] +
//             mat_A[322] * mat_B[85] +
//             mat_A[323] * mat_B[117] +
//             mat_A[324] * mat_B[149] +
//             mat_A[325] * mat_B[181] +
//             mat_A[326] * mat_B[213] +
//             mat_A[327] * mat_B[245] +
//             mat_A[328] * mat_B[277] +
//             mat_A[329] * mat_B[309] +
//             mat_A[330] * mat_B[341] +
//             mat_A[331] * mat_B[373] +
//             mat_A[332] * mat_B[405] +
//             mat_A[333] * mat_B[437] +
//             mat_A[334] * mat_B[469] +
//             mat_A[335] * mat_B[501] +
//             mat_A[336] * mat_B[533] +
//             mat_A[337] * mat_B[565] +
//             mat_A[338] * mat_B[597] +
//             mat_A[339] * mat_B[629] +
//             mat_A[340] * mat_B[661] +
//             mat_A[341] * mat_B[693] +
//             mat_A[342] * mat_B[725] +
//             mat_A[343] * mat_B[757] +
//             mat_A[344] * mat_B[789] +
//             mat_A[345] * mat_B[821] +
//             mat_A[346] * mat_B[853] +
//             mat_A[347] * mat_B[885] +
//             mat_A[348] * mat_B[917] +
//             mat_A[349] * mat_B[949] +
//             mat_A[350] * mat_B[981] +
//             mat_A[351] * mat_B[1013];
//  mat_C[342] <= 
//             mat_A[320] * mat_B[22] +
//             mat_A[321] * mat_B[54] +
//             mat_A[322] * mat_B[86] +
//             mat_A[323] * mat_B[118] +
//             mat_A[324] * mat_B[150] +
//             mat_A[325] * mat_B[182] +
//             mat_A[326] * mat_B[214] +
//             mat_A[327] * mat_B[246] +
//             mat_A[328] * mat_B[278] +
//             mat_A[329] * mat_B[310] +
//             mat_A[330] * mat_B[342] +
//             mat_A[331] * mat_B[374] +
//             mat_A[332] * mat_B[406] +
//             mat_A[333] * mat_B[438] +
//             mat_A[334] * mat_B[470] +
//             mat_A[335] * mat_B[502] +
//             mat_A[336] * mat_B[534] +
//             mat_A[337] * mat_B[566] +
//             mat_A[338] * mat_B[598] +
//             mat_A[339] * mat_B[630] +
//             mat_A[340] * mat_B[662] +
//             mat_A[341] * mat_B[694] +
//             mat_A[342] * mat_B[726] +
//             mat_A[343] * mat_B[758] +
//             mat_A[344] * mat_B[790] +
//             mat_A[345] * mat_B[822] +
//             mat_A[346] * mat_B[854] +
//             mat_A[347] * mat_B[886] +
//             mat_A[348] * mat_B[918] +
//             mat_A[349] * mat_B[950] +
//             mat_A[350] * mat_B[982] +
//             mat_A[351] * mat_B[1014];
//  mat_C[343] <= 
//             mat_A[320] * mat_B[23] +
//             mat_A[321] * mat_B[55] +
//             mat_A[322] * mat_B[87] +
//             mat_A[323] * mat_B[119] +
//             mat_A[324] * mat_B[151] +
//             mat_A[325] * mat_B[183] +
//             mat_A[326] * mat_B[215] +
//             mat_A[327] * mat_B[247] +
//             mat_A[328] * mat_B[279] +
//             mat_A[329] * mat_B[311] +
//             mat_A[330] * mat_B[343] +
//             mat_A[331] * mat_B[375] +
//             mat_A[332] * mat_B[407] +
//             mat_A[333] * mat_B[439] +
//             mat_A[334] * mat_B[471] +
//             mat_A[335] * mat_B[503] +
//             mat_A[336] * mat_B[535] +
//             mat_A[337] * mat_B[567] +
//             mat_A[338] * mat_B[599] +
//             mat_A[339] * mat_B[631] +
//             mat_A[340] * mat_B[663] +
//             mat_A[341] * mat_B[695] +
//             mat_A[342] * mat_B[727] +
//             mat_A[343] * mat_B[759] +
//             mat_A[344] * mat_B[791] +
//             mat_A[345] * mat_B[823] +
//             mat_A[346] * mat_B[855] +
//             mat_A[347] * mat_B[887] +
//             mat_A[348] * mat_B[919] +
//             mat_A[349] * mat_B[951] +
//             mat_A[350] * mat_B[983] +
//             mat_A[351] * mat_B[1015];
//  mat_C[344] <= 
//             mat_A[320] * mat_B[24] +
//             mat_A[321] * mat_B[56] +
//             mat_A[322] * mat_B[88] +
//             mat_A[323] * mat_B[120] +
//             mat_A[324] * mat_B[152] +
//             mat_A[325] * mat_B[184] +
//             mat_A[326] * mat_B[216] +
//             mat_A[327] * mat_B[248] +
//             mat_A[328] * mat_B[280] +
//             mat_A[329] * mat_B[312] +
//             mat_A[330] * mat_B[344] +
//             mat_A[331] * mat_B[376] +
//             mat_A[332] * mat_B[408] +
//             mat_A[333] * mat_B[440] +
//             mat_A[334] * mat_B[472] +
//             mat_A[335] * mat_B[504] +
//             mat_A[336] * mat_B[536] +
//             mat_A[337] * mat_B[568] +
//             mat_A[338] * mat_B[600] +
//             mat_A[339] * mat_B[632] +
//             mat_A[340] * mat_B[664] +
//             mat_A[341] * mat_B[696] +
//             mat_A[342] * mat_B[728] +
//             mat_A[343] * mat_B[760] +
//             mat_A[344] * mat_B[792] +
//             mat_A[345] * mat_B[824] +
//             mat_A[346] * mat_B[856] +
//             mat_A[347] * mat_B[888] +
//             mat_A[348] * mat_B[920] +
//             mat_A[349] * mat_B[952] +
//             mat_A[350] * mat_B[984] +
//             mat_A[351] * mat_B[1016];
//  mat_C[345] <= 
//             mat_A[320] * mat_B[25] +
//             mat_A[321] * mat_B[57] +
//             mat_A[322] * mat_B[89] +
//             mat_A[323] * mat_B[121] +
//             mat_A[324] * mat_B[153] +
//             mat_A[325] * mat_B[185] +
//             mat_A[326] * mat_B[217] +
//             mat_A[327] * mat_B[249] +
//             mat_A[328] * mat_B[281] +
//             mat_A[329] * mat_B[313] +
//             mat_A[330] * mat_B[345] +
//             mat_A[331] * mat_B[377] +
//             mat_A[332] * mat_B[409] +
//             mat_A[333] * mat_B[441] +
//             mat_A[334] * mat_B[473] +
//             mat_A[335] * mat_B[505] +
//             mat_A[336] * mat_B[537] +
//             mat_A[337] * mat_B[569] +
//             mat_A[338] * mat_B[601] +
//             mat_A[339] * mat_B[633] +
//             mat_A[340] * mat_B[665] +
//             mat_A[341] * mat_B[697] +
//             mat_A[342] * mat_B[729] +
//             mat_A[343] * mat_B[761] +
//             mat_A[344] * mat_B[793] +
//             mat_A[345] * mat_B[825] +
//             mat_A[346] * mat_B[857] +
//             mat_A[347] * mat_B[889] +
//             mat_A[348] * mat_B[921] +
//             mat_A[349] * mat_B[953] +
//             mat_A[350] * mat_B[985] +
//             mat_A[351] * mat_B[1017];
//  mat_C[346] <= 
//             mat_A[320] * mat_B[26] +
//             mat_A[321] * mat_B[58] +
//             mat_A[322] * mat_B[90] +
//             mat_A[323] * mat_B[122] +
//             mat_A[324] * mat_B[154] +
//             mat_A[325] * mat_B[186] +
//             mat_A[326] * mat_B[218] +
//             mat_A[327] * mat_B[250] +
//             mat_A[328] * mat_B[282] +
//             mat_A[329] * mat_B[314] +
//             mat_A[330] * mat_B[346] +
//             mat_A[331] * mat_B[378] +
//             mat_A[332] * mat_B[410] +
//             mat_A[333] * mat_B[442] +
//             mat_A[334] * mat_B[474] +
//             mat_A[335] * mat_B[506] +
//             mat_A[336] * mat_B[538] +
//             mat_A[337] * mat_B[570] +
//             mat_A[338] * mat_B[602] +
//             mat_A[339] * mat_B[634] +
//             mat_A[340] * mat_B[666] +
//             mat_A[341] * mat_B[698] +
//             mat_A[342] * mat_B[730] +
//             mat_A[343] * mat_B[762] +
//             mat_A[344] * mat_B[794] +
//             mat_A[345] * mat_B[826] +
//             mat_A[346] * mat_B[858] +
//             mat_A[347] * mat_B[890] +
//             mat_A[348] * mat_B[922] +
//             mat_A[349] * mat_B[954] +
//             mat_A[350] * mat_B[986] +
//             mat_A[351] * mat_B[1018];
//  mat_C[347] <= 
//             mat_A[320] * mat_B[27] +
//             mat_A[321] * mat_B[59] +
//             mat_A[322] * mat_B[91] +
//             mat_A[323] * mat_B[123] +
//             mat_A[324] * mat_B[155] +
//             mat_A[325] * mat_B[187] +
//             mat_A[326] * mat_B[219] +
//             mat_A[327] * mat_B[251] +
//             mat_A[328] * mat_B[283] +
//             mat_A[329] * mat_B[315] +
//             mat_A[330] * mat_B[347] +
//             mat_A[331] * mat_B[379] +
//             mat_A[332] * mat_B[411] +
//             mat_A[333] * mat_B[443] +
//             mat_A[334] * mat_B[475] +
//             mat_A[335] * mat_B[507] +
//             mat_A[336] * mat_B[539] +
//             mat_A[337] * mat_B[571] +
//             mat_A[338] * mat_B[603] +
//             mat_A[339] * mat_B[635] +
//             mat_A[340] * mat_B[667] +
//             mat_A[341] * mat_B[699] +
//             mat_A[342] * mat_B[731] +
//             mat_A[343] * mat_B[763] +
//             mat_A[344] * mat_B[795] +
//             mat_A[345] * mat_B[827] +
//             mat_A[346] * mat_B[859] +
//             mat_A[347] * mat_B[891] +
//             mat_A[348] * mat_B[923] +
//             mat_A[349] * mat_B[955] +
//             mat_A[350] * mat_B[987] +
//             mat_A[351] * mat_B[1019];
//  mat_C[348] <= 
//             mat_A[320] * mat_B[28] +
//             mat_A[321] * mat_B[60] +
//             mat_A[322] * mat_B[92] +
//             mat_A[323] * mat_B[124] +
//             mat_A[324] * mat_B[156] +
//             mat_A[325] * mat_B[188] +
//             mat_A[326] * mat_B[220] +
//             mat_A[327] * mat_B[252] +
//             mat_A[328] * mat_B[284] +
//             mat_A[329] * mat_B[316] +
//             mat_A[330] * mat_B[348] +
//             mat_A[331] * mat_B[380] +
//             mat_A[332] * mat_B[412] +
//             mat_A[333] * mat_B[444] +
//             mat_A[334] * mat_B[476] +
//             mat_A[335] * mat_B[508] +
//             mat_A[336] * mat_B[540] +
//             mat_A[337] * mat_B[572] +
//             mat_A[338] * mat_B[604] +
//             mat_A[339] * mat_B[636] +
//             mat_A[340] * mat_B[668] +
//             mat_A[341] * mat_B[700] +
//             mat_A[342] * mat_B[732] +
//             mat_A[343] * mat_B[764] +
//             mat_A[344] * mat_B[796] +
//             mat_A[345] * mat_B[828] +
//             mat_A[346] * mat_B[860] +
//             mat_A[347] * mat_B[892] +
//             mat_A[348] * mat_B[924] +
//             mat_A[349] * mat_B[956] +
//             mat_A[350] * mat_B[988] +
//             mat_A[351] * mat_B[1020];
//  mat_C[349] <= 
//             mat_A[320] * mat_B[29] +
//             mat_A[321] * mat_B[61] +
//             mat_A[322] * mat_B[93] +
//             mat_A[323] * mat_B[125] +
//             mat_A[324] * mat_B[157] +
//             mat_A[325] * mat_B[189] +
//             mat_A[326] * mat_B[221] +
//             mat_A[327] * mat_B[253] +
//             mat_A[328] * mat_B[285] +
//             mat_A[329] * mat_B[317] +
//             mat_A[330] * mat_B[349] +
//             mat_A[331] * mat_B[381] +
//             mat_A[332] * mat_B[413] +
//             mat_A[333] * mat_B[445] +
//             mat_A[334] * mat_B[477] +
//             mat_A[335] * mat_B[509] +
//             mat_A[336] * mat_B[541] +
//             mat_A[337] * mat_B[573] +
//             mat_A[338] * mat_B[605] +
//             mat_A[339] * mat_B[637] +
//             mat_A[340] * mat_B[669] +
//             mat_A[341] * mat_B[701] +
//             mat_A[342] * mat_B[733] +
//             mat_A[343] * mat_B[765] +
//             mat_A[344] * mat_B[797] +
//             mat_A[345] * mat_B[829] +
//             mat_A[346] * mat_B[861] +
//             mat_A[347] * mat_B[893] +
//             mat_A[348] * mat_B[925] +
//             mat_A[349] * mat_B[957] +
//             mat_A[350] * mat_B[989] +
//             mat_A[351] * mat_B[1021];
//  mat_C[350] <= 
//             mat_A[320] * mat_B[30] +
//             mat_A[321] * mat_B[62] +
//             mat_A[322] * mat_B[94] +
//             mat_A[323] * mat_B[126] +
//             mat_A[324] * mat_B[158] +
//             mat_A[325] * mat_B[190] +
//             mat_A[326] * mat_B[222] +
//             mat_A[327] * mat_B[254] +
//             mat_A[328] * mat_B[286] +
//             mat_A[329] * mat_B[318] +
//             mat_A[330] * mat_B[350] +
//             mat_A[331] * mat_B[382] +
//             mat_A[332] * mat_B[414] +
//             mat_A[333] * mat_B[446] +
//             mat_A[334] * mat_B[478] +
//             mat_A[335] * mat_B[510] +
//             mat_A[336] * mat_B[542] +
//             mat_A[337] * mat_B[574] +
//             mat_A[338] * mat_B[606] +
//             mat_A[339] * mat_B[638] +
//             mat_A[340] * mat_B[670] +
//             mat_A[341] * mat_B[702] +
//             mat_A[342] * mat_B[734] +
//             mat_A[343] * mat_B[766] +
//             mat_A[344] * mat_B[798] +
//             mat_A[345] * mat_B[830] +
//             mat_A[346] * mat_B[862] +
//             mat_A[347] * mat_B[894] +
//             mat_A[348] * mat_B[926] +
//             mat_A[349] * mat_B[958] +
//             mat_A[350] * mat_B[990] +
//             mat_A[351] * mat_B[1022];
//  mat_C[351] <= 
//             mat_A[320] * mat_B[31] +
//             mat_A[321] * mat_B[63] +
//             mat_A[322] * mat_B[95] +
//             mat_A[323] * mat_B[127] +
//             mat_A[324] * mat_B[159] +
//             mat_A[325] * mat_B[191] +
//             mat_A[326] * mat_B[223] +
//             mat_A[327] * mat_B[255] +
//             mat_A[328] * mat_B[287] +
//             mat_A[329] * mat_B[319] +
//             mat_A[330] * mat_B[351] +
//             mat_A[331] * mat_B[383] +
//             mat_A[332] * mat_B[415] +
//             mat_A[333] * mat_B[447] +
//             mat_A[334] * mat_B[479] +
//             mat_A[335] * mat_B[511] +
//             mat_A[336] * mat_B[543] +
//             mat_A[337] * mat_B[575] +
//             mat_A[338] * mat_B[607] +
//             mat_A[339] * mat_B[639] +
//             mat_A[340] * mat_B[671] +
//             mat_A[341] * mat_B[703] +
//             mat_A[342] * mat_B[735] +
//             mat_A[343] * mat_B[767] +
//             mat_A[344] * mat_B[799] +
//             mat_A[345] * mat_B[831] +
//             mat_A[346] * mat_B[863] +
//             mat_A[347] * mat_B[895] +
//             mat_A[348] * mat_B[927] +
//             mat_A[349] * mat_B[959] +
//             mat_A[350] * mat_B[991] +
//             mat_A[351] * mat_B[1023];
//  mat_C[352] <= 
//             mat_A[352] * mat_B[0] +
//             mat_A[353] * mat_B[32] +
//             mat_A[354] * mat_B[64] +
//             mat_A[355] * mat_B[96] +
//             mat_A[356] * mat_B[128] +
//             mat_A[357] * mat_B[160] +
//             mat_A[358] * mat_B[192] +
//             mat_A[359] * mat_B[224] +
//             mat_A[360] * mat_B[256] +
//             mat_A[361] * mat_B[288] +
//             mat_A[362] * mat_B[320] +
//             mat_A[363] * mat_B[352] +
//             mat_A[364] * mat_B[384] +
//             mat_A[365] * mat_B[416] +
//             mat_A[366] * mat_B[448] +
//             mat_A[367] * mat_B[480] +
//             mat_A[368] * mat_B[512] +
//             mat_A[369] * mat_B[544] +
//             mat_A[370] * mat_B[576] +
//             mat_A[371] * mat_B[608] +
//             mat_A[372] * mat_B[640] +
//             mat_A[373] * mat_B[672] +
//             mat_A[374] * mat_B[704] +
//             mat_A[375] * mat_B[736] +
//             mat_A[376] * mat_B[768] +
//             mat_A[377] * mat_B[800] +
//             mat_A[378] * mat_B[832] +
//             mat_A[379] * mat_B[864] +
//             mat_A[380] * mat_B[896] +
//             mat_A[381] * mat_B[928] +
//             mat_A[382] * mat_B[960] +
//             mat_A[383] * mat_B[992];
//  mat_C[353] <= 
//             mat_A[352] * mat_B[1] +
//             mat_A[353] * mat_B[33] +
//             mat_A[354] * mat_B[65] +
//             mat_A[355] * mat_B[97] +
//             mat_A[356] * mat_B[129] +
//             mat_A[357] * mat_B[161] +
//             mat_A[358] * mat_B[193] +
//             mat_A[359] * mat_B[225] +
//             mat_A[360] * mat_B[257] +
//             mat_A[361] * mat_B[289] +
//             mat_A[362] * mat_B[321] +
//             mat_A[363] * mat_B[353] +
//             mat_A[364] * mat_B[385] +
//             mat_A[365] * mat_B[417] +
//             mat_A[366] * mat_B[449] +
//             mat_A[367] * mat_B[481] +
//             mat_A[368] * mat_B[513] +
//             mat_A[369] * mat_B[545] +
//             mat_A[370] * mat_B[577] +
//             mat_A[371] * mat_B[609] +
//             mat_A[372] * mat_B[641] +
//             mat_A[373] * mat_B[673] +
//             mat_A[374] * mat_B[705] +
//             mat_A[375] * mat_B[737] +
//             mat_A[376] * mat_B[769] +
//             mat_A[377] * mat_B[801] +
//             mat_A[378] * mat_B[833] +
//             mat_A[379] * mat_B[865] +
//             mat_A[380] * mat_B[897] +
//             mat_A[381] * mat_B[929] +
//             mat_A[382] * mat_B[961] +
//             mat_A[383] * mat_B[993];
//  mat_C[354] <= 
//             mat_A[352] * mat_B[2] +
//             mat_A[353] * mat_B[34] +
//             mat_A[354] * mat_B[66] +
//             mat_A[355] * mat_B[98] +
//             mat_A[356] * mat_B[130] +
//             mat_A[357] * mat_B[162] +
//             mat_A[358] * mat_B[194] +
//             mat_A[359] * mat_B[226] +
//             mat_A[360] * mat_B[258] +
//             mat_A[361] * mat_B[290] +
//             mat_A[362] * mat_B[322] +
//             mat_A[363] * mat_B[354] +
//             mat_A[364] * mat_B[386] +
//             mat_A[365] * mat_B[418] +
//             mat_A[366] * mat_B[450] +
//             mat_A[367] * mat_B[482] +
//             mat_A[368] * mat_B[514] +
//             mat_A[369] * mat_B[546] +
//             mat_A[370] * mat_B[578] +
//             mat_A[371] * mat_B[610] +
//             mat_A[372] * mat_B[642] +
//             mat_A[373] * mat_B[674] +
//             mat_A[374] * mat_B[706] +
//             mat_A[375] * mat_B[738] +
//             mat_A[376] * mat_B[770] +
//             mat_A[377] * mat_B[802] +
//             mat_A[378] * mat_B[834] +
//             mat_A[379] * mat_B[866] +
//             mat_A[380] * mat_B[898] +
//             mat_A[381] * mat_B[930] +
//             mat_A[382] * mat_B[962] +
//             mat_A[383] * mat_B[994];
//  mat_C[355] <= 
//             mat_A[352] * mat_B[3] +
//             mat_A[353] * mat_B[35] +
//             mat_A[354] * mat_B[67] +
//             mat_A[355] * mat_B[99] +
//             mat_A[356] * mat_B[131] +
//             mat_A[357] * mat_B[163] +
//             mat_A[358] * mat_B[195] +
//             mat_A[359] * mat_B[227] +
//             mat_A[360] * mat_B[259] +
//             mat_A[361] * mat_B[291] +
//             mat_A[362] * mat_B[323] +
//             mat_A[363] * mat_B[355] +
//             mat_A[364] * mat_B[387] +
//             mat_A[365] * mat_B[419] +
//             mat_A[366] * mat_B[451] +
//             mat_A[367] * mat_B[483] +
//             mat_A[368] * mat_B[515] +
//             mat_A[369] * mat_B[547] +
//             mat_A[370] * mat_B[579] +
//             mat_A[371] * mat_B[611] +
//             mat_A[372] * mat_B[643] +
//             mat_A[373] * mat_B[675] +
//             mat_A[374] * mat_B[707] +
//             mat_A[375] * mat_B[739] +
//             mat_A[376] * mat_B[771] +
//             mat_A[377] * mat_B[803] +
//             mat_A[378] * mat_B[835] +
//             mat_A[379] * mat_B[867] +
//             mat_A[380] * mat_B[899] +
//             mat_A[381] * mat_B[931] +
//             mat_A[382] * mat_B[963] +
//             mat_A[383] * mat_B[995];
//  mat_C[356] <= 
//             mat_A[352] * mat_B[4] +
//             mat_A[353] * mat_B[36] +
//             mat_A[354] * mat_B[68] +
//             mat_A[355] * mat_B[100] +
//             mat_A[356] * mat_B[132] +
//             mat_A[357] * mat_B[164] +
//             mat_A[358] * mat_B[196] +
//             mat_A[359] * mat_B[228] +
//             mat_A[360] * mat_B[260] +
//             mat_A[361] * mat_B[292] +
//             mat_A[362] * mat_B[324] +
//             mat_A[363] * mat_B[356] +
//             mat_A[364] * mat_B[388] +
//             mat_A[365] * mat_B[420] +
//             mat_A[366] * mat_B[452] +
//             mat_A[367] * mat_B[484] +
//             mat_A[368] * mat_B[516] +
//             mat_A[369] * mat_B[548] +
//             mat_A[370] * mat_B[580] +
//             mat_A[371] * mat_B[612] +
//             mat_A[372] * mat_B[644] +
//             mat_A[373] * mat_B[676] +
//             mat_A[374] * mat_B[708] +
//             mat_A[375] * mat_B[740] +
//             mat_A[376] * mat_B[772] +
//             mat_A[377] * mat_B[804] +
//             mat_A[378] * mat_B[836] +
//             mat_A[379] * mat_B[868] +
//             mat_A[380] * mat_B[900] +
//             mat_A[381] * mat_B[932] +
//             mat_A[382] * mat_B[964] +
//             mat_A[383] * mat_B[996];
//  mat_C[357] <= 
//             mat_A[352] * mat_B[5] +
//             mat_A[353] * mat_B[37] +
//             mat_A[354] * mat_B[69] +
//             mat_A[355] * mat_B[101] +
//             mat_A[356] * mat_B[133] +
//             mat_A[357] * mat_B[165] +
//             mat_A[358] * mat_B[197] +
//             mat_A[359] * mat_B[229] +
//             mat_A[360] * mat_B[261] +
//             mat_A[361] * mat_B[293] +
//             mat_A[362] * mat_B[325] +
//             mat_A[363] * mat_B[357] +
//             mat_A[364] * mat_B[389] +
//             mat_A[365] * mat_B[421] +
//             mat_A[366] * mat_B[453] +
//             mat_A[367] * mat_B[485] +
//             mat_A[368] * mat_B[517] +
//             mat_A[369] * mat_B[549] +
//             mat_A[370] * mat_B[581] +
//             mat_A[371] * mat_B[613] +
//             mat_A[372] * mat_B[645] +
//             mat_A[373] * mat_B[677] +
//             mat_A[374] * mat_B[709] +
//             mat_A[375] * mat_B[741] +
//             mat_A[376] * mat_B[773] +
//             mat_A[377] * mat_B[805] +
//             mat_A[378] * mat_B[837] +
//             mat_A[379] * mat_B[869] +
//             mat_A[380] * mat_B[901] +
//             mat_A[381] * mat_B[933] +
//             mat_A[382] * mat_B[965] +
//             mat_A[383] * mat_B[997];
//  mat_C[358] <= 
//             mat_A[352] * mat_B[6] +
//             mat_A[353] * mat_B[38] +
//             mat_A[354] * mat_B[70] +
//             mat_A[355] * mat_B[102] +
//             mat_A[356] * mat_B[134] +
//             mat_A[357] * mat_B[166] +
//             mat_A[358] * mat_B[198] +
//             mat_A[359] * mat_B[230] +
//             mat_A[360] * mat_B[262] +
//             mat_A[361] * mat_B[294] +
//             mat_A[362] * mat_B[326] +
//             mat_A[363] * mat_B[358] +
//             mat_A[364] * mat_B[390] +
//             mat_A[365] * mat_B[422] +
//             mat_A[366] * mat_B[454] +
//             mat_A[367] * mat_B[486] +
//             mat_A[368] * mat_B[518] +
//             mat_A[369] * mat_B[550] +
//             mat_A[370] * mat_B[582] +
//             mat_A[371] * mat_B[614] +
//             mat_A[372] * mat_B[646] +
//             mat_A[373] * mat_B[678] +
//             mat_A[374] * mat_B[710] +
//             mat_A[375] * mat_B[742] +
//             mat_A[376] * mat_B[774] +
//             mat_A[377] * mat_B[806] +
//             mat_A[378] * mat_B[838] +
//             mat_A[379] * mat_B[870] +
//             mat_A[380] * mat_B[902] +
//             mat_A[381] * mat_B[934] +
//             mat_A[382] * mat_B[966] +
//             mat_A[383] * mat_B[998];
//  mat_C[359] <= 
//             mat_A[352] * mat_B[7] +
//             mat_A[353] * mat_B[39] +
//             mat_A[354] * mat_B[71] +
//             mat_A[355] * mat_B[103] +
//             mat_A[356] * mat_B[135] +
//             mat_A[357] * mat_B[167] +
//             mat_A[358] * mat_B[199] +
//             mat_A[359] * mat_B[231] +
//             mat_A[360] * mat_B[263] +
//             mat_A[361] * mat_B[295] +
//             mat_A[362] * mat_B[327] +
//             mat_A[363] * mat_B[359] +
//             mat_A[364] * mat_B[391] +
//             mat_A[365] * mat_B[423] +
//             mat_A[366] * mat_B[455] +
//             mat_A[367] * mat_B[487] +
//             mat_A[368] * mat_B[519] +
//             mat_A[369] * mat_B[551] +
//             mat_A[370] * mat_B[583] +
//             mat_A[371] * mat_B[615] +
//             mat_A[372] * mat_B[647] +
//             mat_A[373] * mat_B[679] +
//             mat_A[374] * mat_B[711] +
//             mat_A[375] * mat_B[743] +
//             mat_A[376] * mat_B[775] +
//             mat_A[377] * mat_B[807] +
//             mat_A[378] * mat_B[839] +
//             mat_A[379] * mat_B[871] +
//             mat_A[380] * mat_B[903] +
//             mat_A[381] * mat_B[935] +
//             mat_A[382] * mat_B[967] +
//             mat_A[383] * mat_B[999];
//  mat_C[360] <= 
//             mat_A[352] * mat_B[8] +
//             mat_A[353] * mat_B[40] +
//             mat_A[354] * mat_B[72] +
//             mat_A[355] * mat_B[104] +
//             mat_A[356] * mat_B[136] +
//             mat_A[357] * mat_B[168] +
//             mat_A[358] * mat_B[200] +
//             mat_A[359] * mat_B[232] +
//             mat_A[360] * mat_B[264] +
//             mat_A[361] * mat_B[296] +
//             mat_A[362] * mat_B[328] +
//             mat_A[363] * mat_B[360] +
//             mat_A[364] * mat_B[392] +
//             mat_A[365] * mat_B[424] +
//             mat_A[366] * mat_B[456] +
//             mat_A[367] * mat_B[488] +
//             mat_A[368] * mat_B[520] +
//             mat_A[369] * mat_B[552] +
//             mat_A[370] * mat_B[584] +
//             mat_A[371] * mat_B[616] +
//             mat_A[372] * mat_B[648] +
//             mat_A[373] * mat_B[680] +
//             mat_A[374] * mat_B[712] +
//             mat_A[375] * mat_B[744] +
//             mat_A[376] * mat_B[776] +
//             mat_A[377] * mat_B[808] +
//             mat_A[378] * mat_B[840] +
//             mat_A[379] * mat_B[872] +
//             mat_A[380] * mat_B[904] +
//             mat_A[381] * mat_B[936] +
//             mat_A[382] * mat_B[968] +
//             mat_A[383] * mat_B[1000];
//  mat_C[361] <= 
//             mat_A[352] * mat_B[9] +
//             mat_A[353] * mat_B[41] +
//             mat_A[354] * mat_B[73] +
//             mat_A[355] * mat_B[105] +
//             mat_A[356] * mat_B[137] +
//             mat_A[357] * mat_B[169] +
//             mat_A[358] * mat_B[201] +
//             mat_A[359] * mat_B[233] +
//             mat_A[360] * mat_B[265] +
//             mat_A[361] * mat_B[297] +
//             mat_A[362] * mat_B[329] +
//             mat_A[363] * mat_B[361] +
//             mat_A[364] * mat_B[393] +
//             mat_A[365] * mat_B[425] +
//             mat_A[366] * mat_B[457] +
//             mat_A[367] * mat_B[489] +
//             mat_A[368] * mat_B[521] +
//             mat_A[369] * mat_B[553] +
//             mat_A[370] * mat_B[585] +
//             mat_A[371] * mat_B[617] +
//             mat_A[372] * mat_B[649] +
//             mat_A[373] * mat_B[681] +
//             mat_A[374] * mat_B[713] +
//             mat_A[375] * mat_B[745] +
//             mat_A[376] * mat_B[777] +
//             mat_A[377] * mat_B[809] +
//             mat_A[378] * mat_B[841] +
//             mat_A[379] * mat_B[873] +
//             mat_A[380] * mat_B[905] +
//             mat_A[381] * mat_B[937] +
//             mat_A[382] * mat_B[969] +
//             mat_A[383] * mat_B[1001];
//  mat_C[362] <= 
//             mat_A[352] * mat_B[10] +
//             mat_A[353] * mat_B[42] +
//             mat_A[354] * mat_B[74] +
//             mat_A[355] * mat_B[106] +
//             mat_A[356] * mat_B[138] +
//             mat_A[357] * mat_B[170] +
//             mat_A[358] * mat_B[202] +
//             mat_A[359] * mat_B[234] +
//             mat_A[360] * mat_B[266] +
//             mat_A[361] * mat_B[298] +
//             mat_A[362] * mat_B[330] +
//             mat_A[363] * mat_B[362] +
//             mat_A[364] * mat_B[394] +
//             mat_A[365] * mat_B[426] +
//             mat_A[366] * mat_B[458] +
//             mat_A[367] * mat_B[490] +
//             mat_A[368] * mat_B[522] +
//             mat_A[369] * mat_B[554] +
//             mat_A[370] * mat_B[586] +
//             mat_A[371] * mat_B[618] +
//             mat_A[372] * mat_B[650] +
//             mat_A[373] * mat_B[682] +
//             mat_A[374] * mat_B[714] +
//             mat_A[375] * mat_B[746] +
//             mat_A[376] * mat_B[778] +
//             mat_A[377] * mat_B[810] +
//             mat_A[378] * mat_B[842] +
//             mat_A[379] * mat_B[874] +
//             mat_A[380] * mat_B[906] +
//             mat_A[381] * mat_B[938] +
//             mat_A[382] * mat_B[970] +
//             mat_A[383] * mat_B[1002];
//  mat_C[363] <= 
//             mat_A[352] * mat_B[11] +
//             mat_A[353] * mat_B[43] +
//             mat_A[354] * mat_B[75] +
//             mat_A[355] * mat_B[107] +
//             mat_A[356] * mat_B[139] +
//             mat_A[357] * mat_B[171] +
//             mat_A[358] * mat_B[203] +
//             mat_A[359] * mat_B[235] +
//             mat_A[360] * mat_B[267] +
//             mat_A[361] * mat_B[299] +
//             mat_A[362] * mat_B[331] +
//             mat_A[363] * mat_B[363] +
//             mat_A[364] * mat_B[395] +
//             mat_A[365] * mat_B[427] +
//             mat_A[366] * mat_B[459] +
//             mat_A[367] * mat_B[491] +
//             mat_A[368] * mat_B[523] +
//             mat_A[369] * mat_B[555] +
//             mat_A[370] * mat_B[587] +
//             mat_A[371] * mat_B[619] +
//             mat_A[372] * mat_B[651] +
//             mat_A[373] * mat_B[683] +
//             mat_A[374] * mat_B[715] +
//             mat_A[375] * mat_B[747] +
//             mat_A[376] * mat_B[779] +
//             mat_A[377] * mat_B[811] +
//             mat_A[378] * mat_B[843] +
//             mat_A[379] * mat_B[875] +
//             mat_A[380] * mat_B[907] +
//             mat_A[381] * mat_B[939] +
//             mat_A[382] * mat_B[971] +
//             mat_A[383] * mat_B[1003];
//  mat_C[364] <= 
//             mat_A[352] * mat_B[12] +
//             mat_A[353] * mat_B[44] +
//             mat_A[354] * mat_B[76] +
//             mat_A[355] * mat_B[108] +
//             mat_A[356] * mat_B[140] +
//             mat_A[357] * mat_B[172] +
//             mat_A[358] * mat_B[204] +
//             mat_A[359] * mat_B[236] +
//             mat_A[360] * mat_B[268] +
//             mat_A[361] * mat_B[300] +
//             mat_A[362] * mat_B[332] +
//             mat_A[363] * mat_B[364] +
//             mat_A[364] * mat_B[396] +
//             mat_A[365] * mat_B[428] +
//             mat_A[366] * mat_B[460] +
//             mat_A[367] * mat_B[492] +
//             mat_A[368] * mat_B[524] +
//             mat_A[369] * mat_B[556] +
//             mat_A[370] * mat_B[588] +
//             mat_A[371] * mat_B[620] +
//             mat_A[372] * mat_B[652] +
//             mat_A[373] * mat_B[684] +
//             mat_A[374] * mat_B[716] +
//             mat_A[375] * mat_B[748] +
//             mat_A[376] * mat_B[780] +
//             mat_A[377] * mat_B[812] +
//             mat_A[378] * mat_B[844] +
//             mat_A[379] * mat_B[876] +
//             mat_A[380] * mat_B[908] +
//             mat_A[381] * mat_B[940] +
//             mat_A[382] * mat_B[972] +
//             mat_A[383] * mat_B[1004];
//  mat_C[365] <= 
//             mat_A[352] * mat_B[13] +
//             mat_A[353] * mat_B[45] +
//             mat_A[354] * mat_B[77] +
//             mat_A[355] * mat_B[109] +
//             mat_A[356] * mat_B[141] +
//             mat_A[357] * mat_B[173] +
//             mat_A[358] * mat_B[205] +
//             mat_A[359] * mat_B[237] +
//             mat_A[360] * mat_B[269] +
//             mat_A[361] * mat_B[301] +
//             mat_A[362] * mat_B[333] +
//             mat_A[363] * mat_B[365] +
//             mat_A[364] * mat_B[397] +
//             mat_A[365] * mat_B[429] +
//             mat_A[366] * mat_B[461] +
//             mat_A[367] * mat_B[493] +
//             mat_A[368] * mat_B[525] +
//             mat_A[369] * mat_B[557] +
//             mat_A[370] * mat_B[589] +
//             mat_A[371] * mat_B[621] +
//             mat_A[372] * mat_B[653] +
//             mat_A[373] * mat_B[685] +
//             mat_A[374] * mat_B[717] +
//             mat_A[375] * mat_B[749] +
//             mat_A[376] * mat_B[781] +
//             mat_A[377] * mat_B[813] +
//             mat_A[378] * mat_B[845] +
//             mat_A[379] * mat_B[877] +
//             mat_A[380] * mat_B[909] +
//             mat_A[381] * mat_B[941] +
//             mat_A[382] * mat_B[973] +
//             mat_A[383] * mat_B[1005];
//  mat_C[366] <= 
//             mat_A[352] * mat_B[14] +
//             mat_A[353] * mat_B[46] +
//             mat_A[354] * mat_B[78] +
//             mat_A[355] * mat_B[110] +
//             mat_A[356] * mat_B[142] +
//             mat_A[357] * mat_B[174] +
//             mat_A[358] * mat_B[206] +
//             mat_A[359] * mat_B[238] +
//             mat_A[360] * mat_B[270] +
//             mat_A[361] * mat_B[302] +
//             mat_A[362] * mat_B[334] +
//             mat_A[363] * mat_B[366] +
//             mat_A[364] * mat_B[398] +
//             mat_A[365] * mat_B[430] +
//             mat_A[366] * mat_B[462] +
//             mat_A[367] * mat_B[494] +
//             mat_A[368] * mat_B[526] +
//             mat_A[369] * mat_B[558] +
//             mat_A[370] * mat_B[590] +
//             mat_A[371] * mat_B[622] +
//             mat_A[372] * mat_B[654] +
//             mat_A[373] * mat_B[686] +
//             mat_A[374] * mat_B[718] +
//             mat_A[375] * mat_B[750] +
//             mat_A[376] * mat_B[782] +
//             mat_A[377] * mat_B[814] +
//             mat_A[378] * mat_B[846] +
//             mat_A[379] * mat_B[878] +
//             mat_A[380] * mat_B[910] +
//             mat_A[381] * mat_B[942] +
//             mat_A[382] * mat_B[974] +
//             mat_A[383] * mat_B[1006];
//  mat_C[367] <= 
//             mat_A[352] * mat_B[15] +
//             mat_A[353] * mat_B[47] +
//             mat_A[354] * mat_B[79] +
//             mat_A[355] * mat_B[111] +
//             mat_A[356] * mat_B[143] +
//             mat_A[357] * mat_B[175] +
//             mat_A[358] * mat_B[207] +
//             mat_A[359] * mat_B[239] +
//             mat_A[360] * mat_B[271] +
//             mat_A[361] * mat_B[303] +
//             mat_A[362] * mat_B[335] +
//             mat_A[363] * mat_B[367] +
//             mat_A[364] * mat_B[399] +
//             mat_A[365] * mat_B[431] +
//             mat_A[366] * mat_B[463] +
//             mat_A[367] * mat_B[495] +
//             mat_A[368] * mat_B[527] +
//             mat_A[369] * mat_B[559] +
//             mat_A[370] * mat_B[591] +
//             mat_A[371] * mat_B[623] +
//             mat_A[372] * mat_B[655] +
//             mat_A[373] * mat_B[687] +
//             mat_A[374] * mat_B[719] +
//             mat_A[375] * mat_B[751] +
//             mat_A[376] * mat_B[783] +
//             mat_A[377] * mat_B[815] +
//             mat_A[378] * mat_B[847] +
//             mat_A[379] * mat_B[879] +
//             mat_A[380] * mat_B[911] +
//             mat_A[381] * mat_B[943] +
//             mat_A[382] * mat_B[975] +
//             mat_A[383] * mat_B[1007];
//  mat_C[368] <= 
//             mat_A[352] * mat_B[16] +
//             mat_A[353] * mat_B[48] +
//             mat_A[354] * mat_B[80] +
//             mat_A[355] * mat_B[112] +
//             mat_A[356] * mat_B[144] +
//             mat_A[357] * mat_B[176] +
//             mat_A[358] * mat_B[208] +
//             mat_A[359] * mat_B[240] +
//             mat_A[360] * mat_B[272] +
//             mat_A[361] * mat_B[304] +
//             mat_A[362] * mat_B[336] +
//             mat_A[363] * mat_B[368] +
//             mat_A[364] * mat_B[400] +
//             mat_A[365] * mat_B[432] +
//             mat_A[366] * mat_B[464] +
//             mat_A[367] * mat_B[496] +
//             mat_A[368] * mat_B[528] +
//             mat_A[369] * mat_B[560] +
//             mat_A[370] * mat_B[592] +
//             mat_A[371] * mat_B[624] +
//             mat_A[372] * mat_B[656] +
//             mat_A[373] * mat_B[688] +
//             mat_A[374] * mat_B[720] +
//             mat_A[375] * mat_B[752] +
//             mat_A[376] * mat_B[784] +
//             mat_A[377] * mat_B[816] +
//             mat_A[378] * mat_B[848] +
//             mat_A[379] * mat_B[880] +
//             mat_A[380] * mat_B[912] +
//             mat_A[381] * mat_B[944] +
//             mat_A[382] * mat_B[976] +
//             mat_A[383] * mat_B[1008];
//  mat_C[369] <= 
//             mat_A[352] * mat_B[17] +
//             mat_A[353] * mat_B[49] +
//             mat_A[354] * mat_B[81] +
//             mat_A[355] * mat_B[113] +
//             mat_A[356] * mat_B[145] +
//             mat_A[357] * mat_B[177] +
//             mat_A[358] * mat_B[209] +
//             mat_A[359] * mat_B[241] +
//             mat_A[360] * mat_B[273] +
//             mat_A[361] * mat_B[305] +
//             mat_A[362] * mat_B[337] +
//             mat_A[363] * mat_B[369] +
//             mat_A[364] * mat_B[401] +
//             mat_A[365] * mat_B[433] +
//             mat_A[366] * mat_B[465] +
//             mat_A[367] * mat_B[497] +
//             mat_A[368] * mat_B[529] +
//             mat_A[369] * mat_B[561] +
//             mat_A[370] * mat_B[593] +
//             mat_A[371] * mat_B[625] +
//             mat_A[372] * mat_B[657] +
//             mat_A[373] * mat_B[689] +
//             mat_A[374] * mat_B[721] +
//             mat_A[375] * mat_B[753] +
//             mat_A[376] * mat_B[785] +
//             mat_A[377] * mat_B[817] +
//             mat_A[378] * mat_B[849] +
//             mat_A[379] * mat_B[881] +
//             mat_A[380] * mat_B[913] +
//             mat_A[381] * mat_B[945] +
//             mat_A[382] * mat_B[977] +
//             mat_A[383] * mat_B[1009];
//  mat_C[370] <= 
//             mat_A[352] * mat_B[18] +
//             mat_A[353] * mat_B[50] +
//             mat_A[354] * mat_B[82] +
//             mat_A[355] * mat_B[114] +
//             mat_A[356] * mat_B[146] +
//             mat_A[357] * mat_B[178] +
//             mat_A[358] * mat_B[210] +
//             mat_A[359] * mat_B[242] +
//             mat_A[360] * mat_B[274] +
//             mat_A[361] * mat_B[306] +
//             mat_A[362] * mat_B[338] +
//             mat_A[363] * mat_B[370] +
//             mat_A[364] * mat_B[402] +
//             mat_A[365] * mat_B[434] +
//             mat_A[366] * mat_B[466] +
//             mat_A[367] * mat_B[498] +
//             mat_A[368] * mat_B[530] +
//             mat_A[369] * mat_B[562] +
//             mat_A[370] * mat_B[594] +
//             mat_A[371] * mat_B[626] +
//             mat_A[372] * mat_B[658] +
//             mat_A[373] * mat_B[690] +
//             mat_A[374] * mat_B[722] +
//             mat_A[375] * mat_B[754] +
//             mat_A[376] * mat_B[786] +
//             mat_A[377] * mat_B[818] +
//             mat_A[378] * mat_B[850] +
//             mat_A[379] * mat_B[882] +
//             mat_A[380] * mat_B[914] +
//             mat_A[381] * mat_B[946] +
//             mat_A[382] * mat_B[978] +
//             mat_A[383] * mat_B[1010];
//  mat_C[371] <= 
//             mat_A[352] * mat_B[19] +
//             mat_A[353] * mat_B[51] +
//             mat_A[354] * mat_B[83] +
//             mat_A[355] * mat_B[115] +
//             mat_A[356] * mat_B[147] +
//             mat_A[357] * mat_B[179] +
//             mat_A[358] * mat_B[211] +
//             mat_A[359] * mat_B[243] +
//             mat_A[360] * mat_B[275] +
//             mat_A[361] * mat_B[307] +
//             mat_A[362] * mat_B[339] +
//             mat_A[363] * mat_B[371] +
//             mat_A[364] * mat_B[403] +
//             mat_A[365] * mat_B[435] +
//             mat_A[366] * mat_B[467] +
//             mat_A[367] * mat_B[499] +
//             mat_A[368] * mat_B[531] +
//             mat_A[369] * mat_B[563] +
//             mat_A[370] * mat_B[595] +
//             mat_A[371] * mat_B[627] +
//             mat_A[372] * mat_B[659] +
//             mat_A[373] * mat_B[691] +
//             mat_A[374] * mat_B[723] +
//             mat_A[375] * mat_B[755] +
//             mat_A[376] * mat_B[787] +
//             mat_A[377] * mat_B[819] +
//             mat_A[378] * mat_B[851] +
//             mat_A[379] * mat_B[883] +
//             mat_A[380] * mat_B[915] +
//             mat_A[381] * mat_B[947] +
//             mat_A[382] * mat_B[979] +
//             mat_A[383] * mat_B[1011];
//  mat_C[372] <= 
//             mat_A[352] * mat_B[20] +
//             mat_A[353] * mat_B[52] +
//             mat_A[354] * mat_B[84] +
//             mat_A[355] * mat_B[116] +
//             mat_A[356] * mat_B[148] +
//             mat_A[357] * mat_B[180] +
//             mat_A[358] * mat_B[212] +
//             mat_A[359] * mat_B[244] +
//             mat_A[360] * mat_B[276] +
//             mat_A[361] * mat_B[308] +
//             mat_A[362] * mat_B[340] +
//             mat_A[363] * mat_B[372] +
//             mat_A[364] * mat_B[404] +
//             mat_A[365] * mat_B[436] +
//             mat_A[366] * mat_B[468] +
//             mat_A[367] * mat_B[500] +
//             mat_A[368] * mat_B[532] +
//             mat_A[369] * mat_B[564] +
//             mat_A[370] * mat_B[596] +
//             mat_A[371] * mat_B[628] +
//             mat_A[372] * mat_B[660] +
//             mat_A[373] * mat_B[692] +
//             mat_A[374] * mat_B[724] +
//             mat_A[375] * mat_B[756] +
//             mat_A[376] * mat_B[788] +
//             mat_A[377] * mat_B[820] +
//             mat_A[378] * mat_B[852] +
//             mat_A[379] * mat_B[884] +
//             mat_A[380] * mat_B[916] +
//             mat_A[381] * mat_B[948] +
//             mat_A[382] * mat_B[980] +
//             mat_A[383] * mat_B[1012];
//  mat_C[373] <= 
//             mat_A[352] * mat_B[21] +
//             mat_A[353] * mat_B[53] +
//             mat_A[354] * mat_B[85] +
//             mat_A[355] * mat_B[117] +
//             mat_A[356] * mat_B[149] +
//             mat_A[357] * mat_B[181] +
//             mat_A[358] * mat_B[213] +
//             mat_A[359] * mat_B[245] +
//             mat_A[360] * mat_B[277] +
//             mat_A[361] * mat_B[309] +
//             mat_A[362] * mat_B[341] +
//             mat_A[363] * mat_B[373] +
//             mat_A[364] * mat_B[405] +
//             mat_A[365] * mat_B[437] +
//             mat_A[366] * mat_B[469] +
//             mat_A[367] * mat_B[501] +
//             mat_A[368] * mat_B[533] +
//             mat_A[369] * mat_B[565] +
//             mat_A[370] * mat_B[597] +
//             mat_A[371] * mat_B[629] +
//             mat_A[372] * mat_B[661] +
//             mat_A[373] * mat_B[693] +
//             mat_A[374] * mat_B[725] +
//             mat_A[375] * mat_B[757] +
//             mat_A[376] * mat_B[789] +
//             mat_A[377] * mat_B[821] +
//             mat_A[378] * mat_B[853] +
//             mat_A[379] * mat_B[885] +
//             mat_A[380] * mat_B[917] +
//             mat_A[381] * mat_B[949] +
//             mat_A[382] * mat_B[981] +
//             mat_A[383] * mat_B[1013];
//  mat_C[374] <= 
//             mat_A[352] * mat_B[22] +
//             mat_A[353] * mat_B[54] +
//             mat_A[354] * mat_B[86] +
//             mat_A[355] * mat_B[118] +
//             mat_A[356] * mat_B[150] +
//             mat_A[357] * mat_B[182] +
//             mat_A[358] * mat_B[214] +
//             mat_A[359] * mat_B[246] +
//             mat_A[360] * mat_B[278] +
//             mat_A[361] * mat_B[310] +
//             mat_A[362] * mat_B[342] +
//             mat_A[363] * mat_B[374] +
//             mat_A[364] * mat_B[406] +
//             mat_A[365] * mat_B[438] +
//             mat_A[366] * mat_B[470] +
//             mat_A[367] * mat_B[502] +
//             mat_A[368] * mat_B[534] +
//             mat_A[369] * mat_B[566] +
//             mat_A[370] * mat_B[598] +
//             mat_A[371] * mat_B[630] +
//             mat_A[372] * mat_B[662] +
//             mat_A[373] * mat_B[694] +
//             mat_A[374] * mat_B[726] +
//             mat_A[375] * mat_B[758] +
//             mat_A[376] * mat_B[790] +
//             mat_A[377] * mat_B[822] +
//             mat_A[378] * mat_B[854] +
//             mat_A[379] * mat_B[886] +
//             mat_A[380] * mat_B[918] +
//             mat_A[381] * mat_B[950] +
//             mat_A[382] * mat_B[982] +
//             mat_A[383] * mat_B[1014];
//  mat_C[375] <= 
//             mat_A[352] * mat_B[23] +
//             mat_A[353] * mat_B[55] +
//             mat_A[354] * mat_B[87] +
//             mat_A[355] * mat_B[119] +
//             mat_A[356] * mat_B[151] +
//             mat_A[357] * mat_B[183] +
//             mat_A[358] * mat_B[215] +
//             mat_A[359] * mat_B[247] +
//             mat_A[360] * mat_B[279] +
//             mat_A[361] * mat_B[311] +
//             mat_A[362] * mat_B[343] +
//             mat_A[363] * mat_B[375] +
//             mat_A[364] * mat_B[407] +
//             mat_A[365] * mat_B[439] +
//             mat_A[366] * mat_B[471] +
//             mat_A[367] * mat_B[503] +
//             mat_A[368] * mat_B[535] +
//             mat_A[369] * mat_B[567] +
//             mat_A[370] * mat_B[599] +
//             mat_A[371] * mat_B[631] +
//             mat_A[372] * mat_B[663] +
//             mat_A[373] * mat_B[695] +
//             mat_A[374] * mat_B[727] +
//             mat_A[375] * mat_B[759] +
//             mat_A[376] * mat_B[791] +
//             mat_A[377] * mat_B[823] +
//             mat_A[378] * mat_B[855] +
//             mat_A[379] * mat_B[887] +
//             mat_A[380] * mat_B[919] +
//             mat_A[381] * mat_B[951] +
//             mat_A[382] * mat_B[983] +
//             mat_A[383] * mat_B[1015];
//  mat_C[376] <= 
//             mat_A[352] * mat_B[24] +
//             mat_A[353] * mat_B[56] +
//             mat_A[354] * mat_B[88] +
//             mat_A[355] * mat_B[120] +
//             mat_A[356] * mat_B[152] +
//             mat_A[357] * mat_B[184] +
//             mat_A[358] * mat_B[216] +
//             mat_A[359] * mat_B[248] +
//             mat_A[360] * mat_B[280] +
//             mat_A[361] * mat_B[312] +
//             mat_A[362] * mat_B[344] +
//             mat_A[363] * mat_B[376] +
//             mat_A[364] * mat_B[408] +
//             mat_A[365] * mat_B[440] +
//             mat_A[366] * mat_B[472] +
//             mat_A[367] * mat_B[504] +
//             mat_A[368] * mat_B[536] +
//             mat_A[369] * mat_B[568] +
//             mat_A[370] * mat_B[600] +
//             mat_A[371] * mat_B[632] +
//             mat_A[372] * mat_B[664] +
//             mat_A[373] * mat_B[696] +
//             mat_A[374] * mat_B[728] +
//             mat_A[375] * mat_B[760] +
//             mat_A[376] * mat_B[792] +
//             mat_A[377] * mat_B[824] +
//             mat_A[378] * mat_B[856] +
//             mat_A[379] * mat_B[888] +
//             mat_A[380] * mat_B[920] +
//             mat_A[381] * mat_B[952] +
//             mat_A[382] * mat_B[984] +
//             mat_A[383] * mat_B[1016];
//  mat_C[377] <= 
//             mat_A[352] * mat_B[25] +
//             mat_A[353] * mat_B[57] +
//             mat_A[354] * mat_B[89] +
//             mat_A[355] * mat_B[121] +
//             mat_A[356] * mat_B[153] +
//             mat_A[357] * mat_B[185] +
//             mat_A[358] * mat_B[217] +
//             mat_A[359] * mat_B[249] +
//             mat_A[360] * mat_B[281] +
//             mat_A[361] * mat_B[313] +
//             mat_A[362] * mat_B[345] +
//             mat_A[363] * mat_B[377] +
//             mat_A[364] * mat_B[409] +
//             mat_A[365] * mat_B[441] +
//             mat_A[366] * mat_B[473] +
//             mat_A[367] * mat_B[505] +
//             mat_A[368] * mat_B[537] +
//             mat_A[369] * mat_B[569] +
//             mat_A[370] * mat_B[601] +
//             mat_A[371] * mat_B[633] +
//             mat_A[372] * mat_B[665] +
//             mat_A[373] * mat_B[697] +
//             mat_A[374] * mat_B[729] +
//             mat_A[375] * mat_B[761] +
//             mat_A[376] * mat_B[793] +
//             mat_A[377] * mat_B[825] +
//             mat_A[378] * mat_B[857] +
//             mat_A[379] * mat_B[889] +
//             mat_A[380] * mat_B[921] +
//             mat_A[381] * mat_B[953] +
//             mat_A[382] * mat_B[985] +
//             mat_A[383] * mat_B[1017];
//  mat_C[378] <= 
//             mat_A[352] * mat_B[26] +
//             mat_A[353] * mat_B[58] +
//             mat_A[354] * mat_B[90] +
//             mat_A[355] * mat_B[122] +
//             mat_A[356] * mat_B[154] +
//             mat_A[357] * mat_B[186] +
//             mat_A[358] * mat_B[218] +
//             mat_A[359] * mat_B[250] +
//             mat_A[360] * mat_B[282] +
//             mat_A[361] * mat_B[314] +
//             mat_A[362] * mat_B[346] +
//             mat_A[363] * mat_B[378] +
//             mat_A[364] * mat_B[410] +
//             mat_A[365] * mat_B[442] +
//             mat_A[366] * mat_B[474] +
//             mat_A[367] * mat_B[506] +
//             mat_A[368] * mat_B[538] +
//             mat_A[369] * mat_B[570] +
//             mat_A[370] * mat_B[602] +
//             mat_A[371] * mat_B[634] +
//             mat_A[372] * mat_B[666] +
//             mat_A[373] * mat_B[698] +
//             mat_A[374] * mat_B[730] +
//             mat_A[375] * mat_B[762] +
//             mat_A[376] * mat_B[794] +
//             mat_A[377] * mat_B[826] +
//             mat_A[378] * mat_B[858] +
//             mat_A[379] * mat_B[890] +
//             mat_A[380] * mat_B[922] +
//             mat_A[381] * mat_B[954] +
//             mat_A[382] * mat_B[986] +
//             mat_A[383] * mat_B[1018];
//  mat_C[379] <= 
//             mat_A[352] * mat_B[27] +
//             mat_A[353] * mat_B[59] +
//             mat_A[354] * mat_B[91] +
//             mat_A[355] * mat_B[123] +
//             mat_A[356] * mat_B[155] +
//             mat_A[357] * mat_B[187] +
//             mat_A[358] * mat_B[219] +
//             mat_A[359] * mat_B[251] +
//             mat_A[360] * mat_B[283] +
//             mat_A[361] * mat_B[315] +
//             mat_A[362] * mat_B[347] +
//             mat_A[363] * mat_B[379] +
//             mat_A[364] * mat_B[411] +
//             mat_A[365] * mat_B[443] +
//             mat_A[366] * mat_B[475] +
//             mat_A[367] * mat_B[507] +
//             mat_A[368] * mat_B[539] +
//             mat_A[369] * mat_B[571] +
//             mat_A[370] * mat_B[603] +
//             mat_A[371] * mat_B[635] +
//             mat_A[372] * mat_B[667] +
//             mat_A[373] * mat_B[699] +
//             mat_A[374] * mat_B[731] +
//             mat_A[375] * mat_B[763] +
//             mat_A[376] * mat_B[795] +
//             mat_A[377] * mat_B[827] +
//             mat_A[378] * mat_B[859] +
//             mat_A[379] * mat_B[891] +
//             mat_A[380] * mat_B[923] +
//             mat_A[381] * mat_B[955] +
//             mat_A[382] * mat_B[987] +
//             mat_A[383] * mat_B[1019];
//  mat_C[380] <= 
//             mat_A[352] * mat_B[28] +
//             mat_A[353] * mat_B[60] +
//             mat_A[354] * mat_B[92] +
//             mat_A[355] * mat_B[124] +
//             mat_A[356] * mat_B[156] +
//             mat_A[357] * mat_B[188] +
//             mat_A[358] * mat_B[220] +
//             mat_A[359] * mat_B[252] +
//             mat_A[360] * mat_B[284] +
//             mat_A[361] * mat_B[316] +
//             mat_A[362] * mat_B[348] +
//             mat_A[363] * mat_B[380] +
//             mat_A[364] * mat_B[412] +
//             mat_A[365] * mat_B[444] +
//             mat_A[366] * mat_B[476] +
//             mat_A[367] * mat_B[508] +
//             mat_A[368] * mat_B[540] +
//             mat_A[369] * mat_B[572] +
//             mat_A[370] * mat_B[604] +
//             mat_A[371] * mat_B[636] +
//             mat_A[372] * mat_B[668] +
//             mat_A[373] * mat_B[700] +
//             mat_A[374] * mat_B[732] +
//             mat_A[375] * mat_B[764] +
//             mat_A[376] * mat_B[796] +
//             mat_A[377] * mat_B[828] +
//             mat_A[378] * mat_B[860] +
//             mat_A[379] * mat_B[892] +
//             mat_A[380] * mat_B[924] +
//             mat_A[381] * mat_B[956] +
//             mat_A[382] * mat_B[988] +
//             mat_A[383] * mat_B[1020];
//  mat_C[381] <= 
//             mat_A[352] * mat_B[29] +
//             mat_A[353] * mat_B[61] +
//             mat_A[354] * mat_B[93] +
//             mat_A[355] * mat_B[125] +
//             mat_A[356] * mat_B[157] +
//             mat_A[357] * mat_B[189] +
//             mat_A[358] * mat_B[221] +
//             mat_A[359] * mat_B[253] +
//             mat_A[360] * mat_B[285] +
//             mat_A[361] * mat_B[317] +
//             mat_A[362] * mat_B[349] +
//             mat_A[363] * mat_B[381] +
//             mat_A[364] * mat_B[413] +
//             mat_A[365] * mat_B[445] +
//             mat_A[366] * mat_B[477] +
//             mat_A[367] * mat_B[509] +
//             mat_A[368] * mat_B[541] +
//             mat_A[369] * mat_B[573] +
//             mat_A[370] * mat_B[605] +
//             mat_A[371] * mat_B[637] +
//             mat_A[372] * mat_B[669] +
//             mat_A[373] * mat_B[701] +
//             mat_A[374] * mat_B[733] +
//             mat_A[375] * mat_B[765] +
//             mat_A[376] * mat_B[797] +
//             mat_A[377] * mat_B[829] +
//             mat_A[378] * mat_B[861] +
//             mat_A[379] * mat_B[893] +
//             mat_A[380] * mat_B[925] +
//             mat_A[381] * mat_B[957] +
//             mat_A[382] * mat_B[989] +
//             mat_A[383] * mat_B[1021];
//  mat_C[382] <= 
//             mat_A[352] * mat_B[30] +
//             mat_A[353] * mat_B[62] +
//             mat_A[354] * mat_B[94] +
//             mat_A[355] * mat_B[126] +
//             mat_A[356] * mat_B[158] +
//             mat_A[357] * mat_B[190] +
//             mat_A[358] * mat_B[222] +
//             mat_A[359] * mat_B[254] +
//             mat_A[360] * mat_B[286] +
//             mat_A[361] * mat_B[318] +
//             mat_A[362] * mat_B[350] +
//             mat_A[363] * mat_B[382] +
//             mat_A[364] * mat_B[414] +
//             mat_A[365] * mat_B[446] +
//             mat_A[366] * mat_B[478] +
//             mat_A[367] * mat_B[510] +
//             mat_A[368] * mat_B[542] +
//             mat_A[369] * mat_B[574] +
//             mat_A[370] * mat_B[606] +
//             mat_A[371] * mat_B[638] +
//             mat_A[372] * mat_B[670] +
//             mat_A[373] * mat_B[702] +
//             mat_A[374] * mat_B[734] +
//             mat_A[375] * mat_B[766] +
//             mat_A[376] * mat_B[798] +
//             mat_A[377] * mat_B[830] +
//             mat_A[378] * mat_B[862] +
//             mat_A[379] * mat_B[894] +
//             mat_A[380] * mat_B[926] +
//             mat_A[381] * mat_B[958] +
//             mat_A[382] * mat_B[990] +
//             mat_A[383] * mat_B[1022];
//  mat_C[383] <= 
//             mat_A[352] * mat_B[31] +
//             mat_A[353] * mat_B[63] +
//             mat_A[354] * mat_B[95] +
//             mat_A[355] * mat_B[127] +
//             mat_A[356] * mat_B[159] +
//             mat_A[357] * mat_B[191] +
//             mat_A[358] * mat_B[223] +
//             mat_A[359] * mat_B[255] +
//             mat_A[360] * mat_B[287] +
//             mat_A[361] * mat_B[319] +
//             mat_A[362] * mat_B[351] +
//             mat_A[363] * mat_B[383] +
//             mat_A[364] * mat_B[415] +
//             mat_A[365] * mat_B[447] +
//             mat_A[366] * mat_B[479] +
//             mat_A[367] * mat_B[511] +
//             mat_A[368] * mat_B[543] +
//             mat_A[369] * mat_B[575] +
//             mat_A[370] * mat_B[607] +
//             mat_A[371] * mat_B[639] +
//             mat_A[372] * mat_B[671] +
//             mat_A[373] * mat_B[703] +
//             mat_A[374] * mat_B[735] +
//             mat_A[375] * mat_B[767] +
//             mat_A[376] * mat_B[799] +
//             mat_A[377] * mat_B[831] +
//             mat_A[378] * mat_B[863] +
//             mat_A[379] * mat_B[895] +
//             mat_A[380] * mat_B[927] +
//             mat_A[381] * mat_B[959] +
//             mat_A[382] * mat_B[991] +
//             mat_A[383] * mat_B[1023];
//  mat_C[384] <= 
//             mat_A[384] * mat_B[0] +
//             mat_A[385] * mat_B[32] +
//             mat_A[386] * mat_B[64] +
//             mat_A[387] * mat_B[96] +
//             mat_A[388] * mat_B[128] +
//             mat_A[389] * mat_B[160] +
//             mat_A[390] * mat_B[192] +
//             mat_A[391] * mat_B[224] +
//             mat_A[392] * mat_B[256] +
//             mat_A[393] * mat_B[288] +
//             mat_A[394] * mat_B[320] +
//             mat_A[395] * mat_B[352] +
//             mat_A[396] * mat_B[384] +
//             mat_A[397] * mat_B[416] +
//             mat_A[398] * mat_B[448] +
//             mat_A[399] * mat_B[480] +
//             mat_A[400] * mat_B[512] +
//             mat_A[401] * mat_B[544] +
//             mat_A[402] * mat_B[576] +
//             mat_A[403] * mat_B[608] +
//             mat_A[404] * mat_B[640] +
//             mat_A[405] * mat_B[672] +
//             mat_A[406] * mat_B[704] +
//             mat_A[407] * mat_B[736] +
//             mat_A[408] * mat_B[768] +
//             mat_A[409] * mat_B[800] +
//             mat_A[410] * mat_B[832] +
//             mat_A[411] * mat_B[864] +
//             mat_A[412] * mat_B[896] +
//             mat_A[413] * mat_B[928] +
//             mat_A[414] * mat_B[960] +
//             mat_A[415] * mat_B[992];
//  mat_C[385] <= 
//             mat_A[384] * mat_B[1] +
//             mat_A[385] * mat_B[33] +
//             mat_A[386] * mat_B[65] +
//             mat_A[387] * mat_B[97] +
//             mat_A[388] * mat_B[129] +
//             mat_A[389] * mat_B[161] +
//             mat_A[390] * mat_B[193] +
//             mat_A[391] * mat_B[225] +
//             mat_A[392] * mat_B[257] +
//             mat_A[393] * mat_B[289] +
//             mat_A[394] * mat_B[321] +
//             mat_A[395] * mat_B[353] +
//             mat_A[396] * mat_B[385] +
//             mat_A[397] * mat_B[417] +
//             mat_A[398] * mat_B[449] +
//             mat_A[399] * mat_B[481] +
//             mat_A[400] * mat_B[513] +
//             mat_A[401] * mat_B[545] +
//             mat_A[402] * mat_B[577] +
//             mat_A[403] * mat_B[609] +
//             mat_A[404] * mat_B[641] +
//             mat_A[405] * mat_B[673] +
//             mat_A[406] * mat_B[705] +
//             mat_A[407] * mat_B[737] +
//             mat_A[408] * mat_B[769] +
//             mat_A[409] * mat_B[801] +
//             mat_A[410] * mat_B[833] +
//             mat_A[411] * mat_B[865] +
//             mat_A[412] * mat_B[897] +
//             mat_A[413] * mat_B[929] +
//             mat_A[414] * mat_B[961] +
//             mat_A[415] * mat_B[993];
//  mat_C[386] <= 
//             mat_A[384] * mat_B[2] +
//             mat_A[385] * mat_B[34] +
//             mat_A[386] * mat_B[66] +
//             mat_A[387] * mat_B[98] +
//             mat_A[388] * mat_B[130] +
//             mat_A[389] * mat_B[162] +
//             mat_A[390] * mat_B[194] +
//             mat_A[391] * mat_B[226] +
//             mat_A[392] * mat_B[258] +
//             mat_A[393] * mat_B[290] +
//             mat_A[394] * mat_B[322] +
//             mat_A[395] * mat_B[354] +
//             mat_A[396] * mat_B[386] +
//             mat_A[397] * mat_B[418] +
//             mat_A[398] * mat_B[450] +
//             mat_A[399] * mat_B[482] +
//             mat_A[400] * mat_B[514] +
//             mat_A[401] * mat_B[546] +
//             mat_A[402] * mat_B[578] +
//             mat_A[403] * mat_B[610] +
//             mat_A[404] * mat_B[642] +
//             mat_A[405] * mat_B[674] +
//             mat_A[406] * mat_B[706] +
//             mat_A[407] * mat_B[738] +
//             mat_A[408] * mat_B[770] +
//             mat_A[409] * mat_B[802] +
//             mat_A[410] * mat_B[834] +
//             mat_A[411] * mat_B[866] +
//             mat_A[412] * mat_B[898] +
//             mat_A[413] * mat_B[930] +
//             mat_A[414] * mat_B[962] +
//             mat_A[415] * mat_B[994];
//  mat_C[387] <= 
//             mat_A[384] * mat_B[3] +
//             mat_A[385] * mat_B[35] +
//             mat_A[386] * mat_B[67] +
//             mat_A[387] * mat_B[99] +
//             mat_A[388] * mat_B[131] +
//             mat_A[389] * mat_B[163] +
//             mat_A[390] * mat_B[195] +
//             mat_A[391] * mat_B[227] +
//             mat_A[392] * mat_B[259] +
//             mat_A[393] * mat_B[291] +
//             mat_A[394] * mat_B[323] +
//             mat_A[395] * mat_B[355] +
//             mat_A[396] * mat_B[387] +
//             mat_A[397] * mat_B[419] +
//             mat_A[398] * mat_B[451] +
//             mat_A[399] * mat_B[483] +
//             mat_A[400] * mat_B[515] +
//             mat_A[401] * mat_B[547] +
//             mat_A[402] * mat_B[579] +
//             mat_A[403] * mat_B[611] +
//             mat_A[404] * mat_B[643] +
//             mat_A[405] * mat_B[675] +
//             mat_A[406] * mat_B[707] +
//             mat_A[407] * mat_B[739] +
//             mat_A[408] * mat_B[771] +
//             mat_A[409] * mat_B[803] +
//             mat_A[410] * mat_B[835] +
//             mat_A[411] * mat_B[867] +
//             mat_A[412] * mat_B[899] +
//             mat_A[413] * mat_B[931] +
//             mat_A[414] * mat_B[963] +
//             mat_A[415] * mat_B[995];
//  mat_C[388] <= 
//             mat_A[384] * mat_B[4] +
//             mat_A[385] * mat_B[36] +
//             mat_A[386] * mat_B[68] +
//             mat_A[387] * mat_B[100] +
//             mat_A[388] * mat_B[132] +
//             mat_A[389] * mat_B[164] +
//             mat_A[390] * mat_B[196] +
//             mat_A[391] * mat_B[228] +
//             mat_A[392] * mat_B[260] +
//             mat_A[393] * mat_B[292] +
//             mat_A[394] * mat_B[324] +
//             mat_A[395] * mat_B[356] +
//             mat_A[396] * mat_B[388] +
//             mat_A[397] * mat_B[420] +
//             mat_A[398] * mat_B[452] +
//             mat_A[399] * mat_B[484] +
//             mat_A[400] * mat_B[516] +
//             mat_A[401] * mat_B[548] +
//             mat_A[402] * mat_B[580] +
//             mat_A[403] * mat_B[612] +
//             mat_A[404] * mat_B[644] +
//             mat_A[405] * mat_B[676] +
//             mat_A[406] * mat_B[708] +
//             mat_A[407] * mat_B[740] +
//             mat_A[408] * mat_B[772] +
//             mat_A[409] * mat_B[804] +
//             mat_A[410] * mat_B[836] +
//             mat_A[411] * mat_B[868] +
//             mat_A[412] * mat_B[900] +
//             mat_A[413] * mat_B[932] +
//             mat_A[414] * mat_B[964] +
//             mat_A[415] * mat_B[996];
//  mat_C[389] <= 
//             mat_A[384] * mat_B[5] +
//             mat_A[385] * mat_B[37] +
//             mat_A[386] * mat_B[69] +
//             mat_A[387] * mat_B[101] +
//             mat_A[388] * mat_B[133] +
//             mat_A[389] * mat_B[165] +
//             mat_A[390] * mat_B[197] +
//             mat_A[391] * mat_B[229] +
//             mat_A[392] * mat_B[261] +
//             mat_A[393] * mat_B[293] +
//             mat_A[394] * mat_B[325] +
//             mat_A[395] * mat_B[357] +
//             mat_A[396] * mat_B[389] +
//             mat_A[397] * mat_B[421] +
//             mat_A[398] * mat_B[453] +
//             mat_A[399] * mat_B[485] +
//             mat_A[400] * mat_B[517] +
//             mat_A[401] * mat_B[549] +
//             mat_A[402] * mat_B[581] +
//             mat_A[403] * mat_B[613] +
//             mat_A[404] * mat_B[645] +
//             mat_A[405] * mat_B[677] +
//             mat_A[406] * mat_B[709] +
//             mat_A[407] * mat_B[741] +
//             mat_A[408] * mat_B[773] +
//             mat_A[409] * mat_B[805] +
//             mat_A[410] * mat_B[837] +
//             mat_A[411] * mat_B[869] +
//             mat_A[412] * mat_B[901] +
//             mat_A[413] * mat_B[933] +
//             mat_A[414] * mat_B[965] +
//             mat_A[415] * mat_B[997];
//  mat_C[390] <= 
//             mat_A[384] * mat_B[6] +
//             mat_A[385] * mat_B[38] +
//             mat_A[386] * mat_B[70] +
//             mat_A[387] * mat_B[102] +
//             mat_A[388] * mat_B[134] +
//             mat_A[389] * mat_B[166] +
//             mat_A[390] * mat_B[198] +
//             mat_A[391] * mat_B[230] +
//             mat_A[392] * mat_B[262] +
//             mat_A[393] * mat_B[294] +
//             mat_A[394] * mat_B[326] +
//             mat_A[395] * mat_B[358] +
//             mat_A[396] * mat_B[390] +
//             mat_A[397] * mat_B[422] +
//             mat_A[398] * mat_B[454] +
//             mat_A[399] * mat_B[486] +
//             mat_A[400] * mat_B[518] +
//             mat_A[401] * mat_B[550] +
//             mat_A[402] * mat_B[582] +
//             mat_A[403] * mat_B[614] +
//             mat_A[404] * mat_B[646] +
//             mat_A[405] * mat_B[678] +
//             mat_A[406] * mat_B[710] +
//             mat_A[407] * mat_B[742] +
//             mat_A[408] * mat_B[774] +
//             mat_A[409] * mat_B[806] +
//             mat_A[410] * mat_B[838] +
//             mat_A[411] * mat_B[870] +
//             mat_A[412] * mat_B[902] +
//             mat_A[413] * mat_B[934] +
//             mat_A[414] * mat_B[966] +
//             mat_A[415] * mat_B[998];
//  mat_C[391] <= 
//             mat_A[384] * mat_B[7] +
//             mat_A[385] * mat_B[39] +
//             mat_A[386] * mat_B[71] +
//             mat_A[387] * mat_B[103] +
//             mat_A[388] * mat_B[135] +
//             mat_A[389] * mat_B[167] +
//             mat_A[390] * mat_B[199] +
//             mat_A[391] * mat_B[231] +
//             mat_A[392] * mat_B[263] +
//             mat_A[393] * mat_B[295] +
//             mat_A[394] * mat_B[327] +
//             mat_A[395] * mat_B[359] +
//             mat_A[396] * mat_B[391] +
//             mat_A[397] * mat_B[423] +
//             mat_A[398] * mat_B[455] +
//             mat_A[399] * mat_B[487] +
//             mat_A[400] * mat_B[519] +
//             mat_A[401] * mat_B[551] +
//             mat_A[402] * mat_B[583] +
//             mat_A[403] * mat_B[615] +
//             mat_A[404] * mat_B[647] +
//             mat_A[405] * mat_B[679] +
//             mat_A[406] * mat_B[711] +
//             mat_A[407] * mat_B[743] +
//             mat_A[408] * mat_B[775] +
//             mat_A[409] * mat_B[807] +
//             mat_A[410] * mat_B[839] +
//             mat_A[411] * mat_B[871] +
//             mat_A[412] * mat_B[903] +
//             mat_A[413] * mat_B[935] +
//             mat_A[414] * mat_B[967] +
//             mat_A[415] * mat_B[999];
//  mat_C[392] <= 
//             mat_A[384] * mat_B[8] +
//             mat_A[385] * mat_B[40] +
//             mat_A[386] * mat_B[72] +
//             mat_A[387] * mat_B[104] +
//             mat_A[388] * mat_B[136] +
//             mat_A[389] * mat_B[168] +
//             mat_A[390] * mat_B[200] +
//             mat_A[391] * mat_B[232] +
//             mat_A[392] * mat_B[264] +
//             mat_A[393] * mat_B[296] +
//             mat_A[394] * mat_B[328] +
//             mat_A[395] * mat_B[360] +
//             mat_A[396] * mat_B[392] +
//             mat_A[397] * mat_B[424] +
//             mat_A[398] * mat_B[456] +
//             mat_A[399] * mat_B[488] +
//             mat_A[400] * mat_B[520] +
//             mat_A[401] * mat_B[552] +
//             mat_A[402] * mat_B[584] +
//             mat_A[403] * mat_B[616] +
//             mat_A[404] * mat_B[648] +
//             mat_A[405] * mat_B[680] +
//             mat_A[406] * mat_B[712] +
//             mat_A[407] * mat_B[744] +
//             mat_A[408] * mat_B[776] +
//             mat_A[409] * mat_B[808] +
//             mat_A[410] * mat_B[840] +
//             mat_A[411] * mat_B[872] +
//             mat_A[412] * mat_B[904] +
//             mat_A[413] * mat_B[936] +
//             mat_A[414] * mat_B[968] +
//             mat_A[415] * mat_B[1000];
//  mat_C[393] <= 
//             mat_A[384] * mat_B[9] +
//             mat_A[385] * mat_B[41] +
//             mat_A[386] * mat_B[73] +
//             mat_A[387] * mat_B[105] +
//             mat_A[388] * mat_B[137] +
//             mat_A[389] * mat_B[169] +
//             mat_A[390] * mat_B[201] +
//             mat_A[391] * mat_B[233] +
//             mat_A[392] * mat_B[265] +
//             mat_A[393] * mat_B[297] +
//             mat_A[394] * mat_B[329] +
//             mat_A[395] * mat_B[361] +
//             mat_A[396] * mat_B[393] +
//             mat_A[397] * mat_B[425] +
//             mat_A[398] * mat_B[457] +
//             mat_A[399] * mat_B[489] +
//             mat_A[400] * mat_B[521] +
//             mat_A[401] * mat_B[553] +
//             mat_A[402] * mat_B[585] +
//             mat_A[403] * mat_B[617] +
//             mat_A[404] * mat_B[649] +
//             mat_A[405] * mat_B[681] +
//             mat_A[406] * mat_B[713] +
//             mat_A[407] * mat_B[745] +
//             mat_A[408] * mat_B[777] +
//             mat_A[409] * mat_B[809] +
//             mat_A[410] * mat_B[841] +
//             mat_A[411] * mat_B[873] +
//             mat_A[412] * mat_B[905] +
//             mat_A[413] * mat_B[937] +
//             mat_A[414] * mat_B[969] +
//             mat_A[415] * mat_B[1001];
//  mat_C[394] <= 
//             mat_A[384] * mat_B[10] +
//             mat_A[385] * mat_B[42] +
//             mat_A[386] * mat_B[74] +
//             mat_A[387] * mat_B[106] +
//             mat_A[388] * mat_B[138] +
//             mat_A[389] * mat_B[170] +
//             mat_A[390] * mat_B[202] +
//             mat_A[391] * mat_B[234] +
//             mat_A[392] * mat_B[266] +
//             mat_A[393] * mat_B[298] +
//             mat_A[394] * mat_B[330] +
//             mat_A[395] * mat_B[362] +
//             mat_A[396] * mat_B[394] +
//             mat_A[397] * mat_B[426] +
//             mat_A[398] * mat_B[458] +
//             mat_A[399] * mat_B[490] +
//             mat_A[400] * mat_B[522] +
//             mat_A[401] * mat_B[554] +
//             mat_A[402] * mat_B[586] +
//             mat_A[403] * mat_B[618] +
//             mat_A[404] * mat_B[650] +
//             mat_A[405] * mat_B[682] +
//             mat_A[406] * mat_B[714] +
//             mat_A[407] * mat_B[746] +
//             mat_A[408] * mat_B[778] +
//             mat_A[409] * mat_B[810] +
//             mat_A[410] * mat_B[842] +
//             mat_A[411] * mat_B[874] +
//             mat_A[412] * mat_B[906] +
//             mat_A[413] * mat_B[938] +
//             mat_A[414] * mat_B[970] +
//             mat_A[415] * mat_B[1002];
//  mat_C[395] <= 
//             mat_A[384] * mat_B[11] +
//             mat_A[385] * mat_B[43] +
//             mat_A[386] * mat_B[75] +
//             mat_A[387] * mat_B[107] +
//             mat_A[388] * mat_B[139] +
//             mat_A[389] * mat_B[171] +
//             mat_A[390] * mat_B[203] +
//             mat_A[391] * mat_B[235] +
//             mat_A[392] * mat_B[267] +
//             mat_A[393] * mat_B[299] +
//             mat_A[394] * mat_B[331] +
//             mat_A[395] * mat_B[363] +
//             mat_A[396] * mat_B[395] +
//             mat_A[397] * mat_B[427] +
//             mat_A[398] * mat_B[459] +
//             mat_A[399] * mat_B[491] +
//             mat_A[400] * mat_B[523] +
//             mat_A[401] * mat_B[555] +
//             mat_A[402] * mat_B[587] +
//             mat_A[403] * mat_B[619] +
//             mat_A[404] * mat_B[651] +
//             mat_A[405] * mat_B[683] +
//             mat_A[406] * mat_B[715] +
//             mat_A[407] * mat_B[747] +
//             mat_A[408] * mat_B[779] +
//             mat_A[409] * mat_B[811] +
//             mat_A[410] * mat_B[843] +
//             mat_A[411] * mat_B[875] +
//             mat_A[412] * mat_B[907] +
//             mat_A[413] * mat_B[939] +
//             mat_A[414] * mat_B[971] +
//             mat_A[415] * mat_B[1003];
//  mat_C[396] <= 
//             mat_A[384] * mat_B[12] +
//             mat_A[385] * mat_B[44] +
//             mat_A[386] * mat_B[76] +
//             mat_A[387] * mat_B[108] +
//             mat_A[388] * mat_B[140] +
//             mat_A[389] * mat_B[172] +
//             mat_A[390] * mat_B[204] +
//             mat_A[391] * mat_B[236] +
//             mat_A[392] * mat_B[268] +
//             mat_A[393] * mat_B[300] +
//             mat_A[394] * mat_B[332] +
//             mat_A[395] * mat_B[364] +
//             mat_A[396] * mat_B[396] +
//             mat_A[397] * mat_B[428] +
//             mat_A[398] * mat_B[460] +
//             mat_A[399] * mat_B[492] +
//             mat_A[400] * mat_B[524] +
//             mat_A[401] * mat_B[556] +
//             mat_A[402] * mat_B[588] +
//             mat_A[403] * mat_B[620] +
//             mat_A[404] * mat_B[652] +
//             mat_A[405] * mat_B[684] +
//             mat_A[406] * mat_B[716] +
//             mat_A[407] * mat_B[748] +
//             mat_A[408] * mat_B[780] +
//             mat_A[409] * mat_B[812] +
//             mat_A[410] * mat_B[844] +
//             mat_A[411] * mat_B[876] +
//             mat_A[412] * mat_B[908] +
//             mat_A[413] * mat_B[940] +
//             mat_A[414] * mat_B[972] +
//             mat_A[415] * mat_B[1004];
//  mat_C[397] <= 
//             mat_A[384] * mat_B[13] +
//             mat_A[385] * mat_B[45] +
//             mat_A[386] * mat_B[77] +
//             mat_A[387] * mat_B[109] +
//             mat_A[388] * mat_B[141] +
//             mat_A[389] * mat_B[173] +
//             mat_A[390] * mat_B[205] +
//             mat_A[391] * mat_B[237] +
//             mat_A[392] * mat_B[269] +
//             mat_A[393] * mat_B[301] +
//             mat_A[394] * mat_B[333] +
//             mat_A[395] * mat_B[365] +
//             mat_A[396] * mat_B[397] +
//             mat_A[397] * mat_B[429] +
//             mat_A[398] * mat_B[461] +
//             mat_A[399] * mat_B[493] +
//             mat_A[400] * mat_B[525] +
//             mat_A[401] * mat_B[557] +
//             mat_A[402] * mat_B[589] +
//             mat_A[403] * mat_B[621] +
//             mat_A[404] * mat_B[653] +
//             mat_A[405] * mat_B[685] +
//             mat_A[406] * mat_B[717] +
//             mat_A[407] * mat_B[749] +
//             mat_A[408] * mat_B[781] +
//             mat_A[409] * mat_B[813] +
//             mat_A[410] * mat_B[845] +
//             mat_A[411] * mat_B[877] +
//             mat_A[412] * mat_B[909] +
//             mat_A[413] * mat_B[941] +
//             mat_A[414] * mat_B[973] +
//             mat_A[415] * mat_B[1005];
//  mat_C[398] <= 
//             mat_A[384] * mat_B[14] +
//             mat_A[385] * mat_B[46] +
//             mat_A[386] * mat_B[78] +
//             mat_A[387] * mat_B[110] +
//             mat_A[388] * mat_B[142] +
//             mat_A[389] * mat_B[174] +
//             mat_A[390] * mat_B[206] +
//             mat_A[391] * mat_B[238] +
//             mat_A[392] * mat_B[270] +
//             mat_A[393] * mat_B[302] +
//             mat_A[394] * mat_B[334] +
//             mat_A[395] * mat_B[366] +
//             mat_A[396] * mat_B[398] +
//             mat_A[397] * mat_B[430] +
//             mat_A[398] * mat_B[462] +
//             mat_A[399] * mat_B[494] +
//             mat_A[400] * mat_B[526] +
//             mat_A[401] * mat_B[558] +
//             mat_A[402] * mat_B[590] +
//             mat_A[403] * mat_B[622] +
//             mat_A[404] * mat_B[654] +
//             mat_A[405] * mat_B[686] +
//             mat_A[406] * mat_B[718] +
//             mat_A[407] * mat_B[750] +
//             mat_A[408] * mat_B[782] +
//             mat_A[409] * mat_B[814] +
//             mat_A[410] * mat_B[846] +
//             mat_A[411] * mat_B[878] +
//             mat_A[412] * mat_B[910] +
//             mat_A[413] * mat_B[942] +
//             mat_A[414] * mat_B[974] +
//             mat_A[415] * mat_B[1006];
//  mat_C[399] <= 
//             mat_A[384] * mat_B[15] +
//             mat_A[385] * mat_B[47] +
//             mat_A[386] * mat_B[79] +
//             mat_A[387] * mat_B[111] +
//             mat_A[388] * mat_B[143] +
//             mat_A[389] * mat_B[175] +
//             mat_A[390] * mat_B[207] +
//             mat_A[391] * mat_B[239] +
//             mat_A[392] * mat_B[271] +
//             mat_A[393] * mat_B[303] +
//             mat_A[394] * mat_B[335] +
//             mat_A[395] * mat_B[367] +
//             mat_A[396] * mat_B[399] +
//             mat_A[397] * mat_B[431] +
//             mat_A[398] * mat_B[463] +
//             mat_A[399] * mat_B[495] +
//             mat_A[400] * mat_B[527] +
//             mat_A[401] * mat_B[559] +
//             mat_A[402] * mat_B[591] +
//             mat_A[403] * mat_B[623] +
//             mat_A[404] * mat_B[655] +
//             mat_A[405] * mat_B[687] +
//             mat_A[406] * mat_B[719] +
//             mat_A[407] * mat_B[751] +
//             mat_A[408] * mat_B[783] +
//             mat_A[409] * mat_B[815] +
//             mat_A[410] * mat_B[847] +
//             mat_A[411] * mat_B[879] +
//             mat_A[412] * mat_B[911] +
//             mat_A[413] * mat_B[943] +
//             mat_A[414] * mat_B[975] +
//             mat_A[415] * mat_B[1007];
//  mat_C[400] <= 
//             mat_A[384] * mat_B[16] +
//             mat_A[385] * mat_B[48] +
//             mat_A[386] * mat_B[80] +
//             mat_A[387] * mat_B[112] +
//             mat_A[388] * mat_B[144] +
//             mat_A[389] * mat_B[176] +
//             mat_A[390] * mat_B[208] +
//             mat_A[391] * mat_B[240] +
//             mat_A[392] * mat_B[272] +
//             mat_A[393] * mat_B[304] +
//             mat_A[394] * mat_B[336] +
//             mat_A[395] * mat_B[368] +
//             mat_A[396] * mat_B[400] +
//             mat_A[397] * mat_B[432] +
//             mat_A[398] * mat_B[464] +
//             mat_A[399] * mat_B[496] +
//             mat_A[400] * mat_B[528] +
//             mat_A[401] * mat_B[560] +
//             mat_A[402] * mat_B[592] +
//             mat_A[403] * mat_B[624] +
//             mat_A[404] * mat_B[656] +
//             mat_A[405] * mat_B[688] +
//             mat_A[406] * mat_B[720] +
//             mat_A[407] * mat_B[752] +
//             mat_A[408] * mat_B[784] +
//             mat_A[409] * mat_B[816] +
//             mat_A[410] * mat_B[848] +
//             mat_A[411] * mat_B[880] +
//             mat_A[412] * mat_B[912] +
//             mat_A[413] * mat_B[944] +
//             mat_A[414] * mat_B[976] +
//             mat_A[415] * mat_B[1008];
//  mat_C[401] <= 
//             mat_A[384] * mat_B[17] +
//             mat_A[385] * mat_B[49] +
//             mat_A[386] * mat_B[81] +
//             mat_A[387] * mat_B[113] +
//             mat_A[388] * mat_B[145] +
//             mat_A[389] * mat_B[177] +
//             mat_A[390] * mat_B[209] +
//             mat_A[391] * mat_B[241] +
//             mat_A[392] * mat_B[273] +
//             mat_A[393] * mat_B[305] +
//             mat_A[394] * mat_B[337] +
//             mat_A[395] * mat_B[369] +
//             mat_A[396] * mat_B[401] +
//             mat_A[397] * mat_B[433] +
//             mat_A[398] * mat_B[465] +
//             mat_A[399] * mat_B[497] +
//             mat_A[400] * mat_B[529] +
//             mat_A[401] * mat_B[561] +
//             mat_A[402] * mat_B[593] +
//             mat_A[403] * mat_B[625] +
//             mat_A[404] * mat_B[657] +
//             mat_A[405] * mat_B[689] +
//             mat_A[406] * mat_B[721] +
//             mat_A[407] * mat_B[753] +
//             mat_A[408] * mat_B[785] +
//             mat_A[409] * mat_B[817] +
//             mat_A[410] * mat_B[849] +
//             mat_A[411] * mat_B[881] +
//             mat_A[412] * mat_B[913] +
//             mat_A[413] * mat_B[945] +
//             mat_A[414] * mat_B[977] +
//             mat_A[415] * mat_B[1009];
//  mat_C[402] <= 
//             mat_A[384] * mat_B[18] +
//             mat_A[385] * mat_B[50] +
//             mat_A[386] * mat_B[82] +
//             mat_A[387] * mat_B[114] +
//             mat_A[388] * mat_B[146] +
//             mat_A[389] * mat_B[178] +
//             mat_A[390] * mat_B[210] +
//             mat_A[391] * mat_B[242] +
//             mat_A[392] * mat_B[274] +
//             mat_A[393] * mat_B[306] +
//             mat_A[394] * mat_B[338] +
//             mat_A[395] * mat_B[370] +
//             mat_A[396] * mat_B[402] +
//             mat_A[397] * mat_B[434] +
//             mat_A[398] * mat_B[466] +
//             mat_A[399] * mat_B[498] +
//             mat_A[400] * mat_B[530] +
//             mat_A[401] * mat_B[562] +
//             mat_A[402] * mat_B[594] +
//             mat_A[403] * mat_B[626] +
//             mat_A[404] * mat_B[658] +
//             mat_A[405] * mat_B[690] +
//             mat_A[406] * mat_B[722] +
//             mat_A[407] * mat_B[754] +
//             mat_A[408] * mat_B[786] +
//             mat_A[409] * mat_B[818] +
//             mat_A[410] * mat_B[850] +
//             mat_A[411] * mat_B[882] +
//             mat_A[412] * mat_B[914] +
//             mat_A[413] * mat_B[946] +
//             mat_A[414] * mat_B[978] +
//             mat_A[415] * mat_B[1010];
//  mat_C[403] <= 
//             mat_A[384] * mat_B[19] +
//             mat_A[385] * mat_B[51] +
//             mat_A[386] * mat_B[83] +
//             mat_A[387] * mat_B[115] +
//             mat_A[388] * mat_B[147] +
//             mat_A[389] * mat_B[179] +
//             mat_A[390] * mat_B[211] +
//             mat_A[391] * mat_B[243] +
//             mat_A[392] * mat_B[275] +
//             mat_A[393] * mat_B[307] +
//             mat_A[394] * mat_B[339] +
//             mat_A[395] * mat_B[371] +
//             mat_A[396] * mat_B[403] +
//             mat_A[397] * mat_B[435] +
//             mat_A[398] * mat_B[467] +
//             mat_A[399] * mat_B[499] +
//             mat_A[400] * mat_B[531] +
//             mat_A[401] * mat_B[563] +
//             mat_A[402] * mat_B[595] +
//             mat_A[403] * mat_B[627] +
//             mat_A[404] * mat_B[659] +
//             mat_A[405] * mat_B[691] +
//             mat_A[406] * mat_B[723] +
//             mat_A[407] * mat_B[755] +
//             mat_A[408] * mat_B[787] +
//             mat_A[409] * mat_B[819] +
//             mat_A[410] * mat_B[851] +
//             mat_A[411] * mat_B[883] +
//             mat_A[412] * mat_B[915] +
//             mat_A[413] * mat_B[947] +
//             mat_A[414] * mat_B[979] +
//             mat_A[415] * mat_B[1011];
//  mat_C[404] <= 
//             mat_A[384] * mat_B[20] +
//             mat_A[385] * mat_B[52] +
//             mat_A[386] * mat_B[84] +
//             mat_A[387] * mat_B[116] +
//             mat_A[388] * mat_B[148] +
//             mat_A[389] * mat_B[180] +
//             mat_A[390] * mat_B[212] +
//             mat_A[391] * mat_B[244] +
//             mat_A[392] * mat_B[276] +
//             mat_A[393] * mat_B[308] +
//             mat_A[394] * mat_B[340] +
//             mat_A[395] * mat_B[372] +
//             mat_A[396] * mat_B[404] +
//             mat_A[397] * mat_B[436] +
//             mat_A[398] * mat_B[468] +
//             mat_A[399] * mat_B[500] +
//             mat_A[400] * mat_B[532] +
//             mat_A[401] * mat_B[564] +
//             mat_A[402] * mat_B[596] +
//             mat_A[403] * mat_B[628] +
//             mat_A[404] * mat_B[660] +
//             mat_A[405] * mat_B[692] +
//             mat_A[406] * mat_B[724] +
//             mat_A[407] * mat_B[756] +
//             mat_A[408] * mat_B[788] +
//             mat_A[409] * mat_B[820] +
//             mat_A[410] * mat_B[852] +
//             mat_A[411] * mat_B[884] +
//             mat_A[412] * mat_B[916] +
//             mat_A[413] * mat_B[948] +
//             mat_A[414] * mat_B[980] +
//             mat_A[415] * mat_B[1012];
//  mat_C[405] <= 
//             mat_A[384] * mat_B[21] +
//             mat_A[385] * mat_B[53] +
//             mat_A[386] * mat_B[85] +
//             mat_A[387] * mat_B[117] +
//             mat_A[388] * mat_B[149] +
//             mat_A[389] * mat_B[181] +
//             mat_A[390] * mat_B[213] +
//             mat_A[391] * mat_B[245] +
//             mat_A[392] * mat_B[277] +
//             mat_A[393] * mat_B[309] +
//             mat_A[394] * mat_B[341] +
//             mat_A[395] * mat_B[373] +
//             mat_A[396] * mat_B[405] +
//             mat_A[397] * mat_B[437] +
//             mat_A[398] * mat_B[469] +
//             mat_A[399] * mat_B[501] +
//             mat_A[400] * mat_B[533] +
//             mat_A[401] * mat_B[565] +
//             mat_A[402] * mat_B[597] +
//             mat_A[403] * mat_B[629] +
//             mat_A[404] * mat_B[661] +
//             mat_A[405] * mat_B[693] +
//             mat_A[406] * mat_B[725] +
//             mat_A[407] * mat_B[757] +
//             mat_A[408] * mat_B[789] +
//             mat_A[409] * mat_B[821] +
//             mat_A[410] * mat_B[853] +
//             mat_A[411] * mat_B[885] +
//             mat_A[412] * mat_B[917] +
//             mat_A[413] * mat_B[949] +
//             mat_A[414] * mat_B[981] +
//             mat_A[415] * mat_B[1013];
//  mat_C[406] <= 
//             mat_A[384] * mat_B[22] +
//             mat_A[385] * mat_B[54] +
//             mat_A[386] * mat_B[86] +
//             mat_A[387] * mat_B[118] +
//             mat_A[388] * mat_B[150] +
//             mat_A[389] * mat_B[182] +
//             mat_A[390] * mat_B[214] +
//             mat_A[391] * mat_B[246] +
//             mat_A[392] * mat_B[278] +
//             mat_A[393] * mat_B[310] +
//             mat_A[394] * mat_B[342] +
//             mat_A[395] * mat_B[374] +
//             mat_A[396] * mat_B[406] +
//             mat_A[397] * mat_B[438] +
//             mat_A[398] * mat_B[470] +
//             mat_A[399] * mat_B[502] +
//             mat_A[400] * mat_B[534] +
//             mat_A[401] * mat_B[566] +
//             mat_A[402] * mat_B[598] +
//             mat_A[403] * mat_B[630] +
//             mat_A[404] * mat_B[662] +
//             mat_A[405] * mat_B[694] +
//             mat_A[406] * mat_B[726] +
//             mat_A[407] * mat_B[758] +
//             mat_A[408] * mat_B[790] +
//             mat_A[409] * mat_B[822] +
//             mat_A[410] * mat_B[854] +
//             mat_A[411] * mat_B[886] +
//             mat_A[412] * mat_B[918] +
//             mat_A[413] * mat_B[950] +
//             mat_A[414] * mat_B[982] +
//             mat_A[415] * mat_B[1014];
//  mat_C[407] <= 
//             mat_A[384] * mat_B[23] +
//             mat_A[385] * mat_B[55] +
//             mat_A[386] * mat_B[87] +
//             mat_A[387] * mat_B[119] +
//             mat_A[388] * mat_B[151] +
//             mat_A[389] * mat_B[183] +
//             mat_A[390] * mat_B[215] +
//             mat_A[391] * mat_B[247] +
//             mat_A[392] * mat_B[279] +
//             mat_A[393] * mat_B[311] +
//             mat_A[394] * mat_B[343] +
//             mat_A[395] * mat_B[375] +
//             mat_A[396] * mat_B[407] +
//             mat_A[397] * mat_B[439] +
//             mat_A[398] * mat_B[471] +
//             mat_A[399] * mat_B[503] +
//             mat_A[400] * mat_B[535] +
//             mat_A[401] * mat_B[567] +
//             mat_A[402] * mat_B[599] +
//             mat_A[403] * mat_B[631] +
//             mat_A[404] * mat_B[663] +
//             mat_A[405] * mat_B[695] +
//             mat_A[406] * mat_B[727] +
//             mat_A[407] * mat_B[759] +
//             mat_A[408] * mat_B[791] +
//             mat_A[409] * mat_B[823] +
//             mat_A[410] * mat_B[855] +
//             mat_A[411] * mat_B[887] +
//             mat_A[412] * mat_B[919] +
//             mat_A[413] * mat_B[951] +
//             mat_A[414] * mat_B[983] +
//             mat_A[415] * mat_B[1015];
//  mat_C[408] <= 
//             mat_A[384] * mat_B[24] +
//             mat_A[385] * mat_B[56] +
//             mat_A[386] * mat_B[88] +
//             mat_A[387] * mat_B[120] +
//             mat_A[388] * mat_B[152] +
//             mat_A[389] * mat_B[184] +
//             mat_A[390] * mat_B[216] +
//             mat_A[391] * mat_B[248] +
//             mat_A[392] * mat_B[280] +
//             mat_A[393] * mat_B[312] +
//             mat_A[394] * mat_B[344] +
//             mat_A[395] * mat_B[376] +
//             mat_A[396] * mat_B[408] +
//             mat_A[397] * mat_B[440] +
//             mat_A[398] * mat_B[472] +
//             mat_A[399] * mat_B[504] +
//             mat_A[400] * mat_B[536] +
//             mat_A[401] * mat_B[568] +
//             mat_A[402] * mat_B[600] +
//             mat_A[403] * mat_B[632] +
//             mat_A[404] * mat_B[664] +
//             mat_A[405] * mat_B[696] +
//             mat_A[406] * mat_B[728] +
//             mat_A[407] * mat_B[760] +
//             mat_A[408] * mat_B[792] +
//             mat_A[409] * mat_B[824] +
//             mat_A[410] * mat_B[856] +
//             mat_A[411] * mat_B[888] +
//             mat_A[412] * mat_B[920] +
//             mat_A[413] * mat_B[952] +
//             mat_A[414] * mat_B[984] +
//             mat_A[415] * mat_B[1016];
//  mat_C[409] <= 
//             mat_A[384] * mat_B[25] +
//             mat_A[385] * mat_B[57] +
//             mat_A[386] * mat_B[89] +
//             mat_A[387] * mat_B[121] +
//             mat_A[388] * mat_B[153] +
//             mat_A[389] * mat_B[185] +
//             mat_A[390] * mat_B[217] +
//             mat_A[391] * mat_B[249] +
//             mat_A[392] * mat_B[281] +
//             mat_A[393] * mat_B[313] +
//             mat_A[394] * mat_B[345] +
//             mat_A[395] * mat_B[377] +
//             mat_A[396] * mat_B[409] +
//             mat_A[397] * mat_B[441] +
//             mat_A[398] * mat_B[473] +
//             mat_A[399] * mat_B[505] +
//             mat_A[400] * mat_B[537] +
//             mat_A[401] * mat_B[569] +
//             mat_A[402] * mat_B[601] +
//             mat_A[403] * mat_B[633] +
//             mat_A[404] * mat_B[665] +
//             mat_A[405] * mat_B[697] +
//             mat_A[406] * mat_B[729] +
//             mat_A[407] * mat_B[761] +
//             mat_A[408] * mat_B[793] +
//             mat_A[409] * mat_B[825] +
//             mat_A[410] * mat_B[857] +
//             mat_A[411] * mat_B[889] +
//             mat_A[412] * mat_B[921] +
//             mat_A[413] * mat_B[953] +
//             mat_A[414] * mat_B[985] +
//             mat_A[415] * mat_B[1017];
//  mat_C[410] <= 
//             mat_A[384] * mat_B[26] +
//             mat_A[385] * mat_B[58] +
//             mat_A[386] * mat_B[90] +
//             mat_A[387] * mat_B[122] +
//             mat_A[388] * mat_B[154] +
//             mat_A[389] * mat_B[186] +
//             mat_A[390] * mat_B[218] +
//             mat_A[391] * mat_B[250] +
//             mat_A[392] * mat_B[282] +
//             mat_A[393] * mat_B[314] +
//             mat_A[394] * mat_B[346] +
//             mat_A[395] * mat_B[378] +
//             mat_A[396] * mat_B[410] +
//             mat_A[397] * mat_B[442] +
//             mat_A[398] * mat_B[474] +
//             mat_A[399] * mat_B[506] +
//             mat_A[400] * mat_B[538] +
//             mat_A[401] * mat_B[570] +
//             mat_A[402] * mat_B[602] +
//             mat_A[403] * mat_B[634] +
//             mat_A[404] * mat_B[666] +
//             mat_A[405] * mat_B[698] +
//             mat_A[406] * mat_B[730] +
//             mat_A[407] * mat_B[762] +
//             mat_A[408] * mat_B[794] +
//             mat_A[409] * mat_B[826] +
//             mat_A[410] * mat_B[858] +
//             mat_A[411] * mat_B[890] +
//             mat_A[412] * mat_B[922] +
//             mat_A[413] * mat_B[954] +
//             mat_A[414] * mat_B[986] +
//             mat_A[415] * mat_B[1018];
//  mat_C[411] <= 
//             mat_A[384] * mat_B[27] +
//             mat_A[385] * mat_B[59] +
//             mat_A[386] * mat_B[91] +
//             mat_A[387] * mat_B[123] +
//             mat_A[388] * mat_B[155] +
//             mat_A[389] * mat_B[187] +
//             mat_A[390] * mat_B[219] +
//             mat_A[391] * mat_B[251] +
//             mat_A[392] * mat_B[283] +
//             mat_A[393] * mat_B[315] +
//             mat_A[394] * mat_B[347] +
//             mat_A[395] * mat_B[379] +
//             mat_A[396] * mat_B[411] +
//             mat_A[397] * mat_B[443] +
//             mat_A[398] * mat_B[475] +
//             mat_A[399] * mat_B[507] +
//             mat_A[400] * mat_B[539] +
//             mat_A[401] * mat_B[571] +
//             mat_A[402] * mat_B[603] +
//             mat_A[403] * mat_B[635] +
//             mat_A[404] * mat_B[667] +
//             mat_A[405] * mat_B[699] +
//             mat_A[406] * mat_B[731] +
//             mat_A[407] * mat_B[763] +
//             mat_A[408] * mat_B[795] +
//             mat_A[409] * mat_B[827] +
//             mat_A[410] * mat_B[859] +
//             mat_A[411] * mat_B[891] +
//             mat_A[412] * mat_B[923] +
//             mat_A[413] * mat_B[955] +
//             mat_A[414] * mat_B[987] +
//             mat_A[415] * mat_B[1019];
//  mat_C[412] <= 
//             mat_A[384] * mat_B[28] +
//             mat_A[385] * mat_B[60] +
//             mat_A[386] * mat_B[92] +
//             mat_A[387] * mat_B[124] +
//             mat_A[388] * mat_B[156] +
//             mat_A[389] * mat_B[188] +
//             mat_A[390] * mat_B[220] +
//             mat_A[391] * mat_B[252] +
//             mat_A[392] * mat_B[284] +
//             mat_A[393] * mat_B[316] +
//             mat_A[394] * mat_B[348] +
//             mat_A[395] * mat_B[380] +
//             mat_A[396] * mat_B[412] +
//             mat_A[397] * mat_B[444] +
//             mat_A[398] * mat_B[476] +
//             mat_A[399] * mat_B[508] +
//             mat_A[400] * mat_B[540] +
//             mat_A[401] * mat_B[572] +
//             mat_A[402] * mat_B[604] +
//             mat_A[403] * mat_B[636] +
//             mat_A[404] * mat_B[668] +
//             mat_A[405] * mat_B[700] +
//             mat_A[406] * mat_B[732] +
//             mat_A[407] * mat_B[764] +
//             mat_A[408] * mat_B[796] +
//             mat_A[409] * mat_B[828] +
//             mat_A[410] * mat_B[860] +
//             mat_A[411] * mat_B[892] +
//             mat_A[412] * mat_B[924] +
//             mat_A[413] * mat_B[956] +
//             mat_A[414] * mat_B[988] +
//             mat_A[415] * mat_B[1020];
//  mat_C[413] <= 
//             mat_A[384] * mat_B[29] +
//             mat_A[385] * mat_B[61] +
//             mat_A[386] * mat_B[93] +
//             mat_A[387] * mat_B[125] +
//             mat_A[388] * mat_B[157] +
//             mat_A[389] * mat_B[189] +
//             mat_A[390] * mat_B[221] +
//             mat_A[391] * mat_B[253] +
//             mat_A[392] * mat_B[285] +
//             mat_A[393] * mat_B[317] +
//             mat_A[394] * mat_B[349] +
//             mat_A[395] * mat_B[381] +
//             mat_A[396] * mat_B[413] +
//             mat_A[397] * mat_B[445] +
//             mat_A[398] * mat_B[477] +
//             mat_A[399] * mat_B[509] +
//             mat_A[400] * mat_B[541] +
//             mat_A[401] * mat_B[573] +
//             mat_A[402] * mat_B[605] +
//             mat_A[403] * mat_B[637] +
//             mat_A[404] * mat_B[669] +
//             mat_A[405] * mat_B[701] +
//             mat_A[406] * mat_B[733] +
//             mat_A[407] * mat_B[765] +
//             mat_A[408] * mat_B[797] +
//             mat_A[409] * mat_B[829] +
//             mat_A[410] * mat_B[861] +
//             mat_A[411] * mat_B[893] +
//             mat_A[412] * mat_B[925] +
//             mat_A[413] * mat_B[957] +
//             mat_A[414] * mat_B[989] +
//             mat_A[415] * mat_B[1021];
//  mat_C[414] <= 
//             mat_A[384] * mat_B[30] +
//             mat_A[385] * mat_B[62] +
//             mat_A[386] * mat_B[94] +
//             mat_A[387] * mat_B[126] +
//             mat_A[388] * mat_B[158] +
//             mat_A[389] * mat_B[190] +
//             mat_A[390] * mat_B[222] +
//             mat_A[391] * mat_B[254] +
//             mat_A[392] * mat_B[286] +
//             mat_A[393] * mat_B[318] +
//             mat_A[394] * mat_B[350] +
//             mat_A[395] * mat_B[382] +
//             mat_A[396] * mat_B[414] +
//             mat_A[397] * mat_B[446] +
//             mat_A[398] * mat_B[478] +
//             mat_A[399] * mat_B[510] +
//             mat_A[400] * mat_B[542] +
//             mat_A[401] * mat_B[574] +
//             mat_A[402] * mat_B[606] +
//             mat_A[403] * mat_B[638] +
//             mat_A[404] * mat_B[670] +
//             mat_A[405] * mat_B[702] +
//             mat_A[406] * mat_B[734] +
//             mat_A[407] * mat_B[766] +
//             mat_A[408] * mat_B[798] +
//             mat_A[409] * mat_B[830] +
//             mat_A[410] * mat_B[862] +
//             mat_A[411] * mat_B[894] +
//             mat_A[412] * mat_B[926] +
//             mat_A[413] * mat_B[958] +
//             mat_A[414] * mat_B[990] +
//             mat_A[415] * mat_B[1022];
//  mat_C[415] <= 
//             mat_A[384] * mat_B[31] +
//             mat_A[385] * mat_B[63] +
//             mat_A[386] * mat_B[95] +
//             mat_A[387] * mat_B[127] +
//             mat_A[388] * mat_B[159] +
//             mat_A[389] * mat_B[191] +
//             mat_A[390] * mat_B[223] +
//             mat_A[391] * mat_B[255] +
//             mat_A[392] * mat_B[287] +
//             mat_A[393] * mat_B[319] +
//             mat_A[394] * mat_B[351] +
//             mat_A[395] * mat_B[383] +
//             mat_A[396] * mat_B[415] +
//             mat_A[397] * mat_B[447] +
//             mat_A[398] * mat_B[479] +
//             mat_A[399] * mat_B[511] +
//             mat_A[400] * mat_B[543] +
//             mat_A[401] * mat_B[575] +
//             mat_A[402] * mat_B[607] +
//             mat_A[403] * mat_B[639] +
//             mat_A[404] * mat_B[671] +
//             mat_A[405] * mat_B[703] +
//             mat_A[406] * mat_B[735] +
//             mat_A[407] * mat_B[767] +
//             mat_A[408] * mat_B[799] +
//             mat_A[409] * mat_B[831] +
//             mat_A[410] * mat_B[863] +
//             mat_A[411] * mat_B[895] +
//             mat_A[412] * mat_B[927] +
//             mat_A[413] * mat_B[959] +
//             mat_A[414] * mat_B[991] +
//             mat_A[415] * mat_B[1023];
//  mat_C[416] <= 
//             mat_A[416] * mat_B[0] +
//             mat_A[417] * mat_B[32] +
//             mat_A[418] * mat_B[64] +
//             mat_A[419] * mat_B[96] +
//             mat_A[420] * mat_B[128] +
//             mat_A[421] * mat_B[160] +
//             mat_A[422] * mat_B[192] +
//             mat_A[423] * mat_B[224] +
//             mat_A[424] * mat_B[256] +
//             mat_A[425] * mat_B[288] +
//             mat_A[426] * mat_B[320] +
//             mat_A[427] * mat_B[352] +
//             mat_A[428] * mat_B[384] +
//             mat_A[429] * mat_B[416] +
//             mat_A[430] * mat_B[448] +
//             mat_A[431] * mat_B[480] +
//             mat_A[432] * mat_B[512] +
//             mat_A[433] * mat_B[544] +
//             mat_A[434] * mat_B[576] +
//             mat_A[435] * mat_B[608] +
//             mat_A[436] * mat_B[640] +
//             mat_A[437] * mat_B[672] +
//             mat_A[438] * mat_B[704] +
//             mat_A[439] * mat_B[736] +
//             mat_A[440] * mat_B[768] +
//             mat_A[441] * mat_B[800] +
//             mat_A[442] * mat_B[832] +
//             mat_A[443] * mat_B[864] +
//             mat_A[444] * mat_B[896] +
//             mat_A[445] * mat_B[928] +
//             mat_A[446] * mat_B[960] +
//             mat_A[447] * mat_B[992];
//  mat_C[417] <= 
//             mat_A[416] * mat_B[1] +
//             mat_A[417] * mat_B[33] +
//             mat_A[418] * mat_B[65] +
//             mat_A[419] * mat_B[97] +
//             mat_A[420] * mat_B[129] +
//             mat_A[421] * mat_B[161] +
//             mat_A[422] * mat_B[193] +
//             mat_A[423] * mat_B[225] +
//             mat_A[424] * mat_B[257] +
//             mat_A[425] * mat_B[289] +
//             mat_A[426] * mat_B[321] +
//             mat_A[427] * mat_B[353] +
//             mat_A[428] * mat_B[385] +
//             mat_A[429] * mat_B[417] +
//             mat_A[430] * mat_B[449] +
//             mat_A[431] * mat_B[481] +
//             mat_A[432] * mat_B[513] +
//             mat_A[433] * mat_B[545] +
//             mat_A[434] * mat_B[577] +
//             mat_A[435] * mat_B[609] +
//             mat_A[436] * mat_B[641] +
//             mat_A[437] * mat_B[673] +
//             mat_A[438] * mat_B[705] +
//             mat_A[439] * mat_B[737] +
//             mat_A[440] * mat_B[769] +
//             mat_A[441] * mat_B[801] +
//             mat_A[442] * mat_B[833] +
//             mat_A[443] * mat_B[865] +
//             mat_A[444] * mat_B[897] +
//             mat_A[445] * mat_B[929] +
//             mat_A[446] * mat_B[961] +
//             mat_A[447] * mat_B[993];
//  mat_C[418] <= 
//             mat_A[416] * mat_B[2] +
//             mat_A[417] * mat_B[34] +
//             mat_A[418] * mat_B[66] +
//             mat_A[419] * mat_B[98] +
//             mat_A[420] * mat_B[130] +
//             mat_A[421] * mat_B[162] +
//             mat_A[422] * mat_B[194] +
//             mat_A[423] * mat_B[226] +
//             mat_A[424] * mat_B[258] +
//             mat_A[425] * mat_B[290] +
//             mat_A[426] * mat_B[322] +
//             mat_A[427] * mat_B[354] +
//             mat_A[428] * mat_B[386] +
//             mat_A[429] * mat_B[418] +
//             mat_A[430] * mat_B[450] +
//             mat_A[431] * mat_B[482] +
//             mat_A[432] * mat_B[514] +
//             mat_A[433] * mat_B[546] +
//             mat_A[434] * mat_B[578] +
//             mat_A[435] * mat_B[610] +
//             mat_A[436] * mat_B[642] +
//             mat_A[437] * mat_B[674] +
//             mat_A[438] * mat_B[706] +
//             mat_A[439] * mat_B[738] +
//             mat_A[440] * mat_B[770] +
//             mat_A[441] * mat_B[802] +
//             mat_A[442] * mat_B[834] +
//             mat_A[443] * mat_B[866] +
//             mat_A[444] * mat_B[898] +
//             mat_A[445] * mat_B[930] +
//             mat_A[446] * mat_B[962] +
//             mat_A[447] * mat_B[994];
//  mat_C[419] <= 
//             mat_A[416] * mat_B[3] +
//             mat_A[417] * mat_B[35] +
//             mat_A[418] * mat_B[67] +
//             mat_A[419] * mat_B[99] +
//             mat_A[420] * mat_B[131] +
//             mat_A[421] * mat_B[163] +
//             mat_A[422] * mat_B[195] +
//             mat_A[423] * mat_B[227] +
//             mat_A[424] * mat_B[259] +
//             mat_A[425] * mat_B[291] +
//             mat_A[426] * mat_B[323] +
//             mat_A[427] * mat_B[355] +
//             mat_A[428] * mat_B[387] +
//             mat_A[429] * mat_B[419] +
//             mat_A[430] * mat_B[451] +
//             mat_A[431] * mat_B[483] +
//             mat_A[432] * mat_B[515] +
//             mat_A[433] * mat_B[547] +
//             mat_A[434] * mat_B[579] +
//             mat_A[435] * mat_B[611] +
//             mat_A[436] * mat_B[643] +
//             mat_A[437] * mat_B[675] +
//             mat_A[438] * mat_B[707] +
//             mat_A[439] * mat_B[739] +
//             mat_A[440] * mat_B[771] +
//             mat_A[441] * mat_B[803] +
//             mat_A[442] * mat_B[835] +
//             mat_A[443] * mat_B[867] +
//             mat_A[444] * mat_B[899] +
//             mat_A[445] * mat_B[931] +
//             mat_A[446] * mat_B[963] +
//             mat_A[447] * mat_B[995];
//  mat_C[420] <= 
//             mat_A[416] * mat_B[4] +
//             mat_A[417] * mat_B[36] +
//             mat_A[418] * mat_B[68] +
//             mat_A[419] * mat_B[100] +
//             mat_A[420] * mat_B[132] +
//             mat_A[421] * mat_B[164] +
//             mat_A[422] * mat_B[196] +
//             mat_A[423] * mat_B[228] +
//             mat_A[424] * mat_B[260] +
//             mat_A[425] * mat_B[292] +
//             mat_A[426] * mat_B[324] +
//             mat_A[427] * mat_B[356] +
//             mat_A[428] * mat_B[388] +
//             mat_A[429] * mat_B[420] +
//             mat_A[430] * mat_B[452] +
//             mat_A[431] * mat_B[484] +
//             mat_A[432] * mat_B[516] +
//             mat_A[433] * mat_B[548] +
//             mat_A[434] * mat_B[580] +
//             mat_A[435] * mat_B[612] +
//             mat_A[436] * mat_B[644] +
//             mat_A[437] * mat_B[676] +
//             mat_A[438] * mat_B[708] +
//             mat_A[439] * mat_B[740] +
//             mat_A[440] * mat_B[772] +
//             mat_A[441] * mat_B[804] +
//             mat_A[442] * mat_B[836] +
//             mat_A[443] * mat_B[868] +
//             mat_A[444] * mat_B[900] +
//             mat_A[445] * mat_B[932] +
//             mat_A[446] * mat_B[964] +
//             mat_A[447] * mat_B[996];
//  mat_C[421] <= 
//             mat_A[416] * mat_B[5] +
//             mat_A[417] * mat_B[37] +
//             mat_A[418] * mat_B[69] +
//             mat_A[419] * mat_B[101] +
//             mat_A[420] * mat_B[133] +
//             mat_A[421] * mat_B[165] +
//             mat_A[422] * mat_B[197] +
//             mat_A[423] * mat_B[229] +
//             mat_A[424] * mat_B[261] +
//             mat_A[425] * mat_B[293] +
//             mat_A[426] * mat_B[325] +
//             mat_A[427] * mat_B[357] +
//             mat_A[428] * mat_B[389] +
//             mat_A[429] * mat_B[421] +
//             mat_A[430] * mat_B[453] +
//             mat_A[431] * mat_B[485] +
//             mat_A[432] * mat_B[517] +
//             mat_A[433] * mat_B[549] +
//             mat_A[434] * mat_B[581] +
//             mat_A[435] * mat_B[613] +
//             mat_A[436] * mat_B[645] +
//             mat_A[437] * mat_B[677] +
//             mat_A[438] * mat_B[709] +
//             mat_A[439] * mat_B[741] +
//             mat_A[440] * mat_B[773] +
//             mat_A[441] * mat_B[805] +
//             mat_A[442] * mat_B[837] +
//             mat_A[443] * mat_B[869] +
//             mat_A[444] * mat_B[901] +
//             mat_A[445] * mat_B[933] +
//             mat_A[446] * mat_B[965] +
//             mat_A[447] * mat_B[997];
//  mat_C[422] <= 
//             mat_A[416] * mat_B[6] +
//             mat_A[417] * mat_B[38] +
//             mat_A[418] * mat_B[70] +
//             mat_A[419] * mat_B[102] +
//             mat_A[420] * mat_B[134] +
//             mat_A[421] * mat_B[166] +
//             mat_A[422] * mat_B[198] +
//             mat_A[423] * mat_B[230] +
//             mat_A[424] * mat_B[262] +
//             mat_A[425] * mat_B[294] +
//             mat_A[426] * mat_B[326] +
//             mat_A[427] * mat_B[358] +
//             mat_A[428] * mat_B[390] +
//             mat_A[429] * mat_B[422] +
//             mat_A[430] * mat_B[454] +
//             mat_A[431] * mat_B[486] +
//             mat_A[432] * mat_B[518] +
//             mat_A[433] * mat_B[550] +
//             mat_A[434] * mat_B[582] +
//             mat_A[435] * mat_B[614] +
//             mat_A[436] * mat_B[646] +
//             mat_A[437] * mat_B[678] +
//             mat_A[438] * mat_B[710] +
//             mat_A[439] * mat_B[742] +
//             mat_A[440] * mat_B[774] +
//             mat_A[441] * mat_B[806] +
//             mat_A[442] * mat_B[838] +
//             mat_A[443] * mat_B[870] +
//             mat_A[444] * mat_B[902] +
//             mat_A[445] * mat_B[934] +
//             mat_A[446] * mat_B[966] +
//             mat_A[447] * mat_B[998];
//  mat_C[423] <= 
//             mat_A[416] * mat_B[7] +
//             mat_A[417] * mat_B[39] +
//             mat_A[418] * mat_B[71] +
//             mat_A[419] * mat_B[103] +
//             mat_A[420] * mat_B[135] +
//             mat_A[421] * mat_B[167] +
//             mat_A[422] * mat_B[199] +
//             mat_A[423] * mat_B[231] +
//             mat_A[424] * mat_B[263] +
//             mat_A[425] * mat_B[295] +
//             mat_A[426] * mat_B[327] +
//             mat_A[427] * mat_B[359] +
//             mat_A[428] * mat_B[391] +
//             mat_A[429] * mat_B[423] +
//             mat_A[430] * mat_B[455] +
//             mat_A[431] * mat_B[487] +
//             mat_A[432] * mat_B[519] +
//             mat_A[433] * mat_B[551] +
//             mat_A[434] * mat_B[583] +
//             mat_A[435] * mat_B[615] +
//             mat_A[436] * mat_B[647] +
//             mat_A[437] * mat_B[679] +
//             mat_A[438] * mat_B[711] +
//             mat_A[439] * mat_B[743] +
//             mat_A[440] * mat_B[775] +
//             mat_A[441] * mat_B[807] +
//             mat_A[442] * mat_B[839] +
//             mat_A[443] * mat_B[871] +
//             mat_A[444] * mat_B[903] +
//             mat_A[445] * mat_B[935] +
//             mat_A[446] * mat_B[967] +
//             mat_A[447] * mat_B[999];
//  mat_C[424] <= 
//             mat_A[416] * mat_B[8] +
//             mat_A[417] * mat_B[40] +
//             mat_A[418] * mat_B[72] +
//             mat_A[419] * mat_B[104] +
//             mat_A[420] * mat_B[136] +
//             mat_A[421] * mat_B[168] +
//             mat_A[422] * mat_B[200] +
//             mat_A[423] * mat_B[232] +
//             mat_A[424] * mat_B[264] +
//             mat_A[425] * mat_B[296] +
//             mat_A[426] * mat_B[328] +
//             mat_A[427] * mat_B[360] +
//             mat_A[428] * mat_B[392] +
//             mat_A[429] * mat_B[424] +
//             mat_A[430] * mat_B[456] +
//             mat_A[431] * mat_B[488] +
//             mat_A[432] * mat_B[520] +
//             mat_A[433] * mat_B[552] +
//             mat_A[434] * mat_B[584] +
//             mat_A[435] * mat_B[616] +
//             mat_A[436] * mat_B[648] +
//             mat_A[437] * mat_B[680] +
//             mat_A[438] * mat_B[712] +
//             mat_A[439] * mat_B[744] +
//             mat_A[440] * mat_B[776] +
//             mat_A[441] * mat_B[808] +
//             mat_A[442] * mat_B[840] +
//             mat_A[443] * mat_B[872] +
//             mat_A[444] * mat_B[904] +
//             mat_A[445] * mat_B[936] +
//             mat_A[446] * mat_B[968] +
//             mat_A[447] * mat_B[1000];
//  mat_C[425] <= 
//             mat_A[416] * mat_B[9] +
//             mat_A[417] * mat_B[41] +
//             mat_A[418] * mat_B[73] +
//             mat_A[419] * mat_B[105] +
//             mat_A[420] * mat_B[137] +
//             mat_A[421] * mat_B[169] +
//             mat_A[422] * mat_B[201] +
//             mat_A[423] * mat_B[233] +
//             mat_A[424] * mat_B[265] +
//             mat_A[425] * mat_B[297] +
//             mat_A[426] * mat_B[329] +
//             mat_A[427] * mat_B[361] +
//             mat_A[428] * mat_B[393] +
//             mat_A[429] * mat_B[425] +
//             mat_A[430] * mat_B[457] +
//             mat_A[431] * mat_B[489] +
//             mat_A[432] * mat_B[521] +
//             mat_A[433] * mat_B[553] +
//             mat_A[434] * mat_B[585] +
//             mat_A[435] * mat_B[617] +
//             mat_A[436] * mat_B[649] +
//             mat_A[437] * mat_B[681] +
//             mat_A[438] * mat_B[713] +
//             mat_A[439] * mat_B[745] +
//             mat_A[440] * mat_B[777] +
//             mat_A[441] * mat_B[809] +
//             mat_A[442] * mat_B[841] +
//             mat_A[443] * mat_B[873] +
//             mat_A[444] * mat_B[905] +
//             mat_A[445] * mat_B[937] +
//             mat_A[446] * mat_B[969] +
//             mat_A[447] * mat_B[1001];
//  mat_C[426] <= 
//             mat_A[416] * mat_B[10] +
//             mat_A[417] * mat_B[42] +
//             mat_A[418] * mat_B[74] +
//             mat_A[419] * mat_B[106] +
//             mat_A[420] * mat_B[138] +
//             mat_A[421] * mat_B[170] +
//             mat_A[422] * mat_B[202] +
//             mat_A[423] * mat_B[234] +
//             mat_A[424] * mat_B[266] +
//             mat_A[425] * mat_B[298] +
//             mat_A[426] * mat_B[330] +
//             mat_A[427] * mat_B[362] +
//             mat_A[428] * mat_B[394] +
//             mat_A[429] * mat_B[426] +
//             mat_A[430] * mat_B[458] +
//             mat_A[431] * mat_B[490] +
//             mat_A[432] * mat_B[522] +
//             mat_A[433] * mat_B[554] +
//             mat_A[434] * mat_B[586] +
//             mat_A[435] * mat_B[618] +
//             mat_A[436] * mat_B[650] +
//             mat_A[437] * mat_B[682] +
//             mat_A[438] * mat_B[714] +
//             mat_A[439] * mat_B[746] +
//             mat_A[440] * mat_B[778] +
//             mat_A[441] * mat_B[810] +
//             mat_A[442] * mat_B[842] +
//             mat_A[443] * mat_B[874] +
//             mat_A[444] * mat_B[906] +
//             mat_A[445] * mat_B[938] +
//             mat_A[446] * mat_B[970] +
//             mat_A[447] * mat_B[1002];
//  mat_C[427] <= 
//             mat_A[416] * mat_B[11] +
//             mat_A[417] * mat_B[43] +
//             mat_A[418] * mat_B[75] +
//             mat_A[419] * mat_B[107] +
//             mat_A[420] * mat_B[139] +
//             mat_A[421] * mat_B[171] +
//             mat_A[422] * mat_B[203] +
//             mat_A[423] * mat_B[235] +
//             mat_A[424] * mat_B[267] +
//             mat_A[425] * mat_B[299] +
//             mat_A[426] * mat_B[331] +
//             mat_A[427] * mat_B[363] +
//             mat_A[428] * mat_B[395] +
//             mat_A[429] * mat_B[427] +
//             mat_A[430] * mat_B[459] +
//             mat_A[431] * mat_B[491] +
//             mat_A[432] * mat_B[523] +
//             mat_A[433] * mat_B[555] +
//             mat_A[434] * mat_B[587] +
//             mat_A[435] * mat_B[619] +
//             mat_A[436] * mat_B[651] +
//             mat_A[437] * mat_B[683] +
//             mat_A[438] * mat_B[715] +
//             mat_A[439] * mat_B[747] +
//             mat_A[440] * mat_B[779] +
//             mat_A[441] * mat_B[811] +
//             mat_A[442] * mat_B[843] +
//             mat_A[443] * mat_B[875] +
//             mat_A[444] * mat_B[907] +
//             mat_A[445] * mat_B[939] +
//             mat_A[446] * mat_B[971] +
//             mat_A[447] * mat_B[1003];
//  mat_C[428] <= 
//             mat_A[416] * mat_B[12] +
//             mat_A[417] * mat_B[44] +
//             mat_A[418] * mat_B[76] +
//             mat_A[419] * mat_B[108] +
//             mat_A[420] * mat_B[140] +
//             mat_A[421] * mat_B[172] +
//             mat_A[422] * mat_B[204] +
//             mat_A[423] * mat_B[236] +
//             mat_A[424] * mat_B[268] +
//             mat_A[425] * mat_B[300] +
//             mat_A[426] * mat_B[332] +
//             mat_A[427] * mat_B[364] +
//             mat_A[428] * mat_B[396] +
//             mat_A[429] * mat_B[428] +
//             mat_A[430] * mat_B[460] +
//             mat_A[431] * mat_B[492] +
//             mat_A[432] * mat_B[524] +
//             mat_A[433] * mat_B[556] +
//             mat_A[434] * mat_B[588] +
//             mat_A[435] * mat_B[620] +
//             mat_A[436] * mat_B[652] +
//             mat_A[437] * mat_B[684] +
//             mat_A[438] * mat_B[716] +
//             mat_A[439] * mat_B[748] +
//             mat_A[440] * mat_B[780] +
//             mat_A[441] * mat_B[812] +
//             mat_A[442] * mat_B[844] +
//             mat_A[443] * mat_B[876] +
//             mat_A[444] * mat_B[908] +
//             mat_A[445] * mat_B[940] +
//             mat_A[446] * mat_B[972] +
//             mat_A[447] * mat_B[1004];
//  mat_C[429] <= 
//             mat_A[416] * mat_B[13] +
//             mat_A[417] * mat_B[45] +
//             mat_A[418] * mat_B[77] +
//             mat_A[419] * mat_B[109] +
//             mat_A[420] * mat_B[141] +
//             mat_A[421] * mat_B[173] +
//             mat_A[422] * mat_B[205] +
//             mat_A[423] * mat_B[237] +
//             mat_A[424] * mat_B[269] +
//             mat_A[425] * mat_B[301] +
//             mat_A[426] * mat_B[333] +
//             mat_A[427] * mat_B[365] +
//             mat_A[428] * mat_B[397] +
//             mat_A[429] * mat_B[429] +
//             mat_A[430] * mat_B[461] +
//             mat_A[431] * mat_B[493] +
//             mat_A[432] * mat_B[525] +
//             mat_A[433] * mat_B[557] +
//             mat_A[434] * mat_B[589] +
//             mat_A[435] * mat_B[621] +
//             mat_A[436] * mat_B[653] +
//             mat_A[437] * mat_B[685] +
//             mat_A[438] * mat_B[717] +
//             mat_A[439] * mat_B[749] +
//             mat_A[440] * mat_B[781] +
//             mat_A[441] * mat_B[813] +
//             mat_A[442] * mat_B[845] +
//             mat_A[443] * mat_B[877] +
//             mat_A[444] * mat_B[909] +
//             mat_A[445] * mat_B[941] +
//             mat_A[446] * mat_B[973] +
//             mat_A[447] * mat_B[1005];
//  mat_C[430] <= 
//             mat_A[416] * mat_B[14] +
//             mat_A[417] * mat_B[46] +
//             mat_A[418] * mat_B[78] +
//             mat_A[419] * mat_B[110] +
//             mat_A[420] * mat_B[142] +
//             mat_A[421] * mat_B[174] +
//             mat_A[422] * mat_B[206] +
//             mat_A[423] * mat_B[238] +
//             mat_A[424] * mat_B[270] +
//             mat_A[425] * mat_B[302] +
//             mat_A[426] * mat_B[334] +
//             mat_A[427] * mat_B[366] +
//             mat_A[428] * mat_B[398] +
//             mat_A[429] * mat_B[430] +
//             mat_A[430] * mat_B[462] +
//             mat_A[431] * mat_B[494] +
//             mat_A[432] * mat_B[526] +
//             mat_A[433] * mat_B[558] +
//             mat_A[434] * mat_B[590] +
//             mat_A[435] * mat_B[622] +
//             mat_A[436] * mat_B[654] +
//             mat_A[437] * mat_B[686] +
//             mat_A[438] * mat_B[718] +
//             mat_A[439] * mat_B[750] +
//             mat_A[440] * mat_B[782] +
//             mat_A[441] * mat_B[814] +
//             mat_A[442] * mat_B[846] +
//             mat_A[443] * mat_B[878] +
//             mat_A[444] * mat_B[910] +
//             mat_A[445] * mat_B[942] +
//             mat_A[446] * mat_B[974] +
//             mat_A[447] * mat_B[1006];
//  mat_C[431] <= 
//             mat_A[416] * mat_B[15] +
//             mat_A[417] * mat_B[47] +
//             mat_A[418] * mat_B[79] +
//             mat_A[419] * mat_B[111] +
//             mat_A[420] * mat_B[143] +
//             mat_A[421] * mat_B[175] +
//             mat_A[422] * mat_B[207] +
//             mat_A[423] * mat_B[239] +
//             mat_A[424] * mat_B[271] +
//             mat_A[425] * mat_B[303] +
//             mat_A[426] * mat_B[335] +
//             mat_A[427] * mat_B[367] +
//             mat_A[428] * mat_B[399] +
//             mat_A[429] * mat_B[431] +
//             mat_A[430] * mat_B[463] +
//             mat_A[431] * mat_B[495] +
//             mat_A[432] * mat_B[527] +
//             mat_A[433] * mat_B[559] +
//             mat_A[434] * mat_B[591] +
//             mat_A[435] * mat_B[623] +
//             mat_A[436] * mat_B[655] +
//             mat_A[437] * mat_B[687] +
//             mat_A[438] * mat_B[719] +
//             mat_A[439] * mat_B[751] +
//             mat_A[440] * mat_B[783] +
//             mat_A[441] * mat_B[815] +
//             mat_A[442] * mat_B[847] +
//             mat_A[443] * mat_B[879] +
//             mat_A[444] * mat_B[911] +
//             mat_A[445] * mat_B[943] +
//             mat_A[446] * mat_B[975] +
//             mat_A[447] * mat_B[1007];
//  mat_C[432] <= 
//             mat_A[416] * mat_B[16] +
//             mat_A[417] * mat_B[48] +
//             mat_A[418] * mat_B[80] +
//             mat_A[419] * mat_B[112] +
//             mat_A[420] * mat_B[144] +
//             mat_A[421] * mat_B[176] +
//             mat_A[422] * mat_B[208] +
//             mat_A[423] * mat_B[240] +
//             mat_A[424] * mat_B[272] +
//             mat_A[425] * mat_B[304] +
//             mat_A[426] * mat_B[336] +
//             mat_A[427] * mat_B[368] +
//             mat_A[428] * mat_B[400] +
//             mat_A[429] * mat_B[432] +
//             mat_A[430] * mat_B[464] +
//             mat_A[431] * mat_B[496] +
//             mat_A[432] * mat_B[528] +
//             mat_A[433] * mat_B[560] +
//             mat_A[434] * mat_B[592] +
//             mat_A[435] * mat_B[624] +
//             mat_A[436] * mat_B[656] +
//             mat_A[437] * mat_B[688] +
//             mat_A[438] * mat_B[720] +
//             mat_A[439] * mat_B[752] +
//             mat_A[440] * mat_B[784] +
//             mat_A[441] * mat_B[816] +
//             mat_A[442] * mat_B[848] +
//             mat_A[443] * mat_B[880] +
//             mat_A[444] * mat_B[912] +
//             mat_A[445] * mat_B[944] +
//             mat_A[446] * mat_B[976] +
//             mat_A[447] * mat_B[1008];
//  mat_C[433] <= 
//             mat_A[416] * mat_B[17] +
//             mat_A[417] * mat_B[49] +
//             mat_A[418] * mat_B[81] +
//             mat_A[419] * mat_B[113] +
//             mat_A[420] * mat_B[145] +
//             mat_A[421] * mat_B[177] +
//             mat_A[422] * mat_B[209] +
//             mat_A[423] * mat_B[241] +
//             mat_A[424] * mat_B[273] +
//             mat_A[425] * mat_B[305] +
//             mat_A[426] * mat_B[337] +
//             mat_A[427] * mat_B[369] +
//             mat_A[428] * mat_B[401] +
//             mat_A[429] * mat_B[433] +
//             mat_A[430] * mat_B[465] +
//             mat_A[431] * mat_B[497] +
//             mat_A[432] * mat_B[529] +
//             mat_A[433] * mat_B[561] +
//             mat_A[434] * mat_B[593] +
//             mat_A[435] * mat_B[625] +
//             mat_A[436] * mat_B[657] +
//             mat_A[437] * mat_B[689] +
//             mat_A[438] * mat_B[721] +
//             mat_A[439] * mat_B[753] +
//             mat_A[440] * mat_B[785] +
//             mat_A[441] * mat_B[817] +
//             mat_A[442] * mat_B[849] +
//             mat_A[443] * mat_B[881] +
//             mat_A[444] * mat_B[913] +
//             mat_A[445] * mat_B[945] +
//             mat_A[446] * mat_B[977] +
//             mat_A[447] * mat_B[1009];
//  mat_C[434] <= 
//             mat_A[416] * mat_B[18] +
//             mat_A[417] * mat_B[50] +
//             mat_A[418] * mat_B[82] +
//             mat_A[419] * mat_B[114] +
//             mat_A[420] * mat_B[146] +
//             mat_A[421] * mat_B[178] +
//             mat_A[422] * mat_B[210] +
//             mat_A[423] * mat_B[242] +
//             mat_A[424] * mat_B[274] +
//             mat_A[425] * mat_B[306] +
//             mat_A[426] * mat_B[338] +
//             mat_A[427] * mat_B[370] +
//             mat_A[428] * mat_B[402] +
//             mat_A[429] * mat_B[434] +
//             mat_A[430] * mat_B[466] +
//             mat_A[431] * mat_B[498] +
//             mat_A[432] * mat_B[530] +
//             mat_A[433] * mat_B[562] +
//             mat_A[434] * mat_B[594] +
//             mat_A[435] * mat_B[626] +
//             mat_A[436] * mat_B[658] +
//             mat_A[437] * mat_B[690] +
//             mat_A[438] * mat_B[722] +
//             mat_A[439] * mat_B[754] +
//             mat_A[440] * mat_B[786] +
//             mat_A[441] * mat_B[818] +
//             mat_A[442] * mat_B[850] +
//             mat_A[443] * mat_B[882] +
//             mat_A[444] * mat_B[914] +
//             mat_A[445] * mat_B[946] +
//             mat_A[446] * mat_B[978] +
//             mat_A[447] * mat_B[1010];
//  mat_C[435] <= 
//             mat_A[416] * mat_B[19] +
//             mat_A[417] * mat_B[51] +
//             mat_A[418] * mat_B[83] +
//             mat_A[419] * mat_B[115] +
//             mat_A[420] * mat_B[147] +
//             mat_A[421] * mat_B[179] +
//             mat_A[422] * mat_B[211] +
//             mat_A[423] * mat_B[243] +
//             mat_A[424] * mat_B[275] +
//             mat_A[425] * mat_B[307] +
//             mat_A[426] * mat_B[339] +
//             mat_A[427] * mat_B[371] +
//             mat_A[428] * mat_B[403] +
//             mat_A[429] * mat_B[435] +
//             mat_A[430] * mat_B[467] +
//             mat_A[431] * mat_B[499] +
//             mat_A[432] * mat_B[531] +
//             mat_A[433] * mat_B[563] +
//             mat_A[434] * mat_B[595] +
//             mat_A[435] * mat_B[627] +
//             mat_A[436] * mat_B[659] +
//             mat_A[437] * mat_B[691] +
//             mat_A[438] * mat_B[723] +
//             mat_A[439] * mat_B[755] +
//             mat_A[440] * mat_B[787] +
//             mat_A[441] * mat_B[819] +
//             mat_A[442] * mat_B[851] +
//             mat_A[443] * mat_B[883] +
//             mat_A[444] * mat_B[915] +
//             mat_A[445] * mat_B[947] +
//             mat_A[446] * mat_B[979] +
//             mat_A[447] * mat_B[1011];
//  mat_C[436] <= 
//             mat_A[416] * mat_B[20] +
//             mat_A[417] * mat_B[52] +
//             mat_A[418] * mat_B[84] +
//             mat_A[419] * mat_B[116] +
//             mat_A[420] * mat_B[148] +
//             mat_A[421] * mat_B[180] +
//             mat_A[422] * mat_B[212] +
//             mat_A[423] * mat_B[244] +
//             mat_A[424] * mat_B[276] +
//             mat_A[425] * mat_B[308] +
//             mat_A[426] * mat_B[340] +
//             mat_A[427] * mat_B[372] +
//             mat_A[428] * mat_B[404] +
//             mat_A[429] * mat_B[436] +
//             mat_A[430] * mat_B[468] +
//             mat_A[431] * mat_B[500] +
//             mat_A[432] * mat_B[532] +
//             mat_A[433] * mat_B[564] +
//             mat_A[434] * mat_B[596] +
//             mat_A[435] * mat_B[628] +
//             mat_A[436] * mat_B[660] +
//             mat_A[437] * mat_B[692] +
//             mat_A[438] * mat_B[724] +
//             mat_A[439] * mat_B[756] +
//             mat_A[440] * mat_B[788] +
//             mat_A[441] * mat_B[820] +
//             mat_A[442] * mat_B[852] +
//             mat_A[443] * mat_B[884] +
//             mat_A[444] * mat_B[916] +
//             mat_A[445] * mat_B[948] +
//             mat_A[446] * mat_B[980] +
//             mat_A[447] * mat_B[1012];
//  mat_C[437] <= 
//             mat_A[416] * mat_B[21] +
//             mat_A[417] * mat_B[53] +
//             mat_A[418] * mat_B[85] +
//             mat_A[419] * mat_B[117] +
//             mat_A[420] * mat_B[149] +
//             mat_A[421] * mat_B[181] +
//             mat_A[422] * mat_B[213] +
//             mat_A[423] * mat_B[245] +
//             mat_A[424] * mat_B[277] +
//             mat_A[425] * mat_B[309] +
//             mat_A[426] * mat_B[341] +
//             mat_A[427] * mat_B[373] +
//             mat_A[428] * mat_B[405] +
//             mat_A[429] * mat_B[437] +
//             mat_A[430] * mat_B[469] +
//             mat_A[431] * mat_B[501] +
//             mat_A[432] * mat_B[533] +
//             mat_A[433] * mat_B[565] +
//             mat_A[434] * mat_B[597] +
//             mat_A[435] * mat_B[629] +
//             mat_A[436] * mat_B[661] +
//             mat_A[437] * mat_B[693] +
//             mat_A[438] * mat_B[725] +
//             mat_A[439] * mat_B[757] +
//             mat_A[440] * mat_B[789] +
//             mat_A[441] * mat_B[821] +
//             mat_A[442] * mat_B[853] +
//             mat_A[443] * mat_B[885] +
//             mat_A[444] * mat_B[917] +
//             mat_A[445] * mat_B[949] +
//             mat_A[446] * mat_B[981] +
//             mat_A[447] * mat_B[1013];
//  mat_C[438] <= 
//             mat_A[416] * mat_B[22] +
//             mat_A[417] * mat_B[54] +
//             mat_A[418] * mat_B[86] +
//             mat_A[419] * mat_B[118] +
//             mat_A[420] * mat_B[150] +
//             mat_A[421] * mat_B[182] +
//             mat_A[422] * mat_B[214] +
//             mat_A[423] * mat_B[246] +
//             mat_A[424] * mat_B[278] +
//             mat_A[425] * mat_B[310] +
//             mat_A[426] * mat_B[342] +
//             mat_A[427] * mat_B[374] +
//             mat_A[428] * mat_B[406] +
//             mat_A[429] * mat_B[438] +
//             mat_A[430] * mat_B[470] +
//             mat_A[431] * mat_B[502] +
//             mat_A[432] * mat_B[534] +
//             mat_A[433] * mat_B[566] +
//             mat_A[434] * mat_B[598] +
//             mat_A[435] * mat_B[630] +
//             mat_A[436] * mat_B[662] +
//             mat_A[437] * mat_B[694] +
//             mat_A[438] * mat_B[726] +
//             mat_A[439] * mat_B[758] +
//             mat_A[440] * mat_B[790] +
//             mat_A[441] * mat_B[822] +
//             mat_A[442] * mat_B[854] +
//             mat_A[443] * mat_B[886] +
//             mat_A[444] * mat_B[918] +
//             mat_A[445] * mat_B[950] +
//             mat_A[446] * mat_B[982] +
//             mat_A[447] * mat_B[1014];
//  mat_C[439] <= 
//             mat_A[416] * mat_B[23] +
//             mat_A[417] * mat_B[55] +
//             mat_A[418] * mat_B[87] +
//             mat_A[419] * mat_B[119] +
//             mat_A[420] * mat_B[151] +
//             mat_A[421] * mat_B[183] +
//             mat_A[422] * mat_B[215] +
//             mat_A[423] * mat_B[247] +
//             mat_A[424] * mat_B[279] +
//             mat_A[425] * mat_B[311] +
//             mat_A[426] * mat_B[343] +
//             mat_A[427] * mat_B[375] +
//             mat_A[428] * mat_B[407] +
//             mat_A[429] * mat_B[439] +
//             mat_A[430] * mat_B[471] +
//             mat_A[431] * mat_B[503] +
//             mat_A[432] * mat_B[535] +
//             mat_A[433] * mat_B[567] +
//             mat_A[434] * mat_B[599] +
//             mat_A[435] * mat_B[631] +
//             mat_A[436] * mat_B[663] +
//             mat_A[437] * mat_B[695] +
//             mat_A[438] * mat_B[727] +
//             mat_A[439] * mat_B[759] +
//             mat_A[440] * mat_B[791] +
//             mat_A[441] * mat_B[823] +
//             mat_A[442] * mat_B[855] +
//             mat_A[443] * mat_B[887] +
//             mat_A[444] * mat_B[919] +
//             mat_A[445] * mat_B[951] +
//             mat_A[446] * mat_B[983] +
//             mat_A[447] * mat_B[1015];
//  mat_C[440] <= 
//             mat_A[416] * mat_B[24] +
//             mat_A[417] * mat_B[56] +
//             mat_A[418] * mat_B[88] +
//             mat_A[419] * mat_B[120] +
//             mat_A[420] * mat_B[152] +
//             mat_A[421] * mat_B[184] +
//             mat_A[422] * mat_B[216] +
//             mat_A[423] * mat_B[248] +
//             mat_A[424] * mat_B[280] +
//             mat_A[425] * mat_B[312] +
//             mat_A[426] * mat_B[344] +
//             mat_A[427] * mat_B[376] +
//             mat_A[428] * mat_B[408] +
//             mat_A[429] * mat_B[440] +
//             mat_A[430] * mat_B[472] +
//             mat_A[431] * mat_B[504] +
//             mat_A[432] * mat_B[536] +
//             mat_A[433] * mat_B[568] +
//             mat_A[434] * mat_B[600] +
//             mat_A[435] * mat_B[632] +
//             mat_A[436] * mat_B[664] +
//             mat_A[437] * mat_B[696] +
//             mat_A[438] * mat_B[728] +
//             mat_A[439] * mat_B[760] +
//             mat_A[440] * mat_B[792] +
//             mat_A[441] * mat_B[824] +
//             mat_A[442] * mat_B[856] +
//             mat_A[443] * mat_B[888] +
//             mat_A[444] * mat_B[920] +
//             mat_A[445] * mat_B[952] +
//             mat_A[446] * mat_B[984] +
//             mat_A[447] * mat_B[1016];
//  mat_C[441] <= 
//             mat_A[416] * mat_B[25] +
//             mat_A[417] * mat_B[57] +
//             mat_A[418] * mat_B[89] +
//             mat_A[419] * mat_B[121] +
//             mat_A[420] * mat_B[153] +
//             mat_A[421] * mat_B[185] +
//             mat_A[422] * mat_B[217] +
//             mat_A[423] * mat_B[249] +
//             mat_A[424] * mat_B[281] +
//             mat_A[425] * mat_B[313] +
//             mat_A[426] * mat_B[345] +
//             mat_A[427] * mat_B[377] +
//             mat_A[428] * mat_B[409] +
//             mat_A[429] * mat_B[441] +
//             mat_A[430] * mat_B[473] +
//             mat_A[431] * mat_B[505] +
//             mat_A[432] * mat_B[537] +
//             mat_A[433] * mat_B[569] +
//             mat_A[434] * mat_B[601] +
//             mat_A[435] * mat_B[633] +
//             mat_A[436] * mat_B[665] +
//             mat_A[437] * mat_B[697] +
//             mat_A[438] * mat_B[729] +
//             mat_A[439] * mat_B[761] +
//             mat_A[440] * mat_B[793] +
//             mat_A[441] * mat_B[825] +
//             mat_A[442] * mat_B[857] +
//             mat_A[443] * mat_B[889] +
//             mat_A[444] * mat_B[921] +
//             mat_A[445] * mat_B[953] +
//             mat_A[446] * mat_B[985] +
//             mat_A[447] * mat_B[1017];
//  mat_C[442] <= 
//             mat_A[416] * mat_B[26] +
//             mat_A[417] * mat_B[58] +
//             mat_A[418] * mat_B[90] +
//             mat_A[419] * mat_B[122] +
//             mat_A[420] * mat_B[154] +
//             mat_A[421] * mat_B[186] +
//             mat_A[422] * mat_B[218] +
//             mat_A[423] * mat_B[250] +
//             mat_A[424] * mat_B[282] +
//             mat_A[425] * mat_B[314] +
//             mat_A[426] * mat_B[346] +
//             mat_A[427] * mat_B[378] +
//             mat_A[428] * mat_B[410] +
//             mat_A[429] * mat_B[442] +
//             mat_A[430] * mat_B[474] +
//             mat_A[431] * mat_B[506] +
//             mat_A[432] * mat_B[538] +
//             mat_A[433] * mat_B[570] +
//             mat_A[434] * mat_B[602] +
//             mat_A[435] * mat_B[634] +
//             mat_A[436] * mat_B[666] +
//             mat_A[437] * mat_B[698] +
//             mat_A[438] * mat_B[730] +
//             mat_A[439] * mat_B[762] +
//             mat_A[440] * mat_B[794] +
//             mat_A[441] * mat_B[826] +
//             mat_A[442] * mat_B[858] +
//             mat_A[443] * mat_B[890] +
//             mat_A[444] * mat_B[922] +
//             mat_A[445] * mat_B[954] +
//             mat_A[446] * mat_B[986] +
//             mat_A[447] * mat_B[1018];
//  mat_C[443] <= 
//             mat_A[416] * mat_B[27] +
//             mat_A[417] * mat_B[59] +
//             mat_A[418] * mat_B[91] +
//             mat_A[419] * mat_B[123] +
//             mat_A[420] * mat_B[155] +
//             mat_A[421] * mat_B[187] +
//             mat_A[422] * mat_B[219] +
//             mat_A[423] * mat_B[251] +
//             mat_A[424] * mat_B[283] +
//             mat_A[425] * mat_B[315] +
//             mat_A[426] * mat_B[347] +
//             mat_A[427] * mat_B[379] +
//             mat_A[428] * mat_B[411] +
//             mat_A[429] * mat_B[443] +
//             mat_A[430] * mat_B[475] +
//             mat_A[431] * mat_B[507] +
//             mat_A[432] * mat_B[539] +
//             mat_A[433] * mat_B[571] +
//             mat_A[434] * mat_B[603] +
//             mat_A[435] * mat_B[635] +
//             mat_A[436] * mat_B[667] +
//             mat_A[437] * mat_B[699] +
//             mat_A[438] * mat_B[731] +
//             mat_A[439] * mat_B[763] +
//             mat_A[440] * mat_B[795] +
//             mat_A[441] * mat_B[827] +
//             mat_A[442] * mat_B[859] +
//             mat_A[443] * mat_B[891] +
//             mat_A[444] * mat_B[923] +
//             mat_A[445] * mat_B[955] +
//             mat_A[446] * mat_B[987] +
//             mat_A[447] * mat_B[1019];
//  mat_C[444] <= 
//             mat_A[416] * mat_B[28] +
//             mat_A[417] * mat_B[60] +
//             mat_A[418] * mat_B[92] +
//             mat_A[419] * mat_B[124] +
//             mat_A[420] * mat_B[156] +
//             mat_A[421] * mat_B[188] +
//             mat_A[422] * mat_B[220] +
//             mat_A[423] * mat_B[252] +
//             mat_A[424] * mat_B[284] +
//             mat_A[425] * mat_B[316] +
//             mat_A[426] * mat_B[348] +
//             mat_A[427] * mat_B[380] +
//             mat_A[428] * mat_B[412] +
//             mat_A[429] * mat_B[444] +
//             mat_A[430] * mat_B[476] +
//             mat_A[431] * mat_B[508] +
//             mat_A[432] * mat_B[540] +
//             mat_A[433] * mat_B[572] +
//             mat_A[434] * mat_B[604] +
//             mat_A[435] * mat_B[636] +
//             mat_A[436] * mat_B[668] +
//             mat_A[437] * mat_B[700] +
//             mat_A[438] * mat_B[732] +
//             mat_A[439] * mat_B[764] +
//             mat_A[440] * mat_B[796] +
//             mat_A[441] * mat_B[828] +
//             mat_A[442] * mat_B[860] +
//             mat_A[443] * mat_B[892] +
//             mat_A[444] * mat_B[924] +
//             mat_A[445] * mat_B[956] +
//             mat_A[446] * mat_B[988] +
//             mat_A[447] * mat_B[1020];
//  mat_C[445] <= 
//             mat_A[416] * mat_B[29] +
//             mat_A[417] * mat_B[61] +
//             mat_A[418] * mat_B[93] +
//             mat_A[419] * mat_B[125] +
//             mat_A[420] * mat_B[157] +
//             mat_A[421] * mat_B[189] +
//             mat_A[422] * mat_B[221] +
//             mat_A[423] * mat_B[253] +
//             mat_A[424] * mat_B[285] +
//             mat_A[425] * mat_B[317] +
//             mat_A[426] * mat_B[349] +
//             mat_A[427] * mat_B[381] +
//             mat_A[428] * mat_B[413] +
//             mat_A[429] * mat_B[445] +
//             mat_A[430] * mat_B[477] +
//             mat_A[431] * mat_B[509] +
//             mat_A[432] * mat_B[541] +
//             mat_A[433] * mat_B[573] +
//             mat_A[434] * mat_B[605] +
//             mat_A[435] * mat_B[637] +
//             mat_A[436] * mat_B[669] +
//             mat_A[437] * mat_B[701] +
//             mat_A[438] * mat_B[733] +
//             mat_A[439] * mat_B[765] +
//             mat_A[440] * mat_B[797] +
//             mat_A[441] * mat_B[829] +
//             mat_A[442] * mat_B[861] +
//             mat_A[443] * mat_B[893] +
//             mat_A[444] * mat_B[925] +
//             mat_A[445] * mat_B[957] +
//             mat_A[446] * mat_B[989] +
//             mat_A[447] * mat_B[1021];
//  mat_C[446] <= 
//             mat_A[416] * mat_B[30] +
//             mat_A[417] * mat_B[62] +
//             mat_A[418] * mat_B[94] +
//             mat_A[419] * mat_B[126] +
//             mat_A[420] * mat_B[158] +
//             mat_A[421] * mat_B[190] +
//             mat_A[422] * mat_B[222] +
//             mat_A[423] * mat_B[254] +
//             mat_A[424] * mat_B[286] +
//             mat_A[425] * mat_B[318] +
//             mat_A[426] * mat_B[350] +
//             mat_A[427] * mat_B[382] +
//             mat_A[428] * mat_B[414] +
//             mat_A[429] * mat_B[446] +
//             mat_A[430] * mat_B[478] +
//             mat_A[431] * mat_B[510] +
//             mat_A[432] * mat_B[542] +
//             mat_A[433] * mat_B[574] +
//             mat_A[434] * mat_B[606] +
//             mat_A[435] * mat_B[638] +
//             mat_A[436] * mat_B[670] +
//             mat_A[437] * mat_B[702] +
//             mat_A[438] * mat_B[734] +
//             mat_A[439] * mat_B[766] +
//             mat_A[440] * mat_B[798] +
//             mat_A[441] * mat_B[830] +
//             mat_A[442] * mat_B[862] +
//             mat_A[443] * mat_B[894] +
//             mat_A[444] * mat_B[926] +
//             mat_A[445] * mat_B[958] +
//             mat_A[446] * mat_B[990] +
//             mat_A[447] * mat_B[1022];
//  mat_C[447] <= 
//             mat_A[416] * mat_B[31] +
//             mat_A[417] * mat_B[63] +
//             mat_A[418] * mat_B[95] +
//             mat_A[419] * mat_B[127] +
//             mat_A[420] * mat_B[159] +
//             mat_A[421] * mat_B[191] +
//             mat_A[422] * mat_B[223] +
//             mat_A[423] * mat_B[255] +
//             mat_A[424] * mat_B[287] +
//             mat_A[425] * mat_B[319] +
//             mat_A[426] * mat_B[351] +
//             mat_A[427] * mat_B[383] +
//             mat_A[428] * mat_B[415] +
//             mat_A[429] * mat_B[447] +
//             mat_A[430] * mat_B[479] +
//             mat_A[431] * mat_B[511] +
//             mat_A[432] * mat_B[543] +
//             mat_A[433] * mat_B[575] +
//             mat_A[434] * mat_B[607] +
//             mat_A[435] * mat_B[639] +
//             mat_A[436] * mat_B[671] +
//             mat_A[437] * mat_B[703] +
//             mat_A[438] * mat_B[735] +
//             mat_A[439] * mat_B[767] +
//             mat_A[440] * mat_B[799] +
//             mat_A[441] * mat_B[831] +
//             mat_A[442] * mat_B[863] +
//             mat_A[443] * mat_B[895] +
//             mat_A[444] * mat_B[927] +
//             mat_A[445] * mat_B[959] +
//             mat_A[446] * mat_B[991] +
//             mat_A[447] * mat_B[1023];
//  mat_C[448] <= 
//             mat_A[448] * mat_B[0] +
//             mat_A[449] * mat_B[32] +
//             mat_A[450] * mat_B[64] +
//             mat_A[451] * mat_B[96] +
//             mat_A[452] * mat_B[128] +
//             mat_A[453] * mat_B[160] +
//             mat_A[454] * mat_B[192] +
//             mat_A[455] * mat_B[224] +
//             mat_A[456] * mat_B[256] +
//             mat_A[457] * mat_B[288] +
//             mat_A[458] * mat_B[320] +
//             mat_A[459] * mat_B[352] +
//             mat_A[460] * mat_B[384] +
//             mat_A[461] * mat_B[416] +
//             mat_A[462] * mat_B[448] +
//             mat_A[463] * mat_B[480] +
//             mat_A[464] * mat_B[512] +
//             mat_A[465] * mat_B[544] +
//             mat_A[466] * mat_B[576] +
//             mat_A[467] * mat_B[608] +
//             mat_A[468] * mat_B[640] +
//             mat_A[469] * mat_B[672] +
//             mat_A[470] * mat_B[704] +
//             mat_A[471] * mat_B[736] +
//             mat_A[472] * mat_B[768] +
//             mat_A[473] * mat_B[800] +
//             mat_A[474] * mat_B[832] +
//             mat_A[475] * mat_B[864] +
//             mat_A[476] * mat_B[896] +
//             mat_A[477] * mat_B[928] +
//             mat_A[478] * mat_B[960] +
//             mat_A[479] * mat_B[992];
//  mat_C[449] <= 
//             mat_A[448] * mat_B[1] +
//             mat_A[449] * mat_B[33] +
//             mat_A[450] * mat_B[65] +
//             mat_A[451] * mat_B[97] +
//             mat_A[452] * mat_B[129] +
//             mat_A[453] * mat_B[161] +
//             mat_A[454] * mat_B[193] +
//             mat_A[455] * mat_B[225] +
//             mat_A[456] * mat_B[257] +
//             mat_A[457] * mat_B[289] +
//             mat_A[458] * mat_B[321] +
//             mat_A[459] * mat_B[353] +
//             mat_A[460] * mat_B[385] +
//             mat_A[461] * mat_B[417] +
//             mat_A[462] * mat_B[449] +
//             mat_A[463] * mat_B[481] +
//             mat_A[464] * mat_B[513] +
//             mat_A[465] * mat_B[545] +
//             mat_A[466] * mat_B[577] +
//             mat_A[467] * mat_B[609] +
//             mat_A[468] * mat_B[641] +
//             mat_A[469] * mat_B[673] +
//             mat_A[470] * mat_B[705] +
//             mat_A[471] * mat_B[737] +
//             mat_A[472] * mat_B[769] +
//             mat_A[473] * mat_B[801] +
//             mat_A[474] * mat_B[833] +
//             mat_A[475] * mat_B[865] +
//             mat_A[476] * mat_B[897] +
//             mat_A[477] * mat_B[929] +
//             mat_A[478] * mat_B[961] +
//             mat_A[479] * mat_B[993];
//  mat_C[450] <= 
//             mat_A[448] * mat_B[2] +
//             mat_A[449] * mat_B[34] +
//             mat_A[450] * mat_B[66] +
//             mat_A[451] * mat_B[98] +
//             mat_A[452] * mat_B[130] +
//             mat_A[453] * mat_B[162] +
//             mat_A[454] * mat_B[194] +
//             mat_A[455] * mat_B[226] +
//             mat_A[456] * mat_B[258] +
//             mat_A[457] * mat_B[290] +
//             mat_A[458] * mat_B[322] +
//             mat_A[459] * mat_B[354] +
//             mat_A[460] * mat_B[386] +
//             mat_A[461] * mat_B[418] +
//             mat_A[462] * mat_B[450] +
//             mat_A[463] * mat_B[482] +
//             mat_A[464] * mat_B[514] +
//             mat_A[465] * mat_B[546] +
//             mat_A[466] * mat_B[578] +
//             mat_A[467] * mat_B[610] +
//             mat_A[468] * mat_B[642] +
//             mat_A[469] * mat_B[674] +
//             mat_A[470] * mat_B[706] +
//             mat_A[471] * mat_B[738] +
//             mat_A[472] * mat_B[770] +
//             mat_A[473] * mat_B[802] +
//             mat_A[474] * mat_B[834] +
//             mat_A[475] * mat_B[866] +
//             mat_A[476] * mat_B[898] +
//             mat_A[477] * mat_B[930] +
//             mat_A[478] * mat_B[962] +
//             mat_A[479] * mat_B[994];
//  mat_C[451] <= 
//             mat_A[448] * mat_B[3] +
//             mat_A[449] * mat_B[35] +
//             mat_A[450] * mat_B[67] +
//             mat_A[451] * mat_B[99] +
//             mat_A[452] * mat_B[131] +
//             mat_A[453] * mat_B[163] +
//             mat_A[454] * mat_B[195] +
//             mat_A[455] * mat_B[227] +
//             mat_A[456] * mat_B[259] +
//             mat_A[457] * mat_B[291] +
//             mat_A[458] * mat_B[323] +
//             mat_A[459] * mat_B[355] +
//             mat_A[460] * mat_B[387] +
//             mat_A[461] * mat_B[419] +
//             mat_A[462] * mat_B[451] +
//             mat_A[463] * mat_B[483] +
//             mat_A[464] * mat_B[515] +
//             mat_A[465] * mat_B[547] +
//             mat_A[466] * mat_B[579] +
//             mat_A[467] * mat_B[611] +
//             mat_A[468] * mat_B[643] +
//             mat_A[469] * mat_B[675] +
//             mat_A[470] * mat_B[707] +
//             mat_A[471] * mat_B[739] +
//             mat_A[472] * mat_B[771] +
//             mat_A[473] * mat_B[803] +
//             mat_A[474] * mat_B[835] +
//             mat_A[475] * mat_B[867] +
//             mat_A[476] * mat_B[899] +
//             mat_A[477] * mat_B[931] +
//             mat_A[478] * mat_B[963] +
//             mat_A[479] * mat_B[995];
//  mat_C[452] <= 
//             mat_A[448] * mat_B[4] +
//             mat_A[449] * mat_B[36] +
//             mat_A[450] * mat_B[68] +
//             mat_A[451] * mat_B[100] +
//             mat_A[452] * mat_B[132] +
//             mat_A[453] * mat_B[164] +
//             mat_A[454] * mat_B[196] +
//             mat_A[455] * mat_B[228] +
//             mat_A[456] * mat_B[260] +
//             mat_A[457] * mat_B[292] +
//             mat_A[458] * mat_B[324] +
//             mat_A[459] * mat_B[356] +
//             mat_A[460] * mat_B[388] +
//             mat_A[461] * mat_B[420] +
//             mat_A[462] * mat_B[452] +
//             mat_A[463] * mat_B[484] +
//             mat_A[464] * mat_B[516] +
//             mat_A[465] * mat_B[548] +
//             mat_A[466] * mat_B[580] +
//             mat_A[467] * mat_B[612] +
//             mat_A[468] * mat_B[644] +
//             mat_A[469] * mat_B[676] +
//             mat_A[470] * mat_B[708] +
//             mat_A[471] * mat_B[740] +
//             mat_A[472] * mat_B[772] +
//             mat_A[473] * mat_B[804] +
//             mat_A[474] * mat_B[836] +
//             mat_A[475] * mat_B[868] +
//             mat_A[476] * mat_B[900] +
//             mat_A[477] * mat_B[932] +
//             mat_A[478] * mat_B[964] +
//             mat_A[479] * mat_B[996];
//  mat_C[453] <= 
//             mat_A[448] * mat_B[5] +
//             mat_A[449] * mat_B[37] +
//             mat_A[450] * mat_B[69] +
//             mat_A[451] * mat_B[101] +
//             mat_A[452] * mat_B[133] +
//             mat_A[453] * mat_B[165] +
//             mat_A[454] * mat_B[197] +
//             mat_A[455] * mat_B[229] +
//             mat_A[456] * mat_B[261] +
//             mat_A[457] * mat_B[293] +
//             mat_A[458] * mat_B[325] +
//             mat_A[459] * mat_B[357] +
//             mat_A[460] * mat_B[389] +
//             mat_A[461] * mat_B[421] +
//             mat_A[462] * mat_B[453] +
//             mat_A[463] * mat_B[485] +
//             mat_A[464] * mat_B[517] +
//             mat_A[465] * mat_B[549] +
//             mat_A[466] * mat_B[581] +
//             mat_A[467] * mat_B[613] +
//             mat_A[468] * mat_B[645] +
//             mat_A[469] * mat_B[677] +
//             mat_A[470] * mat_B[709] +
//             mat_A[471] * mat_B[741] +
//             mat_A[472] * mat_B[773] +
//             mat_A[473] * mat_B[805] +
//             mat_A[474] * mat_B[837] +
//             mat_A[475] * mat_B[869] +
//             mat_A[476] * mat_B[901] +
//             mat_A[477] * mat_B[933] +
//             mat_A[478] * mat_B[965] +
//             mat_A[479] * mat_B[997];
//  mat_C[454] <= 
//             mat_A[448] * mat_B[6] +
//             mat_A[449] * mat_B[38] +
//             mat_A[450] * mat_B[70] +
//             mat_A[451] * mat_B[102] +
//             mat_A[452] * mat_B[134] +
//             mat_A[453] * mat_B[166] +
//             mat_A[454] * mat_B[198] +
//             mat_A[455] * mat_B[230] +
//             mat_A[456] * mat_B[262] +
//             mat_A[457] * mat_B[294] +
//             mat_A[458] * mat_B[326] +
//             mat_A[459] * mat_B[358] +
//             mat_A[460] * mat_B[390] +
//             mat_A[461] * mat_B[422] +
//             mat_A[462] * mat_B[454] +
//             mat_A[463] * mat_B[486] +
//             mat_A[464] * mat_B[518] +
//             mat_A[465] * mat_B[550] +
//             mat_A[466] * mat_B[582] +
//             mat_A[467] * mat_B[614] +
//             mat_A[468] * mat_B[646] +
//             mat_A[469] * mat_B[678] +
//             mat_A[470] * mat_B[710] +
//             mat_A[471] * mat_B[742] +
//             mat_A[472] * mat_B[774] +
//             mat_A[473] * mat_B[806] +
//             mat_A[474] * mat_B[838] +
//             mat_A[475] * mat_B[870] +
//             mat_A[476] * mat_B[902] +
//             mat_A[477] * mat_B[934] +
//             mat_A[478] * mat_B[966] +
//             mat_A[479] * mat_B[998];
//  mat_C[455] <= 
//             mat_A[448] * mat_B[7] +
//             mat_A[449] * mat_B[39] +
//             mat_A[450] * mat_B[71] +
//             mat_A[451] * mat_B[103] +
//             mat_A[452] * mat_B[135] +
//             mat_A[453] * mat_B[167] +
//             mat_A[454] * mat_B[199] +
//             mat_A[455] * mat_B[231] +
//             mat_A[456] * mat_B[263] +
//             mat_A[457] * mat_B[295] +
//             mat_A[458] * mat_B[327] +
//             mat_A[459] * mat_B[359] +
//             mat_A[460] * mat_B[391] +
//             mat_A[461] * mat_B[423] +
//             mat_A[462] * mat_B[455] +
//             mat_A[463] * mat_B[487] +
//             mat_A[464] * mat_B[519] +
//             mat_A[465] * mat_B[551] +
//             mat_A[466] * mat_B[583] +
//             mat_A[467] * mat_B[615] +
//             mat_A[468] * mat_B[647] +
//             mat_A[469] * mat_B[679] +
//             mat_A[470] * mat_B[711] +
//             mat_A[471] * mat_B[743] +
//             mat_A[472] * mat_B[775] +
//             mat_A[473] * mat_B[807] +
//             mat_A[474] * mat_B[839] +
//             mat_A[475] * mat_B[871] +
//             mat_A[476] * mat_B[903] +
//             mat_A[477] * mat_B[935] +
//             mat_A[478] * mat_B[967] +
//             mat_A[479] * mat_B[999];
//  mat_C[456] <= 
//             mat_A[448] * mat_B[8] +
//             mat_A[449] * mat_B[40] +
//             mat_A[450] * mat_B[72] +
//             mat_A[451] * mat_B[104] +
//             mat_A[452] * mat_B[136] +
//             mat_A[453] * mat_B[168] +
//             mat_A[454] * mat_B[200] +
//             mat_A[455] * mat_B[232] +
//             mat_A[456] * mat_B[264] +
//             mat_A[457] * mat_B[296] +
//             mat_A[458] * mat_B[328] +
//             mat_A[459] * mat_B[360] +
//             mat_A[460] * mat_B[392] +
//             mat_A[461] * mat_B[424] +
//             mat_A[462] * mat_B[456] +
//             mat_A[463] * mat_B[488] +
//             mat_A[464] * mat_B[520] +
//             mat_A[465] * mat_B[552] +
//             mat_A[466] * mat_B[584] +
//             mat_A[467] * mat_B[616] +
//             mat_A[468] * mat_B[648] +
//             mat_A[469] * mat_B[680] +
//             mat_A[470] * mat_B[712] +
//             mat_A[471] * mat_B[744] +
//             mat_A[472] * mat_B[776] +
//             mat_A[473] * mat_B[808] +
//             mat_A[474] * mat_B[840] +
//             mat_A[475] * mat_B[872] +
//             mat_A[476] * mat_B[904] +
//             mat_A[477] * mat_B[936] +
//             mat_A[478] * mat_B[968] +
//             mat_A[479] * mat_B[1000];
//  mat_C[457] <= 
//             mat_A[448] * mat_B[9] +
//             mat_A[449] * mat_B[41] +
//             mat_A[450] * mat_B[73] +
//             mat_A[451] * mat_B[105] +
//             mat_A[452] * mat_B[137] +
//             mat_A[453] * mat_B[169] +
//             mat_A[454] * mat_B[201] +
//             mat_A[455] * mat_B[233] +
//             mat_A[456] * mat_B[265] +
//             mat_A[457] * mat_B[297] +
//             mat_A[458] * mat_B[329] +
//             mat_A[459] * mat_B[361] +
//             mat_A[460] * mat_B[393] +
//             mat_A[461] * mat_B[425] +
//             mat_A[462] * mat_B[457] +
//             mat_A[463] * mat_B[489] +
//             mat_A[464] * mat_B[521] +
//             mat_A[465] * mat_B[553] +
//             mat_A[466] * mat_B[585] +
//             mat_A[467] * mat_B[617] +
//             mat_A[468] * mat_B[649] +
//             mat_A[469] * mat_B[681] +
//             mat_A[470] * mat_B[713] +
//             mat_A[471] * mat_B[745] +
//             mat_A[472] * mat_B[777] +
//             mat_A[473] * mat_B[809] +
//             mat_A[474] * mat_B[841] +
//             mat_A[475] * mat_B[873] +
//             mat_A[476] * mat_B[905] +
//             mat_A[477] * mat_B[937] +
//             mat_A[478] * mat_B[969] +
//             mat_A[479] * mat_B[1001];
//  mat_C[458] <= 
//             mat_A[448] * mat_B[10] +
//             mat_A[449] * mat_B[42] +
//             mat_A[450] * mat_B[74] +
//             mat_A[451] * mat_B[106] +
//             mat_A[452] * mat_B[138] +
//             mat_A[453] * mat_B[170] +
//             mat_A[454] * mat_B[202] +
//             mat_A[455] * mat_B[234] +
//             mat_A[456] * mat_B[266] +
//             mat_A[457] * mat_B[298] +
//             mat_A[458] * mat_B[330] +
//             mat_A[459] * mat_B[362] +
//             mat_A[460] * mat_B[394] +
//             mat_A[461] * mat_B[426] +
//             mat_A[462] * mat_B[458] +
//             mat_A[463] * mat_B[490] +
//             mat_A[464] * mat_B[522] +
//             mat_A[465] * mat_B[554] +
//             mat_A[466] * mat_B[586] +
//             mat_A[467] * mat_B[618] +
//             mat_A[468] * mat_B[650] +
//             mat_A[469] * mat_B[682] +
//             mat_A[470] * mat_B[714] +
//             mat_A[471] * mat_B[746] +
//             mat_A[472] * mat_B[778] +
//             mat_A[473] * mat_B[810] +
//             mat_A[474] * mat_B[842] +
//             mat_A[475] * mat_B[874] +
//             mat_A[476] * mat_B[906] +
//             mat_A[477] * mat_B[938] +
//             mat_A[478] * mat_B[970] +
//             mat_A[479] * mat_B[1002];
//  mat_C[459] <= 
//             mat_A[448] * mat_B[11] +
//             mat_A[449] * mat_B[43] +
//             mat_A[450] * mat_B[75] +
//             mat_A[451] * mat_B[107] +
//             mat_A[452] * mat_B[139] +
//             mat_A[453] * mat_B[171] +
//             mat_A[454] * mat_B[203] +
//             mat_A[455] * mat_B[235] +
//             mat_A[456] * mat_B[267] +
//             mat_A[457] * mat_B[299] +
//             mat_A[458] * mat_B[331] +
//             mat_A[459] * mat_B[363] +
//             mat_A[460] * mat_B[395] +
//             mat_A[461] * mat_B[427] +
//             mat_A[462] * mat_B[459] +
//             mat_A[463] * mat_B[491] +
//             mat_A[464] * mat_B[523] +
//             mat_A[465] * mat_B[555] +
//             mat_A[466] * mat_B[587] +
//             mat_A[467] * mat_B[619] +
//             mat_A[468] * mat_B[651] +
//             mat_A[469] * mat_B[683] +
//             mat_A[470] * mat_B[715] +
//             mat_A[471] * mat_B[747] +
//             mat_A[472] * mat_B[779] +
//             mat_A[473] * mat_B[811] +
//             mat_A[474] * mat_B[843] +
//             mat_A[475] * mat_B[875] +
//             mat_A[476] * mat_B[907] +
//             mat_A[477] * mat_B[939] +
//             mat_A[478] * mat_B[971] +
//             mat_A[479] * mat_B[1003];
//  mat_C[460] <= 
//             mat_A[448] * mat_B[12] +
//             mat_A[449] * mat_B[44] +
//             mat_A[450] * mat_B[76] +
//             mat_A[451] * mat_B[108] +
//             mat_A[452] * mat_B[140] +
//             mat_A[453] * mat_B[172] +
//             mat_A[454] * mat_B[204] +
//             mat_A[455] * mat_B[236] +
//             mat_A[456] * mat_B[268] +
//             mat_A[457] * mat_B[300] +
//             mat_A[458] * mat_B[332] +
//             mat_A[459] * mat_B[364] +
//             mat_A[460] * mat_B[396] +
//             mat_A[461] * mat_B[428] +
//             mat_A[462] * mat_B[460] +
//             mat_A[463] * mat_B[492] +
//             mat_A[464] * mat_B[524] +
//             mat_A[465] * mat_B[556] +
//             mat_A[466] * mat_B[588] +
//             mat_A[467] * mat_B[620] +
//             mat_A[468] * mat_B[652] +
//             mat_A[469] * mat_B[684] +
//             mat_A[470] * mat_B[716] +
//             mat_A[471] * mat_B[748] +
//             mat_A[472] * mat_B[780] +
//             mat_A[473] * mat_B[812] +
//             mat_A[474] * mat_B[844] +
//             mat_A[475] * mat_B[876] +
//             mat_A[476] * mat_B[908] +
//             mat_A[477] * mat_B[940] +
//             mat_A[478] * mat_B[972] +
//             mat_A[479] * mat_B[1004];
//  mat_C[461] <= 
//             mat_A[448] * mat_B[13] +
//             mat_A[449] * mat_B[45] +
//             mat_A[450] * mat_B[77] +
//             mat_A[451] * mat_B[109] +
//             mat_A[452] * mat_B[141] +
//             mat_A[453] * mat_B[173] +
//             mat_A[454] * mat_B[205] +
//             mat_A[455] * mat_B[237] +
//             mat_A[456] * mat_B[269] +
//             mat_A[457] * mat_B[301] +
//             mat_A[458] * mat_B[333] +
//             mat_A[459] * mat_B[365] +
//             mat_A[460] * mat_B[397] +
//             mat_A[461] * mat_B[429] +
//             mat_A[462] * mat_B[461] +
//             mat_A[463] * mat_B[493] +
//             mat_A[464] * mat_B[525] +
//             mat_A[465] * mat_B[557] +
//             mat_A[466] * mat_B[589] +
//             mat_A[467] * mat_B[621] +
//             mat_A[468] * mat_B[653] +
//             mat_A[469] * mat_B[685] +
//             mat_A[470] * mat_B[717] +
//             mat_A[471] * mat_B[749] +
//             mat_A[472] * mat_B[781] +
//             mat_A[473] * mat_B[813] +
//             mat_A[474] * mat_B[845] +
//             mat_A[475] * mat_B[877] +
//             mat_A[476] * mat_B[909] +
//             mat_A[477] * mat_B[941] +
//             mat_A[478] * mat_B[973] +
//             mat_A[479] * mat_B[1005];
//  mat_C[462] <= 
//             mat_A[448] * mat_B[14] +
//             mat_A[449] * mat_B[46] +
//             mat_A[450] * mat_B[78] +
//             mat_A[451] * mat_B[110] +
//             mat_A[452] * mat_B[142] +
//             mat_A[453] * mat_B[174] +
//             mat_A[454] * mat_B[206] +
//             mat_A[455] * mat_B[238] +
//             mat_A[456] * mat_B[270] +
//             mat_A[457] * mat_B[302] +
//             mat_A[458] * mat_B[334] +
//             mat_A[459] * mat_B[366] +
//             mat_A[460] * mat_B[398] +
//             mat_A[461] * mat_B[430] +
//             mat_A[462] * mat_B[462] +
//             mat_A[463] * mat_B[494] +
//             mat_A[464] * mat_B[526] +
//             mat_A[465] * mat_B[558] +
//             mat_A[466] * mat_B[590] +
//             mat_A[467] * mat_B[622] +
//             mat_A[468] * mat_B[654] +
//             mat_A[469] * mat_B[686] +
//             mat_A[470] * mat_B[718] +
//             mat_A[471] * mat_B[750] +
//             mat_A[472] * mat_B[782] +
//             mat_A[473] * mat_B[814] +
//             mat_A[474] * mat_B[846] +
//             mat_A[475] * mat_B[878] +
//             mat_A[476] * mat_B[910] +
//             mat_A[477] * mat_B[942] +
//             mat_A[478] * mat_B[974] +
//             mat_A[479] * mat_B[1006];
//  mat_C[463] <= 
//             mat_A[448] * mat_B[15] +
//             mat_A[449] * mat_B[47] +
//             mat_A[450] * mat_B[79] +
//             mat_A[451] * mat_B[111] +
//             mat_A[452] * mat_B[143] +
//             mat_A[453] * mat_B[175] +
//             mat_A[454] * mat_B[207] +
//             mat_A[455] * mat_B[239] +
//             mat_A[456] * mat_B[271] +
//             mat_A[457] * mat_B[303] +
//             mat_A[458] * mat_B[335] +
//             mat_A[459] * mat_B[367] +
//             mat_A[460] * mat_B[399] +
//             mat_A[461] * mat_B[431] +
//             mat_A[462] * mat_B[463] +
//             mat_A[463] * mat_B[495] +
//             mat_A[464] * mat_B[527] +
//             mat_A[465] * mat_B[559] +
//             mat_A[466] * mat_B[591] +
//             mat_A[467] * mat_B[623] +
//             mat_A[468] * mat_B[655] +
//             mat_A[469] * mat_B[687] +
//             mat_A[470] * mat_B[719] +
//             mat_A[471] * mat_B[751] +
//             mat_A[472] * mat_B[783] +
//             mat_A[473] * mat_B[815] +
//             mat_A[474] * mat_B[847] +
//             mat_A[475] * mat_B[879] +
//             mat_A[476] * mat_B[911] +
//             mat_A[477] * mat_B[943] +
//             mat_A[478] * mat_B[975] +
//             mat_A[479] * mat_B[1007];
//  mat_C[464] <= 
//             mat_A[448] * mat_B[16] +
//             mat_A[449] * mat_B[48] +
//             mat_A[450] * mat_B[80] +
//             mat_A[451] * mat_B[112] +
//             mat_A[452] * mat_B[144] +
//             mat_A[453] * mat_B[176] +
//             mat_A[454] * mat_B[208] +
//             mat_A[455] * mat_B[240] +
//             mat_A[456] * mat_B[272] +
//             mat_A[457] * mat_B[304] +
//             mat_A[458] * mat_B[336] +
//             mat_A[459] * mat_B[368] +
//             mat_A[460] * mat_B[400] +
//             mat_A[461] * mat_B[432] +
//             mat_A[462] * mat_B[464] +
//             mat_A[463] * mat_B[496] +
//             mat_A[464] * mat_B[528] +
//             mat_A[465] * mat_B[560] +
//             mat_A[466] * mat_B[592] +
//             mat_A[467] * mat_B[624] +
//             mat_A[468] * mat_B[656] +
//             mat_A[469] * mat_B[688] +
//             mat_A[470] * mat_B[720] +
//             mat_A[471] * mat_B[752] +
//             mat_A[472] * mat_B[784] +
//             mat_A[473] * mat_B[816] +
//             mat_A[474] * mat_B[848] +
//             mat_A[475] * mat_B[880] +
//             mat_A[476] * mat_B[912] +
//             mat_A[477] * mat_B[944] +
//             mat_A[478] * mat_B[976] +
//             mat_A[479] * mat_B[1008];
//  mat_C[465] <= 
//             mat_A[448] * mat_B[17] +
//             mat_A[449] * mat_B[49] +
//             mat_A[450] * mat_B[81] +
//             mat_A[451] * mat_B[113] +
//             mat_A[452] * mat_B[145] +
//             mat_A[453] * mat_B[177] +
//             mat_A[454] * mat_B[209] +
//             mat_A[455] * mat_B[241] +
//             mat_A[456] * mat_B[273] +
//             mat_A[457] * mat_B[305] +
//             mat_A[458] * mat_B[337] +
//             mat_A[459] * mat_B[369] +
//             mat_A[460] * mat_B[401] +
//             mat_A[461] * mat_B[433] +
//             mat_A[462] * mat_B[465] +
//             mat_A[463] * mat_B[497] +
//             mat_A[464] * mat_B[529] +
//             mat_A[465] * mat_B[561] +
//             mat_A[466] * mat_B[593] +
//             mat_A[467] * mat_B[625] +
//             mat_A[468] * mat_B[657] +
//             mat_A[469] * mat_B[689] +
//             mat_A[470] * mat_B[721] +
//             mat_A[471] * mat_B[753] +
//             mat_A[472] * mat_B[785] +
//             mat_A[473] * mat_B[817] +
//             mat_A[474] * mat_B[849] +
//             mat_A[475] * mat_B[881] +
//             mat_A[476] * mat_B[913] +
//             mat_A[477] * mat_B[945] +
//             mat_A[478] * mat_B[977] +
//             mat_A[479] * mat_B[1009];
//  mat_C[466] <= 
//             mat_A[448] * mat_B[18] +
//             mat_A[449] * mat_B[50] +
//             mat_A[450] * mat_B[82] +
//             mat_A[451] * mat_B[114] +
//             mat_A[452] * mat_B[146] +
//             mat_A[453] * mat_B[178] +
//             mat_A[454] * mat_B[210] +
//             mat_A[455] * mat_B[242] +
//             mat_A[456] * mat_B[274] +
//             mat_A[457] * mat_B[306] +
//             mat_A[458] * mat_B[338] +
//             mat_A[459] * mat_B[370] +
//             mat_A[460] * mat_B[402] +
//             mat_A[461] * mat_B[434] +
//             mat_A[462] * mat_B[466] +
//             mat_A[463] * mat_B[498] +
//             mat_A[464] * mat_B[530] +
//             mat_A[465] * mat_B[562] +
//             mat_A[466] * mat_B[594] +
//             mat_A[467] * mat_B[626] +
//             mat_A[468] * mat_B[658] +
//             mat_A[469] * mat_B[690] +
//             mat_A[470] * mat_B[722] +
//             mat_A[471] * mat_B[754] +
//             mat_A[472] * mat_B[786] +
//             mat_A[473] * mat_B[818] +
//             mat_A[474] * mat_B[850] +
//             mat_A[475] * mat_B[882] +
//             mat_A[476] * mat_B[914] +
//             mat_A[477] * mat_B[946] +
//             mat_A[478] * mat_B[978] +
//             mat_A[479] * mat_B[1010];
//  mat_C[467] <= 
//             mat_A[448] * mat_B[19] +
//             mat_A[449] * mat_B[51] +
//             mat_A[450] * mat_B[83] +
//             mat_A[451] * mat_B[115] +
//             mat_A[452] * mat_B[147] +
//             mat_A[453] * mat_B[179] +
//             mat_A[454] * mat_B[211] +
//             mat_A[455] * mat_B[243] +
//             mat_A[456] * mat_B[275] +
//             mat_A[457] * mat_B[307] +
//             mat_A[458] * mat_B[339] +
//             mat_A[459] * mat_B[371] +
//             mat_A[460] * mat_B[403] +
//             mat_A[461] * mat_B[435] +
//             mat_A[462] * mat_B[467] +
//             mat_A[463] * mat_B[499] +
//             mat_A[464] * mat_B[531] +
//             mat_A[465] * mat_B[563] +
//             mat_A[466] * mat_B[595] +
//             mat_A[467] * mat_B[627] +
//             mat_A[468] * mat_B[659] +
//             mat_A[469] * mat_B[691] +
//             mat_A[470] * mat_B[723] +
//             mat_A[471] * mat_B[755] +
//             mat_A[472] * mat_B[787] +
//             mat_A[473] * mat_B[819] +
//             mat_A[474] * mat_B[851] +
//             mat_A[475] * mat_B[883] +
//             mat_A[476] * mat_B[915] +
//             mat_A[477] * mat_B[947] +
//             mat_A[478] * mat_B[979] +
//             mat_A[479] * mat_B[1011];
//  mat_C[468] <= 
//             mat_A[448] * mat_B[20] +
//             mat_A[449] * mat_B[52] +
//             mat_A[450] * mat_B[84] +
//             mat_A[451] * mat_B[116] +
//             mat_A[452] * mat_B[148] +
//             mat_A[453] * mat_B[180] +
//             mat_A[454] * mat_B[212] +
//             mat_A[455] * mat_B[244] +
//             mat_A[456] * mat_B[276] +
//             mat_A[457] * mat_B[308] +
//             mat_A[458] * mat_B[340] +
//             mat_A[459] * mat_B[372] +
//             mat_A[460] * mat_B[404] +
//             mat_A[461] * mat_B[436] +
//             mat_A[462] * mat_B[468] +
//             mat_A[463] * mat_B[500] +
//             mat_A[464] * mat_B[532] +
//             mat_A[465] * mat_B[564] +
//             mat_A[466] * mat_B[596] +
//             mat_A[467] * mat_B[628] +
//             mat_A[468] * mat_B[660] +
//             mat_A[469] * mat_B[692] +
//             mat_A[470] * mat_B[724] +
//             mat_A[471] * mat_B[756] +
//             mat_A[472] * mat_B[788] +
//             mat_A[473] * mat_B[820] +
//             mat_A[474] * mat_B[852] +
//             mat_A[475] * mat_B[884] +
//             mat_A[476] * mat_B[916] +
//             mat_A[477] * mat_B[948] +
//             mat_A[478] * mat_B[980] +
//             mat_A[479] * mat_B[1012];
//  mat_C[469] <= 
//             mat_A[448] * mat_B[21] +
//             mat_A[449] * mat_B[53] +
//             mat_A[450] * mat_B[85] +
//             mat_A[451] * mat_B[117] +
//             mat_A[452] * mat_B[149] +
//             mat_A[453] * mat_B[181] +
//             mat_A[454] * mat_B[213] +
//             mat_A[455] * mat_B[245] +
//             mat_A[456] * mat_B[277] +
//             mat_A[457] * mat_B[309] +
//             mat_A[458] * mat_B[341] +
//             mat_A[459] * mat_B[373] +
//             mat_A[460] * mat_B[405] +
//             mat_A[461] * mat_B[437] +
//             mat_A[462] * mat_B[469] +
//             mat_A[463] * mat_B[501] +
//             mat_A[464] * mat_B[533] +
//             mat_A[465] * mat_B[565] +
//             mat_A[466] * mat_B[597] +
//             mat_A[467] * mat_B[629] +
//             mat_A[468] * mat_B[661] +
//             mat_A[469] * mat_B[693] +
//             mat_A[470] * mat_B[725] +
//             mat_A[471] * mat_B[757] +
//             mat_A[472] * mat_B[789] +
//             mat_A[473] * mat_B[821] +
//             mat_A[474] * mat_B[853] +
//             mat_A[475] * mat_B[885] +
//             mat_A[476] * mat_B[917] +
//             mat_A[477] * mat_B[949] +
//             mat_A[478] * mat_B[981] +
//             mat_A[479] * mat_B[1013];
//  mat_C[470] <= 
//             mat_A[448] * mat_B[22] +
//             mat_A[449] * mat_B[54] +
//             mat_A[450] * mat_B[86] +
//             mat_A[451] * mat_B[118] +
//             mat_A[452] * mat_B[150] +
//             mat_A[453] * mat_B[182] +
//             mat_A[454] * mat_B[214] +
//             mat_A[455] * mat_B[246] +
//             mat_A[456] * mat_B[278] +
//             mat_A[457] * mat_B[310] +
//             mat_A[458] * mat_B[342] +
//             mat_A[459] * mat_B[374] +
//             mat_A[460] * mat_B[406] +
//             mat_A[461] * mat_B[438] +
//             mat_A[462] * mat_B[470] +
//             mat_A[463] * mat_B[502] +
//             mat_A[464] * mat_B[534] +
//             mat_A[465] * mat_B[566] +
//             mat_A[466] * mat_B[598] +
//             mat_A[467] * mat_B[630] +
//             mat_A[468] * mat_B[662] +
//             mat_A[469] * mat_B[694] +
//             mat_A[470] * mat_B[726] +
//             mat_A[471] * mat_B[758] +
//             mat_A[472] * mat_B[790] +
//             mat_A[473] * mat_B[822] +
//             mat_A[474] * mat_B[854] +
//             mat_A[475] * mat_B[886] +
//             mat_A[476] * mat_B[918] +
//             mat_A[477] * mat_B[950] +
//             mat_A[478] * mat_B[982] +
//             mat_A[479] * mat_B[1014];
//  mat_C[471] <= 
//             mat_A[448] * mat_B[23] +
//             mat_A[449] * mat_B[55] +
//             mat_A[450] * mat_B[87] +
//             mat_A[451] * mat_B[119] +
//             mat_A[452] * mat_B[151] +
//             mat_A[453] * mat_B[183] +
//             mat_A[454] * mat_B[215] +
//             mat_A[455] * mat_B[247] +
//             mat_A[456] * mat_B[279] +
//             mat_A[457] * mat_B[311] +
//             mat_A[458] * mat_B[343] +
//             mat_A[459] * mat_B[375] +
//             mat_A[460] * mat_B[407] +
//             mat_A[461] * mat_B[439] +
//             mat_A[462] * mat_B[471] +
//             mat_A[463] * mat_B[503] +
//             mat_A[464] * mat_B[535] +
//             mat_A[465] * mat_B[567] +
//             mat_A[466] * mat_B[599] +
//             mat_A[467] * mat_B[631] +
//             mat_A[468] * mat_B[663] +
//             mat_A[469] * mat_B[695] +
//             mat_A[470] * mat_B[727] +
//             mat_A[471] * mat_B[759] +
//             mat_A[472] * mat_B[791] +
//             mat_A[473] * mat_B[823] +
//             mat_A[474] * mat_B[855] +
//             mat_A[475] * mat_B[887] +
//             mat_A[476] * mat_B[919] +
//             mat_A[477] * mat_B[951] +
//             mat_A[478] * mat_B[983] +
//             mat_A[479] * mat_B[1015];
//  mat_C[472] <= 
//             mat_A[448] * mat_B[24] +
//             mat_A[449] * mat_B[56] +
//             mat_A[450] * mat_B[88] +
//             mat_A[451] * mat_B[120] +
//             mat_A[452] * mat_B[152] +
//             mat_A[453] * mat_B[184] +
//             mat_A[454] * mat_B[216] +
//             mat_A[455] * mat_B[248] +
//             mat_A[456] * mat_B[280] +
//             mat_A[457] * mat_B[312] +
//             mat_A[458] * mat_B[344] +
//             mat_A[459] * mat_B[376] +
//             mat_A[460] * mat_B[408] +
//             mat_A[461] * mat_B[440] +
//             mat_A[462] * mat_B[472] +
//             mat_A[463] * mat_B[504] +
//             mat_A[464] * mat_B[536] +
//             mat_A[465] * mat_B[568] +
//             mat_A[466] * mat_B[600] +
//             mat_A[467] * mat_B[632] +
//             mat_A[468] * mat_B[664] +
//             mat_A[469] * mat_B[696] +
//             mat_A[470] * mat_B[728] +
//             mat_A[471] * mat_B[760] +
//             mat_A[472] * mat_B[792] +
//             mat_A[473] * mat_B[824] +
//             mat_A[474] * mat_B[856] +
//             mat_A[475] * mat_B[888] +
//             mat_A[476] * mat_B[920] +
//             mat_A[477] * mat_B[952] +
//             mat_A[478] * mat_B[984] +
//             mat_A[479] * mat_B[1016];
//  mat_C[473] <= 
//             mat_A[448] * mat_B[25] +
//             mat_A[449] * mat_B[57] +
//             mat_A[450] * mat_B[89] +
//             mat_A[451] * mat_B[121] +
//             mat_A[452] * mat_B[153] +
//             mat_A[453] * mat_B[185] +
//             mat_A[454] * mat_B[217] +
//             mat_A[455] * mat_B[249] +
//             mat_A[456] * mat_B[281] +
//             mat_A[457] * mat_B[313] +
//             mat_A[458] * mat_B[345] +
//             mat_A[459] * mat_B[377] +
//             mat_A[460] * mat_B[409] +
//             mat_A[461] * mat_B[441] +
//             mat_A[462] * mat_B[473] +
//             mat_A[463] * mat_B[505] +
//             mat_A[464] * mat_B[537] +
//             mat_A[465] * mat_B[569] +
//             mat_A[466] * mat_B[601] +
//             mat_A[467] * mat_B[633] +
//             mat_A[468] * mat_B[665] +
//             mat_A[469] * mat_B[697] +
//             mat_A[470] * mat_B[729] +
//             mat_A[471] * mat_B[761] +
//             mat_A[472] * mat_B[793] +
//             mat_A[473] * mat_B[825] +
//             mat_A[474] * mat_B[857] +
//             mat_A[475] * mat_B[889] +
//             mat_A[476] * mat_B[921] +
//             mat_A[477] * mat_B[953] +
//             mat_A[478] * mat_B[985] +
//             mat_A[479] * mat_B[1017];
//  mat_C[474] <= 
//             mat_A[448] * mat_B[26] +
//             mat_A[449] * mat_B[58] +
//             mat_A[450] * mat_B[90] +
//             mat_A[451] * mat_B[122] +
//             mat_A[452] * mat_B[154] +
//             mat_A[453] * mat_B[186] +
//             mat_A[454] * mat_B[218] +
//             mat_A[455] * mat_B[250] +
//             mat_A[456] * mat_B[282] +
//             mat_A[457] * mat_B[314] +
//             mat_A[458] * mat_B[346] +
//             mat_A[459] * mat_B[378] +
//             mat_A[460] * mat_B[410] +
//             mat_A[461] * mat_B[442] +
//             mat_A[462] * mat_B[474] +
//             mat_A[463] * mat_B[506] +
//             mat_A[464] * mat_B[538] +
//             mat_A[465] * mat_B[570] +
//             mat_A[466] * mat_B[602] +
//             mat_A[467] * mat_B[634] +
//             mat_A[468] * mat_B[666] +
//             mat_A[469] * mat_B[698] +
//             mat_A[470] * mat_B[730] +
//             mat_A[471] * mat_B[762] +
//             mat_A[472] * mat_B[794] +
//             mat_A[473] * mat_B[826] +
//             mat_A[474] * mat_B[858] +
//             mat_A[475] * mat_B[890] +
//             mat_A[476] * mat_B[922] +
//             mat_A[477] * mat_B[954] +
//             mat_A[478] * mat_B[986] +
//             mat_A[479] * mat_B[1018];
//  mat_C[475] <= 
//             mat_A[448] * mat_B[27] +
//             mat_A[449] * mat_B[59] +
//             mat_A[450] * mat_B[91] +
//             mat_A[451] * mat_B[123] +
//             mat_A[452] * mat_B[155] +
//             mat_A[453] * mat_B[187] +
//             mat_A[454] * mat_B[219] +
//             mat_A[455] * mat_B[251] +
//             mat_A[456] * mat_B[283] +
//             mat_A[457] * mat_B[315] +
//             mat_A[458] * mat_B[347] +
//             mat_A[459] * mat_B[379] +
//             mat_A[460] * mat_B[411] +
//             mat_A[461] * mat_B[443] +
//             mat_A[462] * mat_B[475] +
//             mat_A[463] * mat_B[507] +
//             mat_A[464] * mat_B[539] +
//             mat_A[465] * mat_B[571] +
//             mat_A[466] * mat_B[603] +
//             mat_A[467] * mat_B[635] +
//             mat_A[468] * mat_B[667] +
//             mat_A[469] * mat_B[699] +
//             mat_A[470] * mat_B[731] +
//             mat_A[471] * mat_B[763] +
//             mat_A[472] * mat_B[795] +
//             mat_A[473] * mat_B[827] +
//             mat_A[474] * mat_B[859] +
//             mat_A[475] * mat_B[891] +
//             mat_A[476] * mat_B[923] +
//             mat_A[477] * mat_B[955] +
//             mat_A[478] * mat_B[987] +
//             mat_A[479] * mat_B[1019];
//  mat_C[476] <= 
//             mat_A[448] * mat_B[28] +
//             mat_A[449] * mat_B[60] +
//             mat_A[450] * mat_B[92] +
//             mat_A[451] * mat_B[124] +
//             mat_A[452] * mat_B[156] +
//             mat_A[453] * mat_B[188] +
//             mat_A[454] * mat_B[220] +
//             mat_A[455] * mat_B[252] +
//             mat_A[456] * mat_B[284] +
//             mat_A[457] * mat_B[316] +
//             mat_A[458] * mat_B[348] +
//             mat_A[459] * mat_B[380] +
//             mat_A[460] * mat_B[412] +
//             mat_A[461] * mat_B[444] +
//             mat_A[462] * mat_B[476] +
//             mat_A[463] * mat_B[508] +
//             mat_A[464] * mat_B[540] +
//             mat_A[465] * mat_B[572] +
//             mat_A[466] * mat_B[604] +
//             mat_A[467] * mat_B[636] +
//             mat_A[468] * mat_B[668] +
//             mat_A[469] * mat_B[700] +
//             mat_A[470] * mat_B[732] +
//             mat_A[471] * mat_B[764] +
//             mat_A[472] * mat_B[796] +
//             mat_A[473] * mat_B[828] +
//             mat_A[474] * mat_B[860] +
//             mat_A[475] * mat_B[892] +
//             mat_A[476] * mat_B[924] +
//             mat_A[477] * mat_B[956] +
//             mat_A[478] * mat_B[988] +
//             mat_A[479] * mat_B[1020];
//  mat_C[477] <= 
//             mat_A[448] * mat_B[29] +
//             mat_A[449] * mat_B[61] +
//             mat_A[450] * mat_B[93] +
//             mat_A[451] * mat_B[125] +
//             mat_A[452] * mat_B[157] +
//             mat_A[453] * mat_B[189] +
//             mat_A[454] * mat_B[221] +
//             mat_A[455] * mat_B[253] +
//             mat_A[456] * mat_B[285] +
//             mat_A[457] * mat_B[317] +
//             mat_A[458] * mat_B[349] +
//             mat_A[459] * mat_B[381] +
//             mat_A[460] * mat_B[413] +
//             mat_A[461] * mat_B[445] +
//             mat_A[462] * mat_B[477] +
//             mat_A[463] * mat_B[509] +
//             mat_A[464] * mat_B[541] +
//             mat_A[465] * mat_B[573] +
//             mat_A[466] * mat_B[605] +
//             mat_A[467] * mat_B[637] +
//             mat_A[468] * mat_B[669] +
//             mat_A[469] * mat_B[701] +
//             mat_A[470] * mat_B[733] +
//             mat_A[471] * mat_B[765] +
//             mat_A[472] * mat_B[797] +
//             mat_A[473] * mat_B[829] +
//             mat_A[474] * mat_B[861] +
//             mat_A[475] * mat_B[893] +
//             mat_A[476] * mat_B[925] +
//             mat_A[477] * mat_B[957] +
//             mat_A[478] * mat_B[989] +
//             mat_A[479] * mat_B[1021];
//  mat_C[478] <= 
//             mat_A[448] * mat_B[30] +
//             mat_A[449] * mat_B[62] +
//             mat_A[450] * mat_B[94] +
//             mat_A[451] * mat_B[126] +
//             mat_A[452] * mat_B[158] +
//             mat_A[453] * mat_B[190] +
//             mat_A[454] * mat_B[222] +
//             mat_A[455] * mat_B[254] +
//             mat_A[456] * mat_B[286] +
//             mat_A[457] * mat_B[318] +
//             mat_A[458] * mat_B[350] +
//             mat_A[459] * mat_B[382] +
//             mat_A[460] * mat_B[414] +
//             mat_A[461] * mat_B[446] +
//             mat_A[462] * mat_B[478] +
//             mat_A[463] * mat_B[510] +
//             mat_A[464] * mat_B[542] +
//             mat_A[465] * mat_B[574] +
//             mat_A[466] * mat_B[606] +
//             mat_A[467] * mat_B[638] +
//             mat_A[468] * mat_B[670] +
//             mat_A[469] * mat_B[702] +
//             mat_A[470] * mat_B[734] +
//             mat_A[471] * mat_B[766] +
//             mat_A[472] * mat_B[798] +
//             mat_A[473] * mat_B[830] +
//             mat_A[474] * mat_B[862] +
//             mat_A[475] * mat_B[894] +
//             mat_A[476] * mat_B[926] +
//             mat_A[477] * mat_B[958] +
//             mat_A[478] * mat_B[990] +
//             mat_A[479] * mat_B[1022];
//  mat_C[479] <= 
//             mat_A[448] * mat_B[31] +
//             mat_A[449] * mat_B[63] +
//             mat_A[450] * mat_B[95] +
//             mat_A[451] * mat_B[127] +
//             mat_A[452] * mat_B[159] +
//             mat_A[453] * mat_B[191] +
//             mat_A[454] * mat_B[223] +
//             mat_A[455] * mat_B[255] +
//             mat_A[456] * mat_B[287] +
//             mat_A[457] * mat_B[319] +
//             mat_A[458] * mat_B[351] +
//             mat_A[459] * mat_B[383] +
//             mat_A[460] * mat_B[415] +
//             mat_A[461] * mat_B[447] +
//             mat_A[462] * mat_B[479] +
//             mat_A[463] * mat_B[511] +
//             mat_A[464] * mat_B[543] +
//             mat_A[465] * mat_B[575] +
//             mat_A[466] * mat_B[607] +
//             mat_A[467] * mat_B[639] +
//             mat_A[468] * mat_B[671] +
//             mat_A[469] * mat_B[703] +
//             mat_A[470] * mat_B[735] +
//             mat_A[471] * mat_B[767] +
//             mat_A[472] * mat_B[799] +
//             mat_A[473] * mat_B[831] +
//             mat_A[474] * mat_B[863] +
//             mat_A[475] * mat_B[895] +
//             mat_A[476] * mat_B[927] +
//             mat_A[477] * mat_B[959] +
//             mat_A[478] * mat_B[991] +
//             mat_A[479] * mat_B[1023];
//  mat_C[480] <= 
//             mat_A[480] * mat_B[0] +
//             mat_A[481] * mat_B[32] +
//             mat_A[482] * mat_B[64] +
//             mat_A[483] * mat_B[96] +
//             mat_A[484] * mat_B[128] +
//             mat_A[485] * mat_B[160] +
//             mat_A[486] * mat_B[192] +
//             mat_A[487] * mat_B[224] +
//             mat_A[488] * mat_B[256] +
//             mat_A[489] * mat_B[288] +
//             mat_A[490] * mat_B[320] +
//             mat_A[491] * mat_B[352] +
//             mat_A[492] * mat_B[384] +
//             mat_A[493] * mat_B[416] +
//             mat_A[494] * mat_B[448] +
//             mat_A[495] * mat_B[480] +
//             mat_A[496] * mat_B[512] +
//             mat_A[497] * mat_B[544] +
//             mat_A[498] * mat_B[576] +
//             mat_A[499] * mat_B[608] +
//             mat_A[500] * mat_B[640] +
//             mat_A[501] * mat_B[672] +
//             mat_A[502] * mat_B[704] +
//             mat_A[503] * mat_B[736] +
//             mat_A[504] * mat_B[768] +
//             mat_A[505] * mat_B[800] +
//             mat_A[506] * mat_B[832] +
//             mat_A[507] * mat_B[864] +
//             mat_A[508] * mat_B[896] +
//             mat_A[509] * mat_B[928] +
//             mat_A[510] * mat_B[960] +
//             mat_A[511] * mat_B[992];
//  mat_C[481] <= 
//             mat_A[480] * mat_B[1] +
//             mat_A[481] * mat_B[33] +
//             mat_A[482] * mat_B[65] +
//             mat_A[483] * mat_B[97] +
//             mat_A[484] * mat_B[129] +
//             mat_A[485] * mat_B[161] +
//             mat_A[486] * mat_B[193] +
//             mat_A[487] * mat_B[225] +
//             mat_A[488] * mat_B[257] +
//             mat_A[489] * mat_B[289] +
//             mat_A[490] * mat_B[321] +
//             mat_A[491] * mat_B[353] +
//             mat_A[492] * mat_B[385] +
//             mat_A[493] * mat_B[417] +
//             mat_A[494] * mat_B[449] +
//             mat_A[495] * mat_B[481] +
//             mat_A[496] * mat_B[513] +
//             mat_A[497] * mat_B[545] +
//             mat_A[498] * mat_B[577] +
//             mat_A[499] * mat_B[609] +
//             mat_A[500] * mat_B[641] +
//             mat_A[501] * mat_B[673] +
//             mat_A[502] * mat_B[705] +
//             mat_A[503] * mat_B[737] +
//             mat_A[504] * mat_B[769] +
//             mat_A[505] * mat_B[801] +
//             mat_A[506] * mat_B[833] +
//             mat_A[507] * mat_B[865] +
//             mat_A[508] * mat_B[897] +
//             mat_A[509] * mat_B[929] +
//             mat_A[510] * mat_B[961] +
//             mat_A[511] * mat_B[993];
//  mat_C[482] <= 
//             mat_A[480] * mat_B[2] +
//             mat_A[481] * mat_B[34] +
//             mat_A[482] * mat_B[66] +
//             mat_A[483] * mat_B[98] +
//             mat_A[484] * mat_B[130] +
//             mat_A[485] * mat_B[162] +
//             mat_A[486] * mat_B[194] +
//             mat_A[487] * mat_B[226] +
//             mat_A[488] * mat_B[258] +
//             mat_A[489] * mat_B[290] +
//             mat_A[490] * mat_B[322] +
//             mat_A[491] * mat_B[354] +
//             mat_A[492] * mat_B[386] +
//             mat_A[493] * mat_B[418] +
//             mat_A[494] * mat_B[450] +
//             mat_A[495] * mat_B[482] +
//             mat_A[496] * mat_B[514] +
//             mat_A[497] * mat_B[546] +
//             mat_A[498] * mat_B[578] +
//             mat_A[499] * mat_B[610] +
//             mat_A[500] * mat_B[642] +
//             mat_A[501] * mat_B[674] +
//             mat_A[502] * mat_B[706] +
//             mat_A[503] * mat_B[738] +
//             mat_A[504] * mat_B[770] +
//             mat_A[505] * mat_B[802] +
//             mat_A[506] * mat_B[834] +
//             mat_A[507] * mat_B[866] +
//             mat_A[508] * mat_B[898] +
//             mat_A[509] * mat_B[930] +
//             mat_A[510] * mat_B[962] +
//             mat_A[511] * mat_B[994];
//  mat_C[483] <= 
//             mat_A[480] * mat_B[3] +
//             mat_A[481] * mat_B[35] +
//             mat_A[482] * mat_B[67] +
//             mat_A[483] * mat_B[99] +
//             mat_A[484] * mat_B[131] +
//             mat_A[485] * mat_B[163] +
//             mat_A[486] * mat_B[195] +
//             mat_A[487] * mat_B[227] +
//             mat_A[488] * mat_B[259] +
//             mat_A[489] * mat_B[291] +
//             mat_A[490] * mat_B[323] +
//             mat_A[491] * mat_B[355] +
//             mat_A[492] * mat_B[387] +
//             mat_A[493] * mat_B[419] +
//             mat_A[494] * mat_B[451] +
//             mat_A[495] * mat_B[483] +
//             mat_A[496] * mat_B[515] +
//             mat_A[497] * mat_B[547] +
//             mat_A[498] * mat_B[579] +
//             mat_A[499] * mat_B[611] +
//             mat_A[500] * mat_B[643] +
//             mat_A[501] * mat_B[675] +
//             mat_A[502] * mat_B[707] +
//             mat_A[503] * mat_B[739] +
//             mat_A[504] * mat_B[771] +
//             mat_A[505] * mat_B[803] +
//             mat_A[506] * mat_B[835] +
//             mat_A[507] * mat_B[867] +
//             mat_A[508] * mat_B[899] +
//             mat_A[509] * mat_B[931] +
//             mat_A[510] * mat_B[963] +
//             mat_A[511] * mat_B[995];
//  mat_C[484] <= 
//             mat_A[480] * mat_B[4] +
//             mat_A[481] * mat_B[36] +
//             mat_A[482] * mat_B[68] +
//             mat_A[483] * mat_B[100] +
//             mat_A[484] * mat_B[132] +
//             mat_A[485] * mat_B[164] +
//             mat_A[486] * mat_B[196] +
//             mat_A[487] * mat_B[228] +
//             mat_A[488] * mat_B[260] +
//             mat_A[489] * mat_B[292] +
//             mat_A[490] * mat_B[324] +
//             mat_A[491] * mat_B[356] +
//             mat_A[492] * mat_B[388] +
//             mat_A[493] * mat_B[420] +
//             mat_A[494] * mat_B[452] +
//             mat_A[495] * mat_B[484] +
//             mat_A[496] * mat_B[516] +
//             mat_A[497] * mat_B[548] +
//             mat_A[498] * mat_B[580] +
//             mat_A[499] * mat_B[612] +
//             mat_A[500] * mat_B[644] +
//             mat_A[501] * mat_B[676] +
//             mat_A[502] * mat_B[708] +
//             mat_A[503] * mat_B[740] +
//             mat_A[504] * mat_B[772] +
//             mat_A[505] * mat_B[804] +
//             mat_A[506] * mat_B[836] +
//             mat_A[507] * mat_B[868] +
//             mat_A[508] * mat_B[900] +
//             mat_A[509] * mat_B[932] +
//             mat_A[510] * mat_B[964] +
//             mat_A[511] * mat_B[996];
//  mat_C[485] <= 
//             mat_A[480] * mat_B[5] +
//             mat_A[481] * mat_B[37] +
//             mat_A[482] * mat_B[69] +
//             mat_A[483] * mat_B[101] +
//             mat_A[484] * mat_B[133] +
//             mat_A[485] * mat_B[165] +
//             mat_A[486] * mat_B[197] +
//             mat_A[487] * mat_B[229] +
//             mat_A[488] * mat_B[261] +
//             mat_A[489] * mat_B[293] +
//             mat_A[490] * mat_B[325] +
//             mat_A[491] * mat_B[357] +
//             mat_A[492] * mat_B[389] +
//             mat_A[493] * mat_B[421] +
//             mat_A[494] * mat_B[453] +
//             mat_A[495] * mat_B[485] +
//             mat_A[496] * mat_B[517] +
//             mat_A[497] * mat_B[549] +
//             mat_A[498] * mat_B[581] +
//             mat_A[499] * mat_B[613] +
//             mat_A[500] * mat_B[645] +
//             mat_A[501] * mat_B[677] +
//             mat_A[502] * mat_B[709] +
//             mat_A[503] * mat_B[741] +
//             mat_A[504] * mat_B[773] +
//             mat_A[505] * mat_B[805] +
//             mat_A[506] * mat_B[837] +
//             mat_A[507] * mat_B[869] +
//             mat_A[508] * mat_B[901] +
//             mat_A[509] * mat_B[933] +
//             mat_A[510] * mat_B[965] +
//             mat_A[511] * mat_B[997];
//  mat_C[486] <= 
//             mat_A[480] * mat_B[6] +
//             mat_A[481] * mat_B[38] +
//             mat_A[482] * mat_B[70] +
//             mat_A[483] * mat_B[102] +
//             mat_A[484] * mat_B[134] +
//             mat_A[485] * mat_B[166] +
//             mat_A[486] * mat_B[198] +
//             mat_A[487] * mat_B[230] +
//             mat_A[488] * mat_B[262] +
//             mat_A[489] * mat_B[294] +
//             mat_A[490] * mat_B[326] +
//             mat_A[491] * mat_B[358] +
//             mat_A[492] * mat_B[390] +
//             mat_A[493] * mat_B[422] +
//             mat_A[494] * mat_B[454] +
//             mat_A[495] * mat_B[486] +
//             mat_A[496] * mat_B[518] +
//             mat_A[497] * mat_B[550] +
//             mat_A[498] * mat_B[582] +
//             mat_A[499] * mat_B[614] +
//             mat_A[500] * mat_B[646] +
//             mat_A[501] * mat_B[678] +
//             mat_A[502] * mat_B[710] +
//             mat_A[503] * mat_B[742] +
//             mat_A[504] * mat_B[774] +
//             mat_A[505] * mat_B[806] +
//             mat_A[506] * mat_B[838] +
//             mat_A[507] * mat_B[870] +
//             mat_A[508] * mat_B[902] +
//             mat_A[509] * mat_B[934] +
//             mat_A[510] * mat_B[966] +
//             mat_A[511] * mat_B[998];
//  mat_C[487] <= 
//             mat_A[480] * mat_B[7] +
//             mat_A[481] * mat_B[39] +
//             mat_A[482] * mat_B[71] +
//             mat_A[483] * mat_B[103] +
//             mat_A[484] * mat_B[135] +
//             mat_A[485] * mat_B[167] +
//             mat_A[486] * mat_B[199] +
//             mat_A[487] * mat_B[231] +
//             mat_A[488] * mat_B[263] +
//             mat_A[489] * mat_B[295] +
//             mat_A[490] * mat_B[327] +
//             mat_A[491] * mat_B[359] +
//             mat_A[492] * mat_B[391] +
//             mat_A[493] * mat_B[423] +
//             mat_A[494] * mat_B[455] +
//             mat_A[495] * mat_B[487] +
//             mat_A[496] * mat_B[519] +
//             mat_A[497] * mat_B[551] +
//             mat_A[498] * mat_B[583] +
//             mat_A[499] * mat_B[615] +
//             mat_A[500] * mat_B[647] +
//             mat_A[501] * mat_B[679] +
//             mat_A[502] * mat_B[711] +
//             mat_A[503] * mat_B[743] +
//             mat_A[504] * mat_B[775] +
//             mat_A[505] * mat_B[807] +
//             mat_A[506] * mat_B[839] +
//             mat_A[507] * mat_B[871] +
//             mat_A[508] * mat_B[903] +
//             mat_A[509] * mat_B[935] +
//             mat_A[510] * mat_B[967] +
//             mat_A[511] * mat_B[999];
//  mat_C[488] <= 
//             mat_A[480] * mat_B[8] +
//             mat_A[481] * mat_B[40] +
//             mat_A[482] * mat_B[72] +
//             mat_A[483] * mat_B[104] +
//             mat_A[484] * mat_B[136] +
//             mat_A[485] * mat_B[168] +
//             mat_A[486] * mat_B[200] +
//             mat_A[487] * mat_B[232] +
//             mat_A[488] * mat_B[264] +
//             mat_A[489] * mat_B[296] +
//             mat_A[490] * mat_B[328] +
//             mat_A[491] * mat_B[360] +
//             mat_A[492] * mat_B[392] +
//             mat_A[493] * mat_B[424] +
//             mat_A[494] * mat_B[456] +
//             mat_A[495] * mat_B[488] +
//             mat_A[496] * mat_B[520] +
//             mat_A[497] * mat_B[552] +
//             mat_A[498] * mat_B[584] +
//             mat_A[499] * mat_B[616] +
//             mat_A[500] * mat_B[648] +
//             mat_A[501] * mat_B[680] +
//             mat_A[502] * mat_B[712] +
//             mat_A[503] * mat_B[744] +
//             mat_A[504] * mat_B[776] +
//             mat_A[505] * mat_B[808] +
//             mat_A[506] * mat_B[840] +
//             mat_A[507] * mat_B[872] +
//             mat_A[508] * mat_B[904] +
//             mat_A[509] * mat_B[936] +
//             mat_A[510] * mat_B[968] +
//             mat_A[511] * mat_B[1000];
//  mat_C[489] <= 
//             mat_A[480] * mat_B[9] +
//             mat_A[481] * mat_B[41] +
//             mat_A[482] * mat_B[73] +
//             mat_A[483] * mat_B[105] +
//             mat_A[484] * mat_B[137] +
//             mat_A[485] * mat_B[169] +
//             mat_A[486] * mat_B[201] +
//             mat_A[487] * mat_B[233] +
//             mat_A[488] * mat_B[265] +
//             mat_A[489] * mat_B[297] +
//             mat_A[490] * mat_B[329] +
//             mat_A[491] * mat_B[361] +
//             mat_A[492] * mat_B[393] +
//             mat_A[493] * mat_B[425] +
//             mat_A[494] * mat_B[457] +
//             mat_A[495] * mat_B[489] +
//             mat_A[496] * mat_B[521] +
//             mat_A[497] * mat_B[553] +
//             mat_A[498] * mat_B[585] +
//             mat_A[499] * mat_B[617] +
//             mat_A[500] * mat_B[649] +
//             mat_A[501] * mat_B[681] +
//             mat_A[502] * mat_B[713] +
//             mat_A[503] * mat_B[745] +
//             mat_A[504] * mat_B[777] +
//             mat_A[505] * mat_B[809] +
//             mat_A[506] * mat_B[841] +
//             mat_A[507] * mat_B[873] +
//             mat_A[508] * mat_B[905] +
//             mat_A[509] * mat_B[937] +
//             mat_A[510] * mat_B[969] +
//             mat_A[511] * mat_B[1001];
//  mat_C[490] <= 
//             mat_A[480] * mat_B[10] +
//             mat_A[481] * mat_B[42] +
//             mat_A[482] * mat_B[74] +
//             mat_A[483] * mat_B[106] +
//             mat_A[484] * mat_B[138] +
//             mat_A[485] * mat_B[170] +
//             mat_A[486] * mat_B[202] +
//             mat_A[487] * mat_B[234] +
//             mat_A[488] * mat_B[266] +
//             mat_A[489] * mat_B[298] +
//             mat_A[490] * mat_B[330] +
//             mat_A[491] * mat_B[362] +
//             mat_A[492] * mat_B[394] +
//             mat_A[493] * mat_B[426] +
//             mat_A[494] * mat_B[458] +
//             mat_A[495] * mat_B[490] +
//             mat_A[496] * mat_B[522] +
//             mat_A[497] * mat_B[554] +
//             mat_A[498] * mat_B[586] +
//             mat_A[499] * mat_B[618] +
//             mat_A[500] * mat_B[650] +
//             mat_A[501] * mat_B[682] +
//             mat_A[502] * mat_B[714] +
//             mat_A[503] * mat_B[746] +
//             mat_A[504] * mat_B[778] +
//             mat_A[505] * mat_B[810] +
//             mat_A[506] * mat_B[842] +
//             mat_A[507] * mat_B[874] +
//             mat_A[508] * mat_B[906] +
//             mat_A[509] * mat_B[938] +
//             mat_A[510] * mat_B[970] +
//             mat_A[511] * mat_B[1002];
//  mat_C[491] <= 
//             mat_A[480] * mat_B[11] +
//             mat_A[481] * mat_B[43] +
//             mat_A[482] * mat_B[75] +
//             mat_A[483] * mat_B[107] +
//             mat_A[484] * mat_B[139] +
//             mat_A[485] * mat_B[171] +
//             mat_A[486] * mat_B[203] +
//             mat_A[487] * mat_B[235] +
//             mat_A[488] * mat_B[267] +
//             mat_A[489] * mat_B[299] +
//             mat_A[490] * mat_B[331] +
//             mat_A[491] * mat_B[363] +
//             mat_A[492] * mat_B[395] +
//             mat_A[493] * mat_B[427] +
//             mat_A[494] * mat_B[459] +
//             mat_A[495] * mat_B[491] +
//             mat_A[496] * mat_B[523] +
//             mat_A[497] * mat_B[555] +
//             mat_A[498] * mat_B[587] +
//             mat_A[499] * mat_B[619] +
//             mat_A[500] * mat_B[651] +
//             mat_A[501] * mat_B[683] +
//             mat_A[502] * mat_B[715] +
//             mat_A[503] * mat_B[747] +
//             mat_A[504] * mat_B[779] +
//             mat_A[505] * mat_B[811] +
//             mat_A[506] * mat_B[843] +
//             mat_A[507] * mat_B[875] +
//             mat_A[508] * mat_B[907] +
//             mat_A[509] * mat_B[939] +
//             mat_A[510] * mat_B[971] +
//             mat_A[511] * mat_B[1003];
//  mat_C[492] <= 
//             mat_A[480] * mat_B[12] +
//             mat_A[481] * mat_B[44] +
//             mat_A[482] * mat_B[76] +
//             mat_A[483] * mat_B[108] +
//             mat_A[484] * mat_B[140] +
//             mat_A[485] * mat_B[172] +
//             mat_A[486] * mat_B[204] +
//             mat_A[487] * mat_B[236] +
//             mat_A[488] * mat_B[268] +
//             mat_A[489] * mat_B[300] +
//             mat_A[490] * mat_B[332] +
//             mat_A[491] * mat_B[364] +
//             mat_A[492] * mat_B[396] +
//             mat_A[493] * mat_B[428] +
//             mat_A[494] * mat_B[460] +
//             mat_A[495] * mat_B[492] +
//             mat_A[496] * mat_B[524] +
//             mat_A[497] * mat_B[556] +
//             mat_A[498] * mat_B[588] +
//             mat_A[499] * mat_B[620] +
//             mat_A[500] * mat_B[652] +
//             mat_A[501] * mat_B[684] +
//             mat_A[502] * mat_B[716] +
//             mat_A[503] * mat_B[748] +
//             mat_A[504] * mat_B[780] +
//             mat_A[505] * mat_B[812] +
//             mat_A[506] * mat_B[844] +
//             mat_A[507] * mat_B[876] +
//             mat_A[508] * mat_B[908] +
//             mat_A[509] * mat_B[940] +
//             mat_A[510] * mat_B[972] +
//             mat_A[511] * mat_B[1004];
//  mat_C[493] <= 
//             mat_A[480] * mat_B[13] +
//             mat_A[481] * mat_B[45] +
//             mat_A[482] * mat_B[77] +
//             mat_A[483] * mat_B[109] +
//             mat_A[484] * mat_B[141] +
//             mat_A[485] * mat_B[173] +
//             mat_A[486] * mat_B[205] +
//             mat_A[487] * mat_B[237] +
//             mat_A[488] * mat_B[269] +
//             mat_A[489] * mat_B[301] +
//             mat_A[490] * mat_B[333] +
//             mat_A[491] * mat_B[365] +
//             mat_A[492] * mat_B[397] +
//             mat_A[493] * mat_B[429] +
//             mat_A[494] * mat_B[461] +
//             mat_A[495] * mat_B[493] +
//             mat_A[496] * mat_B[525] +
//             mat_A[497] * mat_B[557] +
//             mat_A[498] * mat_B[589] +
//             mat_A[499] * mat_B[621] +
//             mat_A[500] * mat_B[653] +
//             mat_A[501] * mat_B[685] +
//             mat_A[502] * mat_B[717] +
//             mat_A[503] * mat_B[749] +
//             mat_A[504] * mat_B[781] +
//             mat_A[505] * mat_B[813] +
//             mat_A[506] * mat_B[845] +
//             mat_A[507] * mat_B[877] +
//             mat_A[508] * mat_B[909] +
//             mat_A[509] * mat_B[941] +
//             mat_A[510] * mat_B[973] +
//             mat_A[511] * mat_B[1005];
//  mat_C[494] <= 
//             mat_A[480] * mat_B[14] +
//             mat_A[481] * mat_B[46] +
//             mat_A[482] * mat_B[78] +
//             mat_A[483] * mat_B[110] +
//             mat_A[484] * mat_B[142] +
//             mat_A[485] * mat_B[174] +
//             mat_A[486] * mat_B[206] +
//             mat_A[487] * mat_B[238] +
//             mat_A[488] * mat_B[270] +
//             mat_A[489] * mat_B[302] +
//             mat_A[490] * mat_B[334] +
//             mat_A[491] * mat_B[366] +
//             mat_A[492] * mat_B[398] +
//             mat_A[493] * mat_B[430] +
//             mat_A[494] * mat_B[462] +
//             mat_A[495] * mat_B[494] +
//             mat_A[496] * mat_B[526] +
//             mat_A[497] * mat_B[558] +
//             mat_A[498] * mat_B[590] +
//             mat_A[499] * mat_B[622] +
//             mat_A[500] * mat_B[654] +
//             mat_A[501] * mat_B[686] +
//             mat_A[502] * mat_B[718] +
//             mat_A[503] * mat_B[750] +
//             mat_A[504] * mat_B[782] +
//             mat_A[505] * mat_B[814] +
//             mat_A[506] * mat_B[846] +
//             mat_A[507] * mat_B[878] +
//             mat_A[508] * mat_B[910] +
//             mat_A[509] * mat_B[942] +
//             mat_A[510] * mat_B[974] +
//             mat_A[511] * mat_B[1006];
//  mat_C[495] <= 
//             mat_A[480] * mat_B[15] +
//             mat_A[481] * mat_B[47] +
//             mat_A[482] * mat_B[79] +
//             mat_A[483] * mat_B[111] +
//             mat_A[484] * mat_B[143] +
//             mat_A[485] * mat_B[175] +
//             mat_A[486] * mat_B[207] +
//             mat_A[487] * mat_B[239] +
//             mat_A[488] * mat_B[271] +
//             mat_A[489] * mat_B[303] +
//             mat_A[490] * mat_B[335] +
//             mat_A[491] * mat_B[367] +
//             mat_A[492] * mat_B[399] +
//             mat_A[493] * mat_B[431] +
//             mat_A[494] * mat_B[463] +
//             mat_A[495] * mat_B[495] +
//             mat_A[496] * mat_B[527] +
//             mat_A[497] * mat_B[559] +
//             mat_A[498] * mat_B[591] +
//             mat_A[499] * mat_B[623] +
//             mat_A[500] * mat_B[655] +
//             mat_A[501] * mat_B[687] +
//             mat_A[502] * mat_B[719] +
//             mat_A[503] * mat_B[751] +
//             mat_A[504] * mat_B[783] +
//             mat_A[505] * mat_B[815] +
//             mat_A[506] * mat_B[847] +
//             mat_A[507] * mat_B[879] +
//             mat_A[508] * mat_B[911] +
//             mat_A[509] * mat_B[943] +
//             mat_A[510] * mat_B[975] +
//             mat_A[511] * mat_B[1007];
//  mat_C[496] <= 
//             mat_A[480] * mat_B[16] +
//             mat_A[481] * mat_B[48] +
//             mat_A[482] * mat_B[80] +
//             mat_A[483] * mat_B[112] +
//             mat_A[484] * mat_B[144] +
//             mat_A[485] * mat_B[176] +
//             mat_A[486] * mat_B[208] +
//             mat_A[487] * mat_B[240] +
//             mat_A[488] * mat_B[272] +
//             mat_A[489] * mat_B[304] +
//             mat_A[490] * mat_B[336] +
//             mat_A[491] * mat_B[368] +
//             mat_A[492] * mat_B[400] +
//             mat_A[493] * mat_B[432] +
//             mat_A[494] * mat_B[464] +
//             mat_A[495] * mat_B[496] +
//             mat_A[496] * mat_B[528] +
//             mat_A[497] * mat_B[560] +
//             mat_A[498] * mat_B[592] +
//             mat_A[499] * mat_B[624] +
//             mat_A[500] * mat_B[656] +
//             mat_A[501] * mat_B[688] +
//             mat_A[502] * mat_B[720] +
//             mat_A[503] * mat_B[752] +
//             mat_A[504] * mat_B[784] +
//             mat_A[505] * mat_B[816] +
//             mat_A[506] * mat_B[848] +
//             mat_A[507] * mat_B[880] +
//             mat_A[508] * mat_B[912] +
//             mat_A[509] * mat_B[944] +
//             mat_A[510] * mat_B[976] +
//             mat_A[511] * mat_B[1008];
//  mat_C[497] <= 
//             mat_A[480] * mat_B[17] +
//             mat_A[481] * mat_B[49] +
//             mat_A[482] * mat_B[81] +
//             mat_A[483] * mat_B[113] +
//             mat_A[484] * mat_B[145] +
//             mat_A[485] * mat_B[177] +
//             mat_A[486] * mat_B[209] +
//             mat_A[487] * mat_B[241] +
//             mat_A[488] * mat_B[273] +
//             mat_A[489] * mat_B[305] +
//             mat_A[490] * mat_B[337] +
//             mat_A[491] * mat_B[369] +
//             mat_A[492] * mat_B[401] +
//             mat_A[493] * mat_B[433] +
//             mat_A[494] * mat_B[465] +
//             mat_A[495] * mat_B[497] +
//             mat_A[496] * mat_B[529] +
//             mat_A[497] * mat_B[561] +
//             mat_A[498] * mat_B[593] +
//             mat_A[499] * mat_B[625] +
//             mat_A[500] * mat_B[657] +
//             mat_A[501] * mat_B[689] +
//             mat_A[502] * mat_B[721] +
//             mat_A[503] * mat_B[753] +
//             mat_A[504] * mat_B[785] +
//             mat_A[505] * mat_B[817] +
//             mat_A[506] * mat_B[849] +
//             mat_A[507] * mat_B[881] +
//             mat_A[508] * mat_B[913] +
//             mat_A[509] * mat_B[945] +
//             mat_A[510] * mat_B[977] +
//             mat_A[511] * mat_B[1009];
//  mat_C[498] <= 
//             mat_A[480] * mat_B[18] +
//             mat_A[481] * mat_B[50] +
//             mat_A[482] * mat_B[82] +
//             mat_A[483] * mat_B[114] +
//             mat_A[484] * mat_B[146] +
//             mat_A[485] * mat_B[178] +
//             mat_A[486] * mat_B[210] +
//             mat_A[487] * mat_B[242] +
//             mat_A[488] * mat_B[274] +
//             mat_A[489] * mat_B[306] +
//             mat_A[490] * mat_B[338] +
//             mat_A[491] * mat_B[370] +
//             mat_A[492] * mat_B[402] +
//             mat_A[493] * mat_B[434] +
//             mat_A[494] * mat_B[466] +
//             mat_A[495] * mat_B[498] +
//             mat_A[496] * mat_B[530] +
//             mat_A[497] * mat_B[562] +
//             mat_A[498] * mat_B[594] +
//             mat_A[499] * mat_B[626] +
//             mat_A[500] * mat_B[658] +
//             mat_A[501] * mat_B[690] +
//             mat_A[502] * mat_B[722] +
//             mat_A[503] * mat_B[754] +
//             mat_A[504] * mat_B[786] +
//             mat_A[505] * mat_B[818] +
//             mat_A[506] * mat_B[850] +
//             mat_A[507] * mat_B[882] +
//             mat_A[508] * mat_B[914] +
//             mat_A[509] * mat_B[946] +
//             mat_A[510] * mat_B[978] +
//             mat_A[511] * mat_B[1010];
//  mat_C[499] <= 
//             mat_A[480] * mat_B[19] +
//             mat_A[481] * mat_B[51] +
//             mat_A[482] * mat_B[83] +
//             mat_A[483] * mat_B[115] +
//             mat_A[484] * mat_B[147] +
//             mat_A[485] * mat_B[179] +
//             mat_A[486] * mat_B[211] +
//             mat_A[487] * mat_B[243] +
//             mat_A[488] * mat_B[275] +
//             mat_A[489] * mat_B[307] +
//             mat_A[490] * mat_B[339] +
//             mat_A[491] * mat_B[371] +
//             mat_A[492] * mat_B[403] +
//             mat_A[493] * mat_B[435] +
//             mat_A[494] * mat_B[467] +
//             mat_A[495] * mat_B[499] +
//             mat_A[496] * mat_B[531] +
//             mat_A[497] * mat_B[563] +
//             mat_A[498] * mat_B[595] +
//             mat_A[499] * mat_B[627] +
//             mat_A[500] * mat_B[659] +
//             mat_A[501] * mat_B[691] +
//             mat_A[502] * mat_B[723] +
//             mat_A[503] * mat_B[755] +
//             mat_A[504] * mat_B[787] +
//             mat_A[505] * mat_B[819] +
//             mat_A[506] * mat_B[851] +
//             mat_A[507] * mat_B[883] +
//             mat_A[508] * mat_B[915] +
//             mat_A[509] * mat_B[947] +
//             mat_A[510] * mat_B[979] +
//             mat_A[511] * mat_B[1011];
//  mat_C[500] <= 
//             mat_A[480] * mat_B[20] +
//             mat_A[481] * mat_B[52] +
//             mat_A[482] * mat_B[84] +
//             mat_A[483] * mat_B[116] +
//             mat_A[484] * mat_B[148] +
//             mat_A[485] * mat_B[180] +
//             mat_A[486] * mat_B[212] +
//             mat_A[487] * mat_B[244] +
//             mat_A[488] * mat_B[276] +
//             mat_A[489] * mat_B[308] +
//             mat_A[490] * mat_B[340] +
//             mat_A[491] * mat_B[372] +
//             mat_A[492] * mat_B[404] +
//             mat_A[493] * mat_B[436] +
//             mat_A[494] * mat_B[468] +
//             mat_A[495] * mat_B[500] +
//             mat_A[496] * mat_B[532] +
//             mat_A[497] * mat_B[564] +
//             mat_A[498] * mat_B[596] +
//             mat_A[499] * mat_B[628] +
//             mat_A[500] * mat_B[660] +
//             mat_A[501] * mat_B[692] +
//             mat_A[502] * mat_B[724] +
//             mat_A[503] * mat_B[756] +
//             mat_A[504] * mat_B[788] +
//             mat_A[505] * mat_B[820] +
//             mat_A[506] * mat_B[852] +
//             mat_A[507] * mat_B[884] +
//             mat_A[508] * mat_B[916] +
//             mat_A[509] * mat_B[948] +
//             mat_A[510] * mat_B[980] +
//             mat_A[511] * mat_B[1012];
//  mat_C[501] <= 
//             mat_A[480] * mat_B[21] +
//             mat_A[481] * mat_B[53] +
//             mat_A[482] * mat_B[85] +
//             mat_A[483] * mat_B[117] +
//             mat_A[484] * mat_B[149] +
//             mat_A[485] * mat_B[181] +
//             mat_A[486] * mat_B[213] +
//             mat_A[487] * mat_B[245] +
//             mat_A[488] * mat_B[277] +
//             mat_A[489] * mat_B[309] +
//             mat_A[490] * mat_B[341] +
//             mat_A[491] * mat_B[373] +
//             mat_A[492] * mat_B[405] +
//             mat_A[493] * mat_B[437] +
//             mat_A[494] * mat_B[469] +
//             mat_A[495] * mat_B[501] +
//             mat_A[496] * mat_B[533] +
//             mat_A[497] * mat_B[565] +
//             mat_A[498] * mat_B[597] +
//             mat_A[499] * mat_B[629] +
//             mat_A[500] * mat_B[661] +
//             mat_A[501] * mat_B[693] +
//             mat_A[502] * mat_B[725] +
//             mat_A[503] * mat_B[757] +
//             mat_A[504] * mat_B[789] +
//             mat_A[505] * mat_B[821] +
//             mat_A[506] * mat_B[853] +
//             mat_A[507] * mat_B[885] +
//             mat_A[508] * mat_B[917] +
//             mat_A[509] * mat_B[949] +
//             mat_A[510] * mat_B[981] +
//             mat_A[511] * mat_B[1013];
//  mat_C[502] <= 
//             mat_A[480] * mat_B[22] +
//             mat_A[481] * mat_B[54] +
//             mat_A[482] * mat_B[86] +
//             mat_A[483] * mat_B[118] +
//             mat_A[484] * mat_B[150] +
//             mat_A[485] * mat_B[182] +
//             mat_A[486] * mat_B[214] +
//             mat_A[487] * mat_B[246] +
//             mat_A[488] * mat_B[278] +
//             mat_A[489] * mat_B[310] +
//             mat_A[490] * mat_B[342] +
//             mat_A[491] * mat_B[374] +
//             mat_A[492] * mat_B[406] +
//             mat_A[493] * mat_B[438] +
//             mat_A[494] * mat_B[470] +
//             mat_A[495] * mat_B[502] +
//             mat_A[496] * mat_B[534] +
//             mat_A[497] * mat_B[566] +
//             mat_A[498] * mat_B[598] +
//             mat_A[499] * mat_B[630] +
//             mat_A[500] * mat_B[662] +
//             mat_A[501] * mat_B[694] +
//             mat_A[502] * mat_B[726] +
//             mat_A[503] * mat_B[758] +
//             mat_A[504] * mat_B[790] +
//             mat_A[505] * mat_B[822] +
//             mat_A[506] * mat_B[854] +
//             mat_A[507] * mat_B[886] +
//             mat_A[508] * mat_B[918] +
//             mat_A[509] * mat_B[950] +
//             mat_A[510] * mat_B[982] +
//             mat_A[511] * mat_B[1014];
//  mat_C[503] <= 
//             mat_A[480] * mat_B[23] +
//             mat_A[481] * mat_B[55] +
//             mat_A[482] * mat_B[87] +
//             mat_A[483] * mat_B[119] +
//             mat_A[484] * mat_B[151] +
//             mat_A[485] * mat_B[183] +
//             mat_A[486] * mat_B[215] +
//             mat_A[487] * mat_B[247] +
//             mat_A[488] * mat_B[279] +
//             mat_A[489] * mat_B[311] +
//             mat_A[490] * mat_B[343] +
//             mat_A[491] * mat_B[375] +
//             mat_A[492] * mat_B[407] +
//             mat_A[493] * mat_B[439] +
//             mat_A[494] * mat_B[471] +
//             mat_A[495] * mat_B[503] +
//             mat_A[496] * mat_B[535] +
//             mat_A[497] * mat_B[567] +
//             mat_A[498] * mat_B[599] +
//             mat_A[499] * mat_B[631] +
//             mat_A[500] * mat_B[663] +
//             mat_A[501] * mat_B[695] +
//             mat_A[502] * mat_B[727] +
//             mat_A[503] * mat_B[759] +
//             mat_A[504] * mat_B[791] +
//             mat_A[505] * mat_B[823] +
//             mat_A[506] * mat_B[855] +
//             mat_A[507] * mat_B[887] +
//             mat_A[508] * mat_B[919] +
//             mat_A[509] * mat_B[951] +
//             mat_A[510] * mat_B[983] +
//             mat_A[511] * mat_B[1015];
//  mat_C[504] <= 
//             mat_A[480] * mat_B[24] +
//             mat_A[481] * mat_B[56] +
//             mat_A[482] * mat_B[88] +
//             mat_A[483] * mat_B[120] +
//             mat_A[484] * mat_B[152] +
//             mat_A[485] * mat_B[184] +
//             mat_A[486] * mat_B[216] +
//             mat_A[487] * mat_B[248] +
//             mat_A[488] * mat_B[280] +
//             mat_A[489] * mat_B[312] +
//             mat_A[490] * mat_B[344] +
//             mat_A[491] * mat_B[376] +
//             mat_A[492] * mat_B[408] +
//             mat_A[493] * mat_B[440] +
//             mat_A[494] * mat_B[472] +
//             mat_A[495] * mat_B[504] +
//             mat_A[496] * mat_B[536] +
//             mat_A[497] * mat_B[568] +
//             mat_A[498] * mat_B[600] +
//             mat_A[499] * mat_B[632] +
//             mat_A[500] * mat_B[664] +
//             mat_A[501] * mat_B[696] +
//             mat_A[502] * mat_B[728] +
//             mat_A[503] * mat_B[760] +
//             mat_A[504] * mat_B[792] +
//             mat_A[505] * mat_B[824] +
//             mat_A[506] * mat_B[856] +
//             mat_A[507] * mat_B[888] +
//             mat_A[508] * mat_B[920] +
//             mat_A[509] * mat_B[952] +
//             mat_A[510] * mat_B[984] +
//             mat_A[511] * mat_B[1016];
//  mat_C[505] <= 
//             mat_A[480] * mat_B[25] +
//             mat_A[481] * mat_B[57] +
//             mat_A[482] * mat_B[89] +
//             mat_A[483] * mat_B[121] +
//             mat_A[484] * mat_B[153] +
//             mat_A[485] * mat_B[185] +
//             mat_A[486] * mat_B[217] +
//             mat_A[487] * mat_B[249] +
//             mat_A[488] * mat_B[281] +
//             mat_A[489] * mat_B[313] +
//             mat_A[490] * mat_B[345] +
//             mat_A[491] * mat_B[377] +
//             mat_A[492] * mat_B[409] +
//             mat_A[493] * mat_B[441] +
//             mat_A[494] * mat_B[473] +
//             mat_A[495] * mat_B[505] +
//             mat_A[496] * mat_B[537] +
//             mat_A[497] * mat_B[569] +
//             mat_A[498] * mat_B[601] +
//             mat_A[499] * mat_B[633] +
//             mat_A[500] * mat_B[665] +
//             mat_A[501] * mat_B[697] +
//             mat_A[502] * mat_B[729] +
//             mat_A[503] * mat_B[761] +
//             mat_A[504] * mat_B[793] +
//             mat_A[505] * mat_B[825] +
//             mat_A[506] * mat_B[857] +
//             mat_A[507] * mat_B[889] +
//             mat_A[508] * mat_B[921] +
//             mat_A[509] * mat_B[953] +
//             mat_A[510] * mat_B[985] +
//             mat_A[511] * mat_B[1017];
//  mat_C[506] <= 
//             mat_A[480] * mat_B[26] +
//             mat_A[481] * mat_B[58] +
//             mat_A[482] * mat_B[90] +
//             mat_A[483] * mat_B[122] +
//             mat_A[484] * mat_B[154] +
//             mat_A[485] * mat_B[186] +
//             mat_A[486] * mat_B[218] +
//             mat_A[487] * mat_B[250] +
//             mat_A[488] * mat_B[282] +
//             mat_A[489] * mat_B[314] +
//             mat_A[490] * mat_B[346] +
//             mat_A[491] * mat_B[378] +
//             mat_A[492] * mat_B[410] +
//             mat_A[493] * mat_B[442] +
//             mat_A[494] * mat_B[474] +
//             mat_A[495] * mat_B[506] +
//             mat_A[496] * mat_B[538] +
//             mat_A[497] * mat_B[570] +
//             mat_A[498] * mat_B[602] +
//             mat_A[499] * mat_B[634] +
//             mat_A[500] * mat_B[666] +
//             mat_A[501] * mat_B[698] +
//             mat_A[502] * mat_B[730] +
//             mat_A[503] * mat_B[762] +
//             mat_A[504] * mat_B[794] +
//             mat_A[505] * mat_B[826] +
//             mat_A[506] * mat_B[858] +
//             mat_A[507] * mat_B[890] +
//             mat_A[508] * mat_B[922] +
//             mat_A[509] * mat_B[954] +
//             mat_A[510] * mat_B[986] +
//             mat_A[511] * mat_B[1018];
//  mat_C[507] <= 
//             mat_A[480] * mat_B[27] +
//             mat_A[481] * mat_B[59] +
//             mat_A[482] * mat_B[91] +
//             mat_A[483] * mat_B[123] +
//             mat_A[484] * mat_B[155] +
//             mat_A[485] * mat_B[187] +
//             mat_A[486] * mat_B[219] +
//             mat_A[487] * mat_B[251] +
//             mat_A[488] * mat_B[283] +
//             mat_A[489] * mat_B[315] +
//             mat_A[490] * mat_B[347] +
//             mat_A[491] * mat_B[379] +
//             mat_A[492] * mat_B[411] +
//             mat_A[493] * mat_B[443] +
//             mat_A[494] * mat_B[475] +
//             mat_A[495] * mat_B[507] +
//             mat_A[496] * mat_B[539] +
//             mat_A[497] * mat_B[571] +
//             mat_A[498] * mat_B[603] +
//             mat_A[499] * mat_B[635] +
//             mat_A[500] * mat_B[667] +
//             mat_A[501] * mat_B[699] +
//             mat_A[502] * mat_B[731] +
//             mat_A[503] * mat_B[763] +
//             mat_A[504] * mat_B[795] +
//             mat_A[505] * mat_B[827] +
//             mat_A[506] * mat_B[859] +
//             mat_A[507] * mat_B[891] +
//             mat_A[508] * mat_B[923] +
//             mat_A[509] * mat_B[955] +
//             mat_A[510] * mat_B[987] +
//             mat_A[511] * mat_B[1019];
//  mat_C[508] <= 
//             mat_A[480] * mat_B[28] +
//             mat_A[481] * mat_B[60] +
//             mat_A[482] * mat_B[92] +
//             mat_A[483] * mat_B[124] +
//             mat_A[484] * mat_B[156] +
//             mat_A[485] * mat_B[188] +
//             mat_A[486] * mat_B[220] +
//             mat_A[487] * mat_B[252] +
//             mat_A[488] * mat_B[284] +
//             mat_A[489] * mat_B[316] +
//             mat_A[490] * mat_B[348] +
//             mat_A[491] * mat_B[380] +
//             mat_A[492] * mat_B[412] +
//             mat_A[493] * mat_B[444] +
//             mat_A[494] * mat_B[476] +
//             mat_A[495] * mat_B[508] +
//             mat_A[496] * mat_B[540] +
//             mat_A[497] * mat_B[572] +
//             mat_A[498] * mat_B[604] +
//             mat_A[499] * mat_B[636] +
//             mat_A[500] * mat_B[668] +
//             mat_A[501] * mat_B[700] +
//             mat_A[502] * mat_B[732] +
//             mat_A[503] * mat_B[764] +
//             mat_A[504] * mat_B[796] +
//             mat_A[505] * mat_B[828] +
//             mat_A[506] * mat_B[860] +
//             mat_A[507] * mat_B[892] +
//             mat_A[508] * mat_B[924] +
//             mat_A[509] * mat_B[956] +
//             mat_A[510] * mat_B[988] +
//             mat_A[511] * mat_B[1020];
//  mat_C[509] <= 
//             mat_A[480] * mat_B[29] +
//             mat_A[481] * mat_B[61] +
//             mat_A[482] * mat_B[93] +
//             mat_A[483] * mat_B[125] +
//             mat_A[484] * mat_B[157] +
//             mat_A[485] * mat_B[189] +
//             mat_A[486] * mat_B[221] +
//             mat_A[487] * mat_B[253] +
//             mat_A[488] * mat_B[285] +
//             mat_A[489] * mat_B[317] +
//             mat_A[490] * mat_B[349] +
//             mat_A[491] * mat_B[381] +
//             mat_A[492] * mat_B[413] +
//             mat_A[493] * mat_B[445] +
//             mat_A[494] * mat_B[477] +
//             mat_A[495] * mat_B[509] +
//             mat_A[496] * mat_B[541] +
//             mat_A[497] * mat_B[573] +
//             mat_A[498] * mat_B[605] +
//             mat_A[499] * mat_B[637] +
//             mat_A[500] * mat_B[669] +
//             mat_A[501] * mat_B[701] +
//             mat_A[502] * mat_B[733] +
//             mat_A[503] * mat_B[765] +
//             mat_A[504] * mat_B[797] +
//             mat_A[505] * mat_B[829] +
//             mat_A[506] * mat_B[861] +
//             mat_A[507] * mat_B[893] +
//             mat_A[508] * mat_B[925] +
//             mat_A[509] * mat_B[957] +
//             mat_A[510] * mat_B[989] +
//             mat_A[511] * mat_B[1021];
//  mat_C[510] <= 
//             mat_A[480] * mat_B[30] +
//             mat_A[481] * mat_B[62] +
//             mat_A[482] * mat_B[94] +
//             mat_A[483] * mat_B[126] +
//             mat_A[484] * mat_B[158] +
//             mat_A[485] * mat_B[190] +
//             mat_A[486] * mat_B[222] +
//             mat_A[487] * mat_B[254] +
//             mat_A[488] * mat_B[286] +
//             mat_A[489] * mat_B[318] +
//             mat_A[490] * mat_B[350] +
//             mat_A[491] * mat_B[382] +
//             mat_A[492] * mat_B[414] +
//             mat_A[493] * mat_B[446] +
//             mat_A[494] * mat_B[478] +
//             mat_A[495] * mat_B[510] +
//             mat_A[496] * mat_B[542] +
//             mat_A[497] * mat_B[574] +
//             mat_A[498] * mat_B[606] +
//             mat_A[499] * mat_B[638] +
//             mat_A[500] * mat_B[670] +
//             mat_A[501] * mat_B[702] +
//             mat_A[502] * mat_B[734] +
//             mat_A[503] * mat_B[766] +
//             mat_A[504] * mat_B[798] +
//             mat_A[505] * mat_B[830] +
//             mat_A[506] * mat_B[862] +
//             mat_A[507] * mat_B[894] +
//             mat_A[508] * mat_B[926] +
//             mat_A[509] * mat_B[958] +
//             mat_A[510] * mat_B[990] +
//             mat_A[511] * mat_B[1022];
//  mat_C[511] <= 
//             mat_A[480] * mat_B[31] +
//             mat_A[481] * mat_B[63] +
//             mat_A[482] * mat_B[95] +
//             mat_A[483] * mat_B[127] +
//             mat_A[484] * mat_B[159] +
//             mat_A[485] * mat_B[191] +
//             mat_A[486] * mat_B[223] +
//             mat_A[487] * mat_B[255] +
//             mat_A[488] * mat_B[287] +
//             mat_A[489] * mat_B[319] +
//             mat_A[490] * mat_B[351] +
//             mat_A[491] * mat_B[383] +
//             mat_A[492] * mat_B[415] +
//             mat_A[493] * mat_B[447] +
//             mat_A[494] * mat_B[479] +
//             mat_A[495] * mat_B[511] +
//             mat_A[496] * mat_B[543] +
//             mat_A[497] * mat_B[575] +
//             mat_A[498] * mat_B[607] +
//             mat_A[499] * mat_B[639] +
//             mat_A[500] * mat_B[671] +
//             mat_A[501] * mat_B[703] +
//             mat_A[502] * mat_B[735] +
//             mat_A[503] * mat_B[767] +
//             mat_A[504] * mat_B[799] +
//             mat_A[505] * mat_B[831] +
//             mat_A[506] * mat_B[863] +
//             mat_A[507] * mat_B[895] +
//             mat_A[508] * mat_B[927] +
//             mat_A[509] * mat_B[959] +
//             mat_A[510] * mat_B[991] +
//             mat_A[511] * mat_B[1023];
//  mat_C[512] <= 
//             mat_A[512] * mat_B[0] +
//             mat_A[513] * mat_B[32] +
//             mat_A[514] * mat_B[64] +
//             mat_A[515] * mat_B[96] +
//             mat_A[516] * mat_B[128] +
//             mat_A[517] * mat_B[160] +
//             mat_A[518] * mat_B[192] +
//             mat_A[519] * mat_B[224] +
//             mat_A[520] * mat_B[256] +
//             mat_A[521] * mat_B[288] +
//             mat_A[522] * mat_B[320] +
//             mat_A[523] * mat_B[352] +
//             mat_A[524] * mat_B[384] +
//             mat_A[525] * mat_B[416] +
//             mat_A[526] * mat_B[448] +
//             mat_A[527] * mat_B[480] +
//             mat_A[528] * mat_B[512] +
//             mat_A[529] * mat_B[544] +
//             mat_A[530] * mat_B[576] +
//             mat_A[531] * mat_B[608] +
//             mat_A[532] * mat_B[640] +
//             mat_A[533] * mat_B[672] +
//             mat_A[534] * mat_B[704] +
//             mat_A[535] * mat_B[736] +
//             mat_A[536] * mat_B[768] +
//             mat_A[537] * mat_B[800] +
//             mat_A[538] * mat_B[832] +
//             mat_A[539] * mat_B[864] +
//             mat_A[540] * mat_B[896] +
//             mat_A[541] * mat_B[928] +
//             mat_A[542] * mat_B[960] +
//             mat_A[543] * mat_B[992];
//  mat_C[513] <= 
//             mat_A[512] * mat_B[1] +
//             mat_A[513] * mat_B[33] +
//             mat_A[514] * mat_B[65] +
//             mat_A[515] * mat_B[97] +
//             mat_A[516] * mat_B[129] +
//             mat_A[517] * mat_B[161] +
//             mat_A[518] * mat_B[193] +
//             mat_A[519] * mat_B[225] +
//             mat_A[520] * mat_B[257] +
//             mat_A[521] * mat_B[289] +
//             mat_A[522] * mat_B[321] +
//             mat_A[523] * mat_B[353] +
//             mat_A[524] * mat_B[385] +
//             mat_A[525] * mat_B[417] +
//             mat_A[526] * mat_B[449] +
//             mat_A[527] * mat_B[481] +
//             mat_A[528] * mat_B[513] +
//             mat_A[529] * mat_B[545] +
//             mat_A[530] * mat_B[577] +
//             mat_A[531] * mat_B[609] +
//             mat_A[532] * mat_B[641] +
//             mat_A[533] * mat_B[673] +
//             mat_A[534] * mat_B[705] +
//             mat_A[535] * mat_B[737] +
//             mat_A[536] * mat_B[769] +
//             mat_A[537] * mat_B[801] +
//             mat_A[538] * mat_B[833] +
//             mat_A[539] * mat_B[865] +
//             mat_A[540] * mat_B[897] +
//             mat_A[541] * mat_B[929] +
//             mat_A[542] * mat_B[961] +
//             mat_A[543] * mat_B[993];
//  mat_C[514] <= 
//             mat_A[512] * mat_B[2] +
//             mat_A[513] * mat_B[34] +
//             mat_A[514] * mat_B[66] +
//             mat_A[515] * mat_B[98] +
//             mat_A[516] * mat_B[130] +
//             mat_A[517] * mat_B[162] +
//             mat_A[518] * mat_B[194] +
//             mat_A[519] * mat_B[226] +
//             mat_A[520] * mat_B[258] +
//             mat_A[521] * mat_B[290] +
//             mat_A[522] * mat_B[322] +
//             mat_A[523] * mat_B[354] +
//             mat_A[524] * mat_B[386] +
//             mat_A[525] * mat_B[418] +
//             mat_A[526] * mat_B[450] +
//             mat_A[527] * mat_B[482] +
//             mat_A[528] * mat_B[514] +
//             mat_A[529] * mat_B[546] +
//             mat_A[530] * mat_B[578] +
//             mat_A[531] * mat_B[610] +
//             mat_A[532] * mat_B[642] +
//             mat_A[533] * mat_B[674] +
//             mat_A[534] * mat_B[706] +
//             mat_A[535] * mat_B[738] +
//             mat_A[536] * mat_B[770] +
//             mat_A[537] * mat_B[802] +
//             mat_A[538] * mat_B[834] +
//             mat_A[539] * mat_B[866] +
//             mat_A[540] * mat_B[898] +
//             mat_A[541] * mat_B[930] +
//             mat_A[542] * mat_B[962] +
//             mat_A[543] * mat_B[994];
//  mat_C[515] <= 
//             mat_A[512] * mat_B[3] +
//             mat_A[513] * mat_B[35] +
//             mat_A[514] * mat_B[67] +
//             mat_A[515] * mat_B[99] +
//             mat_A[516] * mat_B[131] +
//             mat_A[517] * mat_B[163] +
//             mat_A[518] * mat_B[195] +
//             mat_A[519] * mat_B[227] +
//             mat_A[520] * mat_B[259] +
//             mat_A[521] * mat_B[291] +
//             mat_A[522] * mat_B[323] +
//             mat_A[523] * mat_B[355] +
//             mat_A[524] * mat_B[387] +
//             mat_A[525] * mat_B[419] +
//             mat_A[526] * mat_B[451] +
//             mat_A[527] * mat_B[483] +
//             mat_A[528] * mat_B[515] +
//             mat_A[529] * mat_B[547] +
//             mat_A[530] * mat_B[579] +
//             mat_A[531] * mat_B[611] +
//             mat_A[532] * mat_B[643] +
//             mat_A[533] * mat_B[675] +
//             mat_A[534] * mat_B[707] +
//             mat_A[535] * mat_B[739] +
//             mat_A[536] * mat_B[771] +
//             mat_A[537] * mat_B[803] +
//             mat_A[538] * mat_B[835] +
//             mat_A[539] * mat_B[867] +
//             mat_A[540] * mat_B[899] +
//             mat_A[541] * mat_B[931] +
//             mat_A[542] * mat_B[963] +
//             mat_A[543] * mat_B[995];
//  mat_C[516] <= 
//             mat_A[512] * mat_B[4] +
//             mat_A[513] * mat_B[36] +
//             mat_A[514] * mat_B[68] +
//             mat_A[515] * mat_B[100] +
//             mat_A[516] * mat_B[132] +
//             mat_A[517] * mat_B[164] +
//             mat_A[518] * mat_B[196] +
//             mat_A[519] * mat_B[228] +
//             mat_A[520] * mat_B[260] +
//             mat_A[521] * mat_B[292] +
//             mat_A[522] * mat_B[324] +
//             mat_A[523] * mat_B[356] +
//             mat_A[524] * mat_B[388] +
//             mat_A[525] * mat_B[420] +
//             mat_A[526] * mat_B[452] +
//             mat_A[527] * mat_B[484] +
//             mat_A[528] * mat_B[516] +
//             mat_A[529] * mat_B[548] +
//             mat_A[530] * mat_B[580] +
//             mat_A[531] * mat_B[612] +
//             mat_A[532] * mat_B[644] +
//             mat_A[533] * mat_B[676] +
//             mat_A[534] * mat_B[708] +
//             mat_A[535] * mat_B[740] +
//             mat_A[536] * mat_B[772] +
//             mat_A[537] * mat_B[804] +
//             mat_A[538] * mat_B[836] +
//             mat_A[539] * mat_B[868] +
//             mat_A[540] * mat_B[900] +
//             mat_A[541] * mat_B[932] +
//             mat_A[542] * mat_B[964] +
//             mat_A[543] * mat_B[996];
//  mat_C[517] <= 
//             mat_A[512] * mat_B[5] +
//             mat_A[513] * mat_B[37] +
//             mat_A[514] * mat_B[69] +
//             mat_A[515] * mat_B[101] +
//             mat_A[516] * mat_B[133] +
//             mat_A[517] * mat_B[165] +
//             mat_A[518] * mat_B[197] +
//             mat_A[519] * mat_B[229] +
//             mat_A[520] * mat_B[261] +
//             mat_A[521] * mat_B[293] +
//             mat_A[522] * mat_B[325] +
//             mat_A[523] * mat_B[357] +
//             mat_A[524] * mat_B[389] +
//             mat_A[525] * mat_B[421] +
//             mat_A[526] * mat_B[453] +
//             mat_A[527] * mat_B[485] +
//             mat_A[528] * mat_B[517] +
//             mat_A[529] * mat_B[549] +
//             mat_A[530] * mat_B[581] +
//             mat_A[531] * mat_B[613] +
//             mat_A[532] * mat_B[645] +
//             mat_A[533] * mat_B[677] +
//             mat_A[534] * mat_B[709] +
//             mat_A[535] * mat_B[741] +
//             mat_A[536] * mat_B[773] +
//             mat_A[537] * mat_B[805] +
//             mat_A[538] * mat_B[837] +
//             mat_A[539] * mat_B[869] +
//             mat_A[540] * mat_B[901] +
//             mat_A[541] * mat_B[933] +
//             mat_A[542] * mat_B[965] +
//             mat_A[543] * mat_B[997];
//  mat_C[518] <= 
//             mat_A[512] * mat_B[6] +
//             mat_A[513] * mat_B[38] +
//             mat_A[514] * mat_B[70] +
//             mat_A[515] * mat_B[102] +
//             mat_A[516] * mat_B[134] +
//             mat_A[517] * mat_B[166] +
//             mat_A[518] * mat_B[198] +
//             mat_A[519] * mat_B[230] +
//             mat_A[520] * mat_B[262] +
//             mat_A[521] * mat_B[294] +
//             mat_A[522] * mat_B[326] +
//             mat_A[523] * mat_B[358] +
//             mat_A[524] * mat_B[390] +
//             mat_A[525] * mat_B[422] +
//             mat_A[526] * mat_B[454] +
//             mat_A[527] * mat_B[486] +
//             mat_A[528] * mat_B[518] +
//             mat_A[529] * mat_B[550] +
//             mat_A[530] * mat_B[582] +
//             mat_A[531] * mat_B[614] +
//             mat_A[532] * mat_B[646] +
//             mat_A[533] * mat_B[678] +
//             mat_A[534] * mat_B[710] +
//             mat_A[535] * mat_B[742] +
//             mat_A[536] * mat_B[774] +
//             mat_A[537] * mat_B[806] +
//             mat_A[538] * mat_B[838] +
//             mat_A[539] * mat_B[870] +
//             mat_A[540] * mat_B[902] +
//             mat_A[541] * mat_B[934] +
//             mat_A[542] * mat_B[966] +
//             mat_A[543] * mat_B[998];
//  mat_C[519] <= 
//             mat_A[512] * mat_B[7] +
//             mat_A[513] * mat_B[39] +
//             mat_A[514] * mat_B[71] +
//             mat_A[515] * mat_B[103] +
//             mat_A[516] * mat_B[135] +
//             mat_A[517] * mat_B[167] +
//             mat_A[518] * mat_B[199] +
//             mat_A[519] * mat_B[231] +
//             mat_A[520] * mat_B[263] +
//             mat_A[521] * mat_B[295] +
//             mat_A[522] * mat_B[327] +
//             mat_A[523] * mat_B[359] +
//             mat_A[524] * mat_B[391] +
//             mat_A[525] * mat_B[423] +
//             mat_A[526] * mat_B[455] +
//             mat_A[527] * mat_B[487] +
//             mat_A[528] * mat_B[519] +
//             mat_A[529] * mat_B[551] +
//             mat_A[530] * mat_B[583] +
//             mat_A[531] * mat_B[615] +
//             mat_A[532] * mat_B[647] +
//             mat_A[533] * mat_B[679] +
//             mat_A[534] * mat_B[711] +
//             mat_A[535] * mat_B[743] +
//             mat_A[536] * mat_B[775] +
//             mat_A[537] * mat_B[807] +
//             mat_A[538] * mat_B[839] +
//             mat_A[539] * mat_B[871] +
//             mat_A[540] * mat_B[903] +
//             mat_A[541] * mat_B[935] +
//             mat_A[542] * mat_B[967] +
//             mat_A[543] * mat_B[999];
//  mat_C[520] <= 
//             mat_A[512] * mat_B[8] +
//             mat_A[513] * mat_B[40] +
//             mat_A[514] * mat_B[72] +
//             mat_A[515] * mat_B[104] +
//             mat_A[516] * mat_B[136] +
//             mat_A[517] * mat_B[168] +
//             mat_A[518] * mat_B[200] +
//             mat_A[519] * mat_B[232] +
//             mat_A[520] * mat_B[264] +
//             mat_A[521] * mat_B[296] +
//             mat_A[522] * mat_B[328] +
//             mat_A[523] * mat_B[360] +
//             mat_A[524] * mat_B[392] +
//             mat_A[525] * mat_B[424] +
//             mat_A[526] * mat_B[456] +
//             mat_A[527] * mat_B[488] +
//             mat_A[528] * mat_B[520] +
//             mat_A[529] * mat_B[552] +
//             mat_A[530] * mat_B[584] +
//             mat_A[531] * mat_B[616] +
//             mat_A[532] * mat_B[648] +
//             mat_A[533] * mat_B[680] +
//             mat_A[534] * mat_B[712] +
//             mat_A[535] * mat_B[744] +
//             mat_A[536] * mat_B[776] +
//             mat_A[537] * mat_B[808] +
//             mat_A[538] * mat_B[840] +
//             mat_A[539] * mat_B[872] +
//             mat_A[540] * mat_B[904] +
//             mat_A[541] * mat_B[936] +
//             mat_A[542] * mat_B[968] +
//             mat_A[543] * mat_B[1000];
//  mat_C[521] <= 
//             mat_A[512] * mat_B[9] +
//             mat_A[513] * mat_B[41] +
//             mat_A[514] * mat_B[73] +
//             mat_A[515] * mat_B[105] +
//             mat_A[516] * mat_B[137] +
//             mat_A[517] * mat_B[169] +
//             mat_A[518] * mat_B[201] +
//             mat_A[519] * mat_B[233] +
//             mat_A[520] * mat_B[265] +
//             mat_A[521] * mat_B[297] +
//             mat_A[522] * mat_B[329] +
//             mat_A[523] * mat_B[361] +
//             mat_A[524] * mat_B[393] +
//             mat_A[525] * mat_B[425] +
//             mat_A[526] * mat_B[457] +
//             mat_A[527] * mat_B[489] +
//             mat_A[528] * mat_B[521] +
//             mat_A[529] * mat_B[553] +
//             mat_A[530] * mat_B[585] +
//             mat_A[531] * mat_B[617] +
//             mat_A[532] * mat_B[649] +
//             mat_A[533] * mat_B[681] +
//             mat_A[534] * mat_B[713] +
//             mat_A[535] * mat_B[745] +
//             mat_A[536] * mat_B[777] +
//             mat_A[537] * mat_B[809] +
//             mat_A[538] * mat_B[841] +
//             mat_A[539] * mat_B[873] +
//             mat_A[540] * mat_B[905] +
//             mat_A[541] * mat_B[937] +
//             mat_A[542] * mat_B[969] +
//             mat_A[543] * mat_B[1001];
//  mat_C[522] <= 
//             mat_A[512] * mat_B[10] +
//             mat_A[513] * mat_B[42] +
//             mat_A[514] * mat_B[74] +
//             mat_A[515] * mat_B[106] +
//             mat_A[516] * mat_B[138] +
//             mat_A[517] * mat_B[170] +
//             mat_A[518] * mat_B[202] +
//             mat_A[519] * mat_B[234] +
//             mat_A[520] * mat_B[266] +
//             mat_A[521] * mat_B[298] +
//             mat_A[522] * mat_B[330] +
//             mat_A[523] * mat_B[362] +
//             mat_A[524] * mat_B[394] +
//             mat_A[525] * mat_B[426] +
//             mat_A[526] * mat_B[458] +
//             mat_A[527] * mat_B[490] +
//             mat_A[528] * mat_B[522] +
//             mat_A[529] * mat_B[554] +
//             mat_A[530] * mat_B[586] +
//             mat_A[531] * mat_B[618] +
//             mat_A[532] * mat_B[650] +
//             mat_A[533] * mat_B[682] +
//             mat_A[534] * mat_B[714] +
//             mat_A[535] * mat_B[746] +
//             mat_A[536] * mat_B[778] +
//             mat_A[537] * mat_B[810] +
//             mat_A[538] * mat_B[842] +
//             mat_A[539] * mat_B[874] +
//             mat_A[540] * mat_B[906] +
//             mat_A[541] * mat_B[938] +
//             mat_A[542] * mat_B[970] +
//             mat_A[543] * mat_B[1002];
//  mat_C[523] <= 
//             mat_A[512] * mat_B[11] +
//             mat_A[513] * mat_B[43] +
//             mat_A[514] * mat_B[75] +
//             mat_A[515] * mat_B[107] +
//             mat_A[516] * mat_B[139] +
//             mat_A[517] * mat_B[171] +
//             mat_A[518] * mat_B[203] +
//             mat_A[519] * mat_B[235] +
//             mat_A[520] * mat_B[267] +
//             mat_A[521] * mat_B[299] +
//             mat_A[522] * mat_B[331] +
//             mat_A[523] * mat_B[363] +
//             mat_A[524] * mat_B[395] +
//             mat_A[525] * mat_B[427] +
//             mat_A[526] * mat_B[459] +
//             mat_A[527] * mat_B[491] +
//             mat_A[528] * mat_B[523] +
//             mat_A[529] * mat_B[555] +
//             mat_A[530] * mat_B[587] +
//             mat_A[531] * mat_B[619] +
//             mat_A[532] * mat_B[651] +
//             mat_A[533] * mat_B[683] +
//             mat_A[534] * mat_B[715] +
//             mat_A[535] * mat_B[747] +
//             mat_A[536] * mat_B[779] +
//             mat_A[537] * mat_B[811] +
//             mat_A[538] * mat_B[843] +
//             mat_A[539] * mat_B[875] +
//             mat_A[540] * mat_B[907] +
//             mat_A[541] * mat_B[939] +
//             mat_A[542] * mat_B[971] +
//             mat_A[543] * mat_B[1003];
//  mat_C[524] <= 
//             mat_A[512] * mat_B[12] +
//             mat_A[513] * mat_B[44] +
//             mat_A[514] * mat_B[76] +
//             mat_A[515] * mat_B[108] +
//             mat_A[516] * mat_B[140] +
//             mat_A[517] * mat_B[172] +
//             mat_A[518] * mat_B[204] +
//             mat_A[519] * mat_B[236] +
//             mat_A[520] * mat_B[268] +
//             mat_A[521] * mat_B[300] +
//             mat_A[522] * mat_B[332] +
//             mat_A[523] * mat_B[364] +
//             mat_A[524] * mat_B[396] +
//             mat_A[525] * mat_B[428] +
//             mat_A[526] * mat_B[460] +
//             mat_A[527] * mat_B[492] +
//             mat_A[528] * mat_B[524] +
//             mat_A[529] * mat_B[556] +
//             mat_A[530] * mat_B[588] +
//             mat_A[531] * mat_B[620] +
//             mat_A[532] * mat_B[652] +
//             mat_A[533] * mat_B[684] +
//             mat_A[534] * mat_B[716] +
//             mat_A[535] * mat_B[748] +
//             mat_A[536] * mat_B[780] +
//             mat_A[537] * mat_B[812] +
//             mat_A[538] * mat_B[844] +
//             mat_A[539] * mat_B[876] +
//             mat_A[540] * mat_B[908] +
//             mat_A[541] * mat_B[940] +
//             mat_A[542] * mat_B[972] +
//             mat_A[543] * mat_B[1004];
//  mat_C[525] <= 
//             mat_A[512] * mat_B[13] +
//             mat_A[513] * mat_B[45] +
//             mat_A[514] * mat_B[77] +
//             mat_A[515] * mat_B[109] +
//             mat_A[516] * mat_B[141] +
//             mat_A[517] * mat_B[173] +
//             mat_A[518] * mat_B[205] +
//             mat_A[519] * mat_B[237] +
//             mat_A[520] * mat_B[269] +
//             mat_A[521] * mat_B[301] +
//             mat_A[522] * mat_B[333] +
//             mat_A[523] * mat_B[365] +
//             mat_A[524] * mat_B[397] +
//             mat_A[525] * mat_B[429] +
//             mat_A[526] * mat_B[461] +
//             mat_A[527] * mat_B[493] +
//             mat_A[528] * mat_B[525] +
//             mat_A[529] * mat_B[557] +
//             mat_A[530] * mat_B[589] +
//             mat_A[531] * mat_B[621] +
//             mat_A[532] * mat_B[653] +
//             mat_A[533] * mat_B[685] +
//             mat_A[534] * mat_B[717] +
//             mat_A[535] * mat_B[749] +
//             mat_A[536] * mat_B[781] +
//             mat_A[537] * mat_B[813] +
//             mat_A[538] * mat_B[845] +
//             mat_A[539] * mat_B[877] +
//             mat_A[540] * mat_B[909] +
//             mat_A[541] * mat_B[941] +
//             mat_A[542] * mat_B[973] +
//             mat_A[543] * mat_B[1005];
//  mat_C[526] <= 
//             mat_A[512] * mat_B[14] +
//             mat_A[513] * mat_B[46] +
//             mat_A[514] * mat_B[78] +
//             mat_A[515] * mat_B[110] +
//             mat_A[516] * mat_B[142] +
//             mat_A[517] * mat_B[174] +
//             mat_A[518] * mat_B[206] +
//             mat_A[519] * mat_B[238] +
//             mat_A[520] * mat_B[270] +
//             mat_A[521] * mat_B[302] +
//             mat_A[522] * mat_B[334] +
//             mat_A[523] * mat_B[366] +
//             mat_A[524] * mat_B[398] +
//             mat_A[525] * mat_B[430] +
//             mat_A[526] * mat_B[462] +
//             mat_A[527] * mat_B[494] +
//             mat_A[528] * mat_B[526] +
//             mat_A[529] * mat_B[558] +
//             mat_A[530] * mat_B[590] +
//             mat_A[531] * mat_B[622] +
//             mat_A[532] * mat_B[654] +
//             mat_A[533] * mat_B[686] +
//             mat_A[534] * mat_B[718] +
//             mat_A[535] * mat_B[750] +
//             mat_A[536] * mat_B[782] +
//             mat_A[537] * mat_B[814] +
//             mat_A[538] * mat_B[846] +
//             mat_A[539] * mat_B[878] +
//             mat_A[540] * mat_B[910] +
//             mat_A[541] * mat_B[942] +
//             mat_A[542] * mat_B[974] +
//             mat_A[543] * mat_B[1006];
//  mat_C[527] <= 
//             mat_A[512] * mat_B[15] +
//             mat_A[513] * mat_B[47] +
//             mat_A[514] * mat_B[79] +
//             mat_A[515] * mat_B[111] +
//             mat_A[516] * mat_B[143] +
//             mat_A[517] * mat_B[175] +
//             mat_A[518] * mat_B[207] +
//             mat_A[519] * mat_B[239] +
//             mat_A[520] * mat_B[271] +
//             mat_A[521] * mat_B[303] +
//             mat_A[522] * mat_B[335] +
//             mat_A[523] * mat_B[367] +
//             mat_A[524] * mat_B[399] +
//             mat_A[525] * mat_B[431] +
//             mat_A[526] * mat_B[463] +
//             mat_A[527] * mat_B[495] +
//             mat_A[528] * mat_B[527] +
//             mat_A[529] * mat_B[559] +
//             mat_A[530] * mat_B[591] +
//             mat_A[531] * mat_B[623] +
//             mat_A[532] * mat_B[655] +
//             mat_A[533] * mat_B[687] +
//             mat_A[534] * mat_B[719] +
//             mat_A[535] * mat_B[751] +
//             mat_A[536] * mat_B[783] +
//             mat_A[537] * mat_B[815] +
//             mat_A[538] * mat_B[847] +
//             mat_A[539] * mat_B[879] +
//             mat_A[540] * mat_B[911] +
//             mat_A[541] * mat_B[943] +
//             mat_A[542] * mat_B[975] +
//             mat_A[543] * mat_B[1007];
//  mat_C[528] <= 
//             mat_A[512] * mat_B[16] +
//             mat_A[513] * mat_B[48] +
//             mat_A[514] * mat_B[80] +
//             mat_A[515] * mat_B[112] +
//             mat_A[516] * mat_B[144] +
//             mat_A[517] * mat_B[176] +
//             mat_A[518] * mat_B[208] +
//             mat_A[519] * mat_B[240] +
//             mat_A[520] * mat_B[272] +
//             mat_A[521] * mat_B[304] +
//             mat_A[522] * mat_B[336] +
//             mat_A[523] * mat_B[368] +
//             mat_A[524] * mat_B[400] +
//             mat_A[525] * mat_B[432] +
//             mat_A[526] * mat_B[464] +
//             mat_A[527] * mat_B[496] +
//             mat_A[528] * mat_B[528] +
//             mat_A[529] * mat_B[560] +
//             mat_A[530] * mat_B[592] +
//             mat_A[531] * mat_B[624] +
//             mat_A[532] * mat_B[656] +
//             mat_A[533] * mat_B[688] +
//             mat_A[534] * mat_B[720] +
//             mat_A[535] * mat_B[752] +
//             mat_A[536] * mat_B[784] +
//             mat_A[537] * mat_B[816] +
//             mat_A[538] * mat_B[848] +
//             mat_A[539] * mat_B[880] +
//             mat_A[540] * mat_B[912] +
//             mat_A[541] * mat_B[944] +
//             mat_A[542] * mat_B[976] +
//             mat_A[543] * mat_B[1008];
//  mat_C[529] <= 
//             mat_A[512] * mat_B[17] +
//             mat_A[513] * mat_B[49] +
//             mat_A[514] * mat_B[81] +
//             mat_A[515] * mat_B[113] +
//             mat_A[516] * mat_B[145] +
//             mat_A[517] * mat_B[177] +
//             mat_A[518] * mat_B[209] +
//             mat_A[519] * mat_B[241] +
//             mat_A[520] * mat_B[273] +
//             mat_A[521] * mat_B[305] +
//             mat_A[522] * mat_B[337] +
//             mat_A[523] * mat_B[369] +
//             mat_A[524] * mat_B[401] +
//             mat_A[525] * mat_B[433] +
//             mat_A[526] * mat_B[465] +
//             mat_A[527] * mat_B[497] +
//             mat_A[528] * mat_B[529] +
//             mat_A[529] * mat_B[561] +
//             mat_A[530] * mat_B[593] +
//             mat_A[531] * mat_B[625] +
//             mat_A[532] * mat_B[657] +
//             mat_A[533] * mat_B[689] +
//             mat_A[534] * mat_B[721] +
//             mat_A[535] * mat_B[753] +
//             mat_A[536] * mat_B[785] +
//             mat_A[537] * mat_B[817] +
//             mat_A[538] * mat_B[849] +
//             mat_A[539] * mat_B[881] +
//             mat_A[540] * mat_B[913] +
//             mat_A[541] * mat_B[945] +
//             mat_A[542] * mat_B[977] +
//             mat_A[543] * mat_B[1009];
//  mat_C[530] <= 
//             mat_A[512] * mat_B[18] +
//             mat_A[513] * mat_B[50] +
//             mat_A[514] * mat_B[82] +
//             mat_A[515] * mat_B[114] +
//             mat_A[516] * mat_B[146] +
//             mat_A[517] * mat_B[178] +
//             mat_A[518] * mat_B[210] +
//             mat_A[519] * mat_B[242] +
//             mat_A[520] * mat_B[274] +
//             mat_A[521] * mat_B[306] +
//             mat_A[522] * mat_B[338] +
//             mat_A[523] * mat_B[370] +
//             mat_A[524] * mat_B[402] +
//             mat_A[525] * mat_B[434] +
//             mat_A[526] * mat_B[466] +
//             mat_A[527] * mat_B[498] +
//             mat_A[528] * mat_B[530] +
//             mat_A[529] * mat_B[562] +
//             mat_A[530] * mat_B[594] +
//             mat_A[531] * mat_B[626] +
//             mat_A[532] * mat_B[658] +
//             mat_A[533] * mat_B[690] +
//             mat_A[534] * mat_B[722] +
//             mat_A[535] * mat_B[754] +
//             mat_A[536] * mat_B[786] +
//             mat_A[537] * mat_B[818] +
//             mat_A[538] * mat_B[850] +
//             mat_A[539] * mat_B[882] +
//             mat_A[540] * mat_B[914] +
//             mat_A[541] * mat_B[946] +
//             mat_A[542] * mat_B[978] +
//             mat_A[543] * mat_B[1010];
//  mat_C[531] <= 
//             mat_A[512] * mat_B[19] +
//             mat_A[513] * mat_B[51] +
//             mat_A[514] * mat_B[83] +
//             mat_A[515] * mat_B[115] +
//             mat_A[516] * mat_B[147] +
//             mat_A[517] * mat_B[179] +
//             mat_A[518] * mat_B[211] +
//             mat_A[519] * mat_B[243] +
//             mat_A[520] * mat_B[275] +
//             mat_A[521] * mat_B[307] +
//             mat_A[522] * mat_B[339] +
//             mat_A[523] * mat_B[371] +
//             mat_A[524] * mat_B[403] +
//             mat_A[525] * mat_B[435] +
//             mat_A[526] * mat_B[467] +
//             mat_A[527] * mat_B[499] +
//             mat_A[528] * mat_B[531] +
//             mat_A[529] * mat_B[563] +
//             mat_A[530] * mat_B[595] +
//             mat_A[531] * mat_B[627] +
//             mat_A[532] * mat_B[659] +
//             mat_A[533] * mat_B[691] +
//             mat_A[534] * mat_B[723] +
//             mat_A[535] * mat_B[755] +
//             mat_A[536] * mat_B[787] +
//             mat_A[537] * mat_B[819] +
//             mat_A[538] * mat_B[851] +
//             mat_A[539] * mat_B[883] +
//             mat_A[540] * mat_B[915] +
//             mat_A[541] * mat_B[947] +
//             mat_A[542] * mat_B[979] +
//             mat_A[543] * mat_B[1011];
//  mat_C[532] <= 
//             mat_A[512] * mat_B[20] +
//             mat_A[513] * mat_B[52] +
//             mat_A[514] * mat_B[84] +
//             mat_A[515] * mat_B[116] +
//             mat_A[516] * mat_B[148] +
//             mat_A[517] * mat_B[180] +
//             mat_A[518] * mat_B[212] +
//             mat_A[519] * mat_B[244] +
//             mat_A[520] * mat_B[276] +
//             mat_A[521] * mat_B[308] +
//             mat_A[522] * mat_B[340] +
//             mat_A[523] * mat_B[372] +
//             mat_A[524] * mat_B[404] +
//             mat_A[525] * mat_B[436] +
//             mat_A[526] * mat_B[468] +
//             mat_A[527] * mat_B[500] +
//             mat_A[528] * mat_B[532] +
//             mat_A[529] * mat_B[564] +
//             mat_A[530] * mat_B[596] +
//             mat_A[531] * mat_B[628] +
//             mat_A[532] * mat_B[660] +
//             mat_A[533] * mat_B[692] +
//             mat_A[534] * mat_B[724] +
//             mat_A[535] * mat_B[756] +
//             mat_A[536] * mat_B[788] +
//             mat_A[537] * mat_B[820] +
//             mat_A[538] * mat_B[852] +
//             mat_A[539] * mat_B[884] +
//             mat_A[540] * mat_B[916] +
//             mat_A[541] * mat_B[948] +
//             mat_A[542] * mat_B[980] +
//             mat_A[543] * mat_B[1012];
//  mat_C[533] <= 
//             mat_A[512] * mat_B[21] +
//             mat_A[513] * mat_B[53] +
//             mat_A[514] * mat_B[85] +
//             mat_A[515] * mat_B[117] +
//             mat_A[516] * mat_B[149] +
//             mat_A[517] * mat_B[181] +
//             mat_A[518] * mat_B[213] +
//             mat_A[519] * mat_B[245] +
//             mat_A[520] * mat_B[277] +
//             mat_A[521] * mat_B[309] +
//             mat_A[522] * mat_B[341] +
//             mat_A[523] * mat_B[373] +
//             mat_A[524] * mat_B[405] +
//             mat_A[525] * mat_B[437] +
//             mat_A[526] * mat_B[469] +
//             mat_A[527] * mat_B[501] +
//             mat_A[528] * mat_B[533] +
//             mat_A[529] * mat_B[565] +
//             mat_A[530] * mat_B[597] +
//             mat_A[531] * mat_B[629] +
//             mat_A[532] * mat_B[661] +
//             mat_A[533] * mat_B[693] +
//             mat_A[534] * mat_B[725] +
//             mat_A[535] * mat_B[757] +
//             mat_A[536] * mat_B[789] +
//             mat_A[537] * mat_B[821] +
//             mat_A[538] * mat_B[853] +
//             mat_A[539] * mat_B[885] +
//             mat_A[540] * mat_B[917] +
//             mat_A[541] * mat_B[949] +
//             mat_A[542] * mat_B[981] +
//             mat_A[543] * mat_B[1013];
//  mat_C[534] <= 
//             mat_A[512] * mat_B[22] +
//             mat_A[513] * mat_B[54] +
//             mat_A[514] * mat_B[86] +
//             mat_A[515] * mat_B[118] +
//             mat_A[516] * mat_B[150] +
//             mat_A[517] * mat_B[182] +
//             mat_A[518] * mat_B[214] +
//             mat_A[519] * mat_B[246] +
//             mat_A[520] * mat_B[278] +
//             mat_A[521] * mat_B[310] +
//             mat_A[522] * mat_B[342] +
//             mat_A[523] * mat_B[374] +
//             mat_A[524] * mat_B[406] +
//             mat_A[525] * mat_B[438] +
//             mat_A[526] * mat_B[470] +
//             mat_A[527] * mat_B[502] +
//             mat_A[528] * mat_B[534] +
//             mat_A[529] * mat_B[566] +
//             mat_A[530] * mat_B[598] +
//             mat_A[531] * mat_B[630] +
//             mat_A[532] * mat_B[662] +
//             mat_A[533] * mat_B[694] +
//             mat_A[534] * mat_B[726] +
//             mat_A[535] * mat_B[758] +
//             mat_A[536] * mat_B[790] +
//             mat_A[537] * mat_B[822] +
//             mat_A[538] * mat_B[854] +
//             mat_A[539] * mat_B[886] +
//             mat_A[540] * mat_B[918] +
//             mat_A[541] * mat_B[950] +
//             mat_A[542] * mat_B[982] +
//             mat_A[543] * mat_B[1014];
//  mat_C[535] <= 
//             mat_A[512] * mat_B[23] +
//             mat_A[513] * mat_B[55] +
//             mat_A[514] * mat_B[87] +
//             mat_A[515] * mat_B[119] +
//             mat_A[516] * mat_B[151] +
//             mat_A[517] * mat_B[183] +
//             mat_A[518] * mat_B[215] +
//             mat_A[519] * mat_B[247] +
//             mat_A[520] * mat_B[279] +
//             mat_A[521] * mat_B[311] +
//             mat_A[522] * mat_B[343] +
//             mat_A[523] * mat_B[375] +
//             mat_A[524] * mat_B[407] +
//             mat_A[525] * mat_B[439] +
//             mat_A[526] * mat_B[471] +
//             mat_A[527] * mat_B[503] +
//             mat_A[528] * mat_B[535] +
//             mat_A[529] * mat_B[567] +
//             mat_A[530] * mat_B[599] +
//             mat_A[531] * mat_B[631] +
//             mat_A[532] * mat_B[663] +
//             mat_A[533] * mat_B[695] +
//             mat_A[534] * mat_B[727] +
//             mat_A[535] * mat_B[759] +
//             mat_A[536] * mat_B[791] +
//             mat_A[537] * mat_B[823] +
//             mat_A[538] * mat_B[855] +
//             mat_A[539] * mat_B[887] +
//             mat_A[540] * mat_B[919] +
//             mat_A[541] * mat_B[951] +
//             mat_A[542] * mat_B[983] +
//             mat_A[543] * mat_B[1015];
//  mat_C[536] <= 
//             mat_A[512] * mat_B[24] +
//             mat_A[513] * mat_B[56] +
//             mat_A[514] * mat_B[88] +
//             mat_A[515] * mat_B[120] +
//             mat_A[516] * mat_B[152] +
//             mat_A[517] * mat_B[184] +
//             mat_A[518] * mat_B[216] +
//             mat_A[519] * mat_B[248] +
//             mat_A[520] * mat_B[280] +
//             mat_A[521] * mat_B[312] +
//             mat_A[522] * mat_B[344] +
//             mat_A[523] * mat_B[376] +
//             mat_A[524] * mat_B[408] +
//             mat_A[525] * mat_B[440] +
//             mat_A[526] * mat_B[472] +
//             mat_A[527] * mat_B[504] +
//             mat_A[528] * mat_B[536] +
//             mat_A[529] * mat_B[568] +
//             mat_A[530] * mat_B[600] +
//             mat_A[531] * mat_B[632] +
//             mat_A[532] * mat_B[664] +
//             mat_A[533] * mat_B[696] +
//             mat_A[534] * mat_B[728] +
//             mat_A[535] * mat_B[760] +
//             mat_A[536] * mat_B[792] +
//             mat_A[537] * mat_B[824] +
//             mat_A[538] * mat_B[856] +
//             mat_A[539] * mat_B[888] +
//             mat_A[540] * mat_B[920] +
//             mat_A[541] * mat_B[952] +
//             mat_A[542] * mat_B[984] +
//             mat_A[543] * mat_B[1016];
//  mat_C[537] <= 
//             mat_A[512] * mat_B[25] +
//             mat_A[513] * mat_B[57] +
//             mat_A[514] * mat_B[89] +
//             mat_A[515] * mat_B[121] +
//             mat_A[516] * mat_B[153] +
//             mat_A[517] * mat_B[185] +
//             mat_A[518] * mat_B[217] +
//             mat_A[519] * mat_B[249] +
//             mat_A[520] * mat_B[281] +
//             mat_A[521] * mat_B[313] +
//             mat_A[522] * mat_B[345] +
//             mat_A[523] * mat_B[377] +
//             mat_A[524] * mat_B[409] +
//             mat_A[525] * mat_B[441] +
//             mat_A[526] * mat_B[473] +
//             mat_A[527] * mat_B[505] +
//             mat_A[528] * mat_B[537] +
//             mat_A[529] * mat_B[569] +
//             mat_A[530] * mat_B[601] +
//             mat_A[531] * mat_B[633] +
//             mat_A[532] * mat_B[665] +
//             mat_A[533] * mat_B[697] +
//             mat_A[534] * mat_B[729] +
//             mat_A[535] * mat_B[761] +
//             mat_A[536] * mat_B[793] +
//             mat_A[537] * mat_B[825] +
//             mat_A[538] * mat_B[857] +
//             mat_A[539] * mat_B[889] +
//             mat_A[540] * mat_B[921] +
//             mat_A[541] * mat_B[953] +
//             mat_A[542] * mat_B[985] +
//             mat_A[543] * mat_B[1017];
//  mat_C[538] <= 
//             mat_A[512] * mat_B[26] +
//             mat_A[513] * mat_B[58] +
//             mat_A[514] * mat_B[90] +
//             mat_A[515] * mat_B[122] +
//             mat_A[516] * mat_B[154] +
//             mat_A[517] * mat_B[186] +
//             mat_A[518] * mat_B[218] +
//             mat_A[519] * mat_B[250] +
//             mat_A[520] * mat_B[282] +
//             mat_A[521] * mat_B[314] +
//             mat_A[522] * mat_B[346] +
//             mat_A[523] * mat_B[378] +
//             mat_A[524] * mat_B[410] +
//             mat_A[525] * mat_B[442] +
//             mat_A[526] * mat_B[474] +
//             mat_A[527] * mat_B[506] +
//             mat_A[528] * mat_B[538] +
//             mat_A[529] * mat_B[570] +
//             mat_A[530] * mat_B[602] +
//             mat_A[531] * mat_B[634] +
//             mat_A[532] * mat_B[666] +
//             mat_A[533] * mat_B[698] +
//             mat_A[534] * mat_B[730] +
//             mat_A[535] * mat_B[762] +
//             mat_A[536] * mat_B[794] +
//             mat_A[537] * mat_B[826] +
//             mat_A[538] * mat_B[858] +
//             mat_A[539] * mat_B[890] +
//             mat_A[540] * mat_B[922] +
//             mat_A[541] * mat_B[954] +
//             mat_A[542] * mat_B[986] +
//             mat_A[543] * mat_B[1018];
//  mat_C[539] <= 
//             mat_A[512] * mat_B[27] +
//             mat_A[513] * mat_B[59] +
//             mat_A[514] * mat_B[91] +
//             mat_A[515] * mat_B[123] +
//             mat_A[516] * mat_B[155] +
//             mat_A[517] * mat_B[187] +
//             mat_A[518] * mat_B[219] +
//             mat_A[519] * mat_B[251] +
//             mat_A[520] * mat_B[283] +
//             mat_A[521] * mat_B[315] +
//             mat_A[522] * mat_B[347] +
//             mat_A[523] * mat_B[379] +
//             mat_A[524] * mat_B[411] +
//             mat_A[525] * mat_B[443] +
//             mat_A[526] * mat_B[475] +
//             mat_A[527] * mat_B[507] +
//             mat_A[528] * mat_B[539] +
//             mat_A[529] * mat_B[571] +
//             mat_A[530] * mat_B[603] +
//             mat_A[531] * mat_B[635] +
//             mat_A[532] * mat_B[667] +
//             mat_A[533] * mat_B[699] +
//             mat_A[534] * mat_B[731] +
//             mat_A[535] * mat_B[763] +
//             mat_A[536] * mat_B[795] +
//             mat_A[537] * mat_B[827] +
//             mat_A[538] * mat_B[859] +
//             mat_A[539] * mat_B[891] +
//             mat_A[540] * mat_B[923] +
//             mat_A[541] * mat_B[955] +
//             mat_A[542] * mat_B[987] +
//             mat_A[543] * mat_B[1019];
//  mat_C[540] <= 
//             mat_A[512] * mat_B[28] +
//             mat_A[513] * mat_B[60] +
//             mat_A[514] * mat_B[92] +
//             mat_A[515] * mat_B[124] +
//             mat_A[516] * mat_B[156] +
//             mat_A[517] * mat_B[188] +
//             mat_A[518] * mat_B[220] +
//             mat_A[519] * mat_B[252] +
//             mat_A[520] * mat_B[284] +
//             mat_A[521] * mat_B[316] +
//             mat_A[522] * mat_B[348] +
//             mat_A[523] * mat_B[380] +
//             mat_A[524] * mat_B[412] +
//             mat_A[525] * mat_B[444] +
//             mat_A[526] * mat_B[476] +
//             mat_A[527] * mat_B[508] +
//             mat_A[528] * mat_B[540] +
//             mat_A[529] * mat_B[572] +
//             mat_A[530] * mat_B[604] +
//             mat_A[531] * mat_B[636] +
//             mat_A[532] * mat_B[668] +
//             mat_A[533] * mat_B[700] +
//             mat_A[534] * mat_B[732] +
//             mat_A[535] * mat_B[764] +
//             mat_A[536] * mat_B[796] +
//             mat_A[537] * mat_B[828] +
//             mat_A[538] * mat_B[860] +
//             mat_A[539] * mat_B[892] +
//             mat_A[540] * mat_B[924] +
//             mat_A[541] * mat_B[956] +
//             mat_A[542] * mat_B[988] +
//             mat_A[543] * mat_B[1020];
//  mat_C[541] <= 
//             mat_A[512] * mat_B[29] +
//             mat_A[513] * mat_B[61] +
//             mat_A[514] * mat_B[93] +
//             mat_A[515] * mat_B[125] +
//             mat_A[516] * mat_B[157] +
//             mat_A[517] * mat_B[189] +
//             mat_A[518] * mat_B[221] +
//             mat_A[519] * mat_B[253] +
//             mat_A[520] * mat_B[285] +
//             mat_A[521] * mat_B[317] +
//             mat_A[522] * mat_B[349] +
//             mat_A[523] * mat_B[381] +
//             mat_A[524] * mat_B[413] +
//             mat_A[525] * mat_B[445] +
//             mat_A[526] * mat_B[477] +
//             mat_A[527] * mat_B[509] +
//             mat_A[528] * mat_B[541] +
//             mat_A[529] * mat_B[573] +
//             mat_A[530] * mat_B[605] +
//             mat_A[531] * mat_B[637] +
//             mat_A[532] * mat_B[669] +
//             mat_A[533] * mat_B[701] +
//             mat_A[534] * mat_B[733] +
//             mat_A[535] * mat_B[765] +
//             mat_A[536] * mat_B[797] +
//             mat_A[537] * mat_B[829] +
//             mat_A[538] * mat_B[861] +
//             mat_A[539] * mat_B[893] +
//             mat_A[540] * mat_B[925] +
//             mat_A[541] * mat_B[957] +
//             mat_A[542] * mat_B[989] +
//             mat_A[543] * mat_B[1021];
//  mat_C[542] <= 
//             mat_A[512] * mat_B[30] +
//             mat_A[513] * mat_B[62] +
//             mat_A[514] * mat_B[94] +
//             mat_A[515] * mat_B[126] +
//             mat_A[516] * mat_B[158] +
//             mat_A[517] * mat_B[190] +
//             mat_A[518] * mat_B[222] +
//             mat_A[519] * mat_B[254] +
//             mat_A[520] * mat_B[286] +
//             mat_A[521] * mat_B[318] +
//             mat_A[522] * mat_B[350] +
//             mat_A[523] * mat_B[382] +
//             mat_A[524] * mat_B[414] +
//             mat_A[525] * mat_B[446] +
//             mat_A[526] * mat_B[478] +
//             mat_A[527] * mat_B[510] +
//             mat_A[528] * mat_B[542] +
//             mat_A[529] * mat_B[574] +
//             mat_A[530] * mat_B[606] +
//             mat_A[531] * mat_B[638] +
//             mat_A[532] * mat_B[670] +
//             mat_A[533] * mat_B[702] +
//             mat_A[534] * mat_B[734] +
//             mat_A[535] * mat_B[766] +
//             mat_A[536] * mat_B[798] +
//             mat_A[537] * mat_B[830] +
//             mat_A[538] * mat_B[862] +
//             mat_A[539] * mat_B[894] +
//             mat_A[540] * mat_B[926] +
//             mat_A[541] * mat_B[958] +
//             mat_A[542] * mat_B[990] +
//             mat_A[543] * mat_B[1022];
//  mat_C[543] <= 
//             mat_A[512] * mat_B[31] +
//             mat_A[513] * mat_B[63] +
//             mat_A[514] * mat_B[95] +
//             mat_A[515] * mat_B[127] +
//             mat_A[516] * mat_B[159] +
//             mat_A[517] * mat_B[191] +
//             mat_A[518] * mat_B[223] +
//             mat_A[519] * mat_B[255] +
//             mat_A[520] * mat_B[287] +
//             mat_A[521] * mat_B[319] +
//             mat_A[522] * mat_B[351] +
//             mat_A[523] * mat_B[383] +
//             mat_A[524] * mat_B[415] +
//             mat_A[525] * mat_B[447] +
//             mat_A[526] * mat_B[479] +
//             mat_A[527] * mat_B[511] +
//             mat_A[528] * mat_B[543] +
//             mat_A[529] * mat_B[575] +
//             mat_A[530] * mat_B[607] +
//             mat_A[531] * mat_B[639] +
//             mat_A[532] * mat_B[671] +
//             mat_A[533] * mat_B[703] +
//             mat_A[534] * mat_B[735] +
//             mat_A[535] * mat_B[767] +
//             mat_A[536] * mat_B[799] +
//             mat_A[537] * mat_B[831] +
//             mat_A[538] * mat_B[863] +
//             mat_A[539] * mat_B[895] +
//             mat_A[540] * mat_B[927] +
//             mat_A[541] * mat_B[959] +
//             mat_A[542] * mat_B[991] +
//             mat_A[543] * mat_B[1023];
//  mat_C[544] <= 
//             mat_A[544] * mat_B[0] +
//             mat_A[545] * mat_B[32] +
//             mat_A[546] * mat_B[64] +
//             mat_A[547] * mat_B[96] +
//             mat_A[548] * mat_B[128] +
//             mat_A[549] * mat_B[160] +
//             mat_A[550] * mat_B[192] +
//             mat_A[551] * mat_B[224] +
//             mat_A[552] * mat_B[256] +
//             mat_A[553] * mat_B[288] +
//             mat_A[554] * mat_B[320] +
//             mat_A[555] * mat_B[352] +
//             mat_A[556] * mat_B[384] +
//             mat_A[557] * mat_B[416] +
//             mat_A[558] * mat_B[448] +
//             mat_A[559] * mat_B[480] +
//             mat_A[560] * mat_B[512] +
//             mat_A[561] * mat_B[544] +
//             mat_A[562] * mat_B[576] +
//             mat_A[563] * mat_B[608] +
//             mat_A[564] * mat_B[640] +
//             mat_A[565] * mat_B[672] +
//             mat_A[566] * mat_B[704] +
//             mat_A[567] * mat_B[736] +
//             mat_A[568] * mat_B[768] +
//             mat_A[569] * mat_B[800] +
//             mat_A[570] * mat_B[832] +
//             mat_A[571] * mat_B[864] +
//             mat_A[572] * mat_B[896] +
//             mat_A[573] * mat_B[928] +
//             mat_A[574] * mat_B[960] +
//             mat_A[575] * mat_B[992];
//  mat_C[545] <= 
//             mat_A[544] * mat_B[1] +
//             mat_A[545] * mat_B[33] +
//             mat_A[546] * mat_B[65] +
//             mat_A[547] * mat_B[97] +
//             mat_A[548] * mat_B[129] +
//             mat_A[549] * mat_B[161] +
//             mat_A[550] * mat_B[193] +
//             mat_A[551] * mat_B[225] +
//             mat_A[552] * mat_B[257] +
//             mat_A[553] * mat_B[289] +
//             mat_A[554] * mat_B[321] +
//             mat_A[555] * mat_B[353] +
//             mat_A[556] * mat_B[385] +
//             mat_A[557] * mat_B[417] +
//             mat_A[558] * mat_B[449] +
//             mat_A[559] * mat_B[481] +
//             mat_A[560] * mat_B[513] +
//             mat_A[561] * mat_B[545] +
//             mat_A[562] * mat_B[577] +
//             mat_A[563] * mat_B[609] +
//             mat_A[564] * mat_B[641] +
//             mat_A[565] * mat_B[673] +
//             mat_A[566] * mat_B[705] +
//             mat_A[567] * mat_B[737] +
//             mat_A[568] * mat_B[769] +
//             mat_A[569] * mat_B[801] +
//             mat_A[570] * mat_B[833] +
//             mat_A[571] * mat_B[865] +
//             mat_A[572] * mat_B[897] +
//             mat_A[573] * mat_B[929] +
//             mat_A[574] * mat_B[961] +
//             mat_A[575] * mat_B[993];
//  mat_C[546] <= 
//             mat_A[544] * mat_B[2] +
//             mat_A[545] * mat_B[34] +
//             mat_A[546] * mat_B[66] +
//             mat_A[547] * mat_B[98] +
//             mat_A[548] * mat_B[130] +
//             mat_A[549] * mat_B[162] +
//             mat_A[550] * mat_B[194] +
//             mat_A[551] * mat_B[226] +
//             mat_A[552] * mat_B[258] +
//             mat_A[553] * mat_B[290] +
//             mat_A[554] * mat_B[322] +
//             mat_A[555] * mat_B[354] +
//             mat_A[556] * mat_B[386] +
//             mat_A[557] * mat_B[418] +
//             mat_A[558] * mat_B[450] +
//             mat_A[559] * mat_B[482] +
//             mat_A[560] * mat_B[514] +
//             mat_A[561] * mat_B[546] +
//             mat_A[562] * mat_B[578] +
//             mat_A[563] * mat_B[610] +
//             mat_A[564] * mat_B[642] +
//             mat_A[565] * mat_B[674] +
//             mat_A[566] * mat_B[706] +
//             mat_A[567] * mat_B[738] +
//             mat_A[568] * mat_B[770] +
//             mat_A[569] * mat_B[802] +
//             mat_A[570] * mat_B[834] +
//             mat_A[571] * mat_B[866] +
//             mat_A[572] * mat_B[898] +
//             mat_A[573] * mat_B[930] +
//             mat_A[574] * mat_B[962] +
//             mat_A[575] * mat_B[994];
//  mat_C[547] <= 
//             mat_A[544] * mat_B[3] +
//             mat_A[545] * mat_B[35] +
//             mat_A[546] * mat_B[67] +
//             mat_A[547] * mat_B[99] +
//             mat_A[548] * mat_B[131] +
//             mat_A[549] * mat_B[163] +
//             mat_A[550] * mat_B[195] +
//             mat_A[551] * mat_B[227] +
//             mat_A[552] * mat_B[259] +
//             mat_A[553] * mat_B[291] +
//             mat_A[554] * mat_B[323] +
//             mat_A[555] * mat_B[355] +
//             mat_A[556] * mat_B[387] +
//             mat_A[557] * mat_B[419] +
//             mat_A[558] * mat_B[451] +
//             mat_A[559] * mat_B[483] +
//             mat_A[560] * mat_B[515] +
//             mat_A[561] * mat_B[547] +
//             mat_A[562] * mat_B[579] +
//             mat_A[563] * mat_B[611] +
//             mat_A[564] * mat_B[643] +
//             mat_A[565] * mat_B[675] +
//             mat_A[566] * mat_B[707] +
//             mat_A[567] * mat_B[739] +
//             mat_A[568] * mat_B[771] +
//             mat_A[569] * mat_B[803] +
//             mat_A[570] * mat_B[835] +
//             mat_A[571] * mat_B[867] +
//             mat_A[572] * mat_B[899] +
//             mat_A[573] * mat_B[931] +
//             mat_A[574] * mat_B[963] +
//             mat_A[575] * mat_B[995];
//  mat_C[548] <= 
//             mat_A[544] * mat_B[4] +
//             mat_A[545] * mat_B[36] +
//             mat_A[546] * mat_B[68] +
//             mat_A[547] * mat_B[100] +
//             mat_A[548] * mat_B[132] +
//             mat_A[549] * mat_B[164] +
//             mat_A[550] * mat_B[196] +
//             mat_A[551] * mat_B[228] +
//             mat_A[552] * mat_B[260] +
//             mat_A[553] * mat_B[292] +
//             mat_A[554] * mat_B[324] +
//             mat_A[555] * mat_B[356] +
//             mat_A[556] * mat_B[388] +
//             mat_A[557] * mat_B[420] +
//             mat_A[558] * mat_B[452] +
//             mat_A[559] * mat_B[484] +
//             mat_A[560] * mat_B[516] +
//             mat_A[561] * mat_B[548] +
//             mat_A[562] * mat_B[580] +
//             mat_A[563] * mat_B[612] +
//             mat_A[564] * mat_B[644] +
//             mat_A[565] * mat_B[676] +
//             mat_A[566] * mat_B[708] +
//             mat_A[567] * mat_B[740] +
//             mat_A[568] * mat_B[772] +
//             mat_A[569] * mat_B[804] +
//             mat_A[570] * mat_B[836] +
//             mat_A[571] * mat_B[868] +
//             mat_A[572] * mat_B[900] +
//             mat_A[573] * mat_B[932] +
//             mat_A[574] * mat_B[964] +
//             mat_A[575] * mat_B[996];
//  mat_C[549] <= 
//             mat_A[544] * mat_B[5] +
//             mat_A[545] * mat_B[37] +
//             mat_A[546] * mat_B[69] +
//             mat_A[547] * mat_B[101] +
//             mat_A[548] * mat_B[133] +
//             mat_A[549] * mat_B[165] +
//             mat_A[550] * mat_B[197] +
//             mat_A[551] * mat_B[229] +
//             mat_A[552] * mat_B[261] +
//             mat_A[553] * mat_B[293] +
//             mat_A[554] * mat_B[325] +
//             mat_A[555] * mat_B[357] +
//             mat_A[556] * mat_B[389] +
//             mat_A[557] * mat_B[421] +
//             mat_A[558] * mat_B[453] +
//             mat_A[559] * mat_B[485] +
//             mat_A[560] * mat_B[517] +
//             mat_A[561] * mat_B[549] +
//             mat_A[562] * mat_B[581] +
//             mat_A[563] * mat_B[613] +
//             mat_A[564] * mat_B[645] +
//             mat_A[565] * mat_B[677] +
//             mat_A[566] * mat_B[709] +
//             mat_A[567] * mat_B[741] +
//             mat_A[568] * mat_B[773] +
//             mat_A[569] * mat_B[805] +
//             mat_A[570] * mat_B[837] +
//             mat_A[571] * mat_B[869] +
//             mat_A[572] * mat_B[901] +
//             mat_A[573] * mat_B[933] +
//             mat_A[574] * mat_B[965] +
//             mat_A[575] * mat_B[997];
//  mat_C[550] <= 
//             mat_A[544] * mat_B[6] +
//             mat_A[545] * mat_B[38] +
//             mat_A[546] * mat_B[70] +
//             mat_A[547] * mat_B[102] +
//             mat_A[548] * mat_B[134] +
//             mat_A[549] * mat_B[166] +
//             mat_A[550] * mat_B[198] +
//             mat_A[551] * mat_B[230] +
//             mat_A[552] * mat_B[262] +
//             mat_A[553] * mat_B[294] +
//             mat_A[554] * mat_B[326] +
//             mat_A[555] * mat_B[358] +
//             mat_A[556] * mat_B[390] +
//             mat_A[557] * mat_B[422] +
//             mat_A[558] * mat_B[454] +
//             mat_A[559] * mat_B[486] +
//             mat_A[560] * mat_B[518] +
//             mat_A[561] * mat_B[550] +
//             mat_A[562] * mat_B[582] +
//             mat_A[563] * mat_B[614] +
//             mat_A[564] * mat_B[646] +
//             mat_A[565] * mat_B[678] +
//             mat_A[566] * mat_B[710] +
//             mat_A[567] * mat_B[742] +
//             mat_A[568] * mat_B[774] +
//             mat_A[569] * mat_B[806] +
//             mat_A[570] * mat_B[838] +
//             mat_A[571] * mat_B[870] +
//             mat_A[572] * mat_B[902] +
//             mat_A[573] * mat_B[934] +
//             mat_A[574] * mat_B[966] +
//             mat_A[575] * mat_B[998];
//  mat_C[551] <= 
//             mat_A[544] * mat_B[7] +
//             mat_A[545] * mat_B[39] +
//             mat_A[546] * mat_B[71] +
//             mat_A[547] * mat_B[103] +
//             mat_A[548] * mat_B[135] +
//             mat_A[549] * mat_B[167] +
//             mat_A[550] * mat_B[199] +
//             mat_A[551] * mat_B[231] +
//             mat_A[552] * mat_B[263] +
//             mat_A[553] * mat_B[295] +
//             mat_A[554] * mat_B[327] +
//             mat_A[555] * mat_B[359] +
//             mat_A[556] * mat_B[391] +
//             mat_A[557] * mat_B[423] +
//             mat_A[558] * mat_B[455] +
//             mat_A[559] * mat_B[487] +
//             mat_A[560] * mat_B[519] +
//             mat_A[561] * mat_B[551] +
//             mat_A[562] * mat_B[583] +
//             mat_A[563] * mat_B[615] +
//             mat_A[564] * mat_B[647] +
//             mat_A[565] * mat_B[679] +
//             mat_A[566] * mat_B[711] +
//             mat_A[567] * mat_B[743] +
//             mat_A[568] * mat_B[775] +
//             mat_A[569] * mat_B[807] +
//             mat_A[570] * mat_B[839] +
//             mat_A[571] * mat_B[871] +
//             mat_A[572] * mat_B[903] +
//             mat_A[573] * mat_B[935] +
//             mat_A[574] * mat_B[967] +
//             mat_A[575] * mat_B[999];
//  mat_C[552] <= 
//             mat_A[544] * mat_B[8] +
//             mat_A[545] * mat_B[40] +
//             mat_A[546] * mat_B[72] +
//             mat_A[547] * mat_B[104] +
//             mat_A[548] * mat_B[136] +
//             mat_A[549] * mat_B[168] +
//             mat_A[550] * mat_B[200] +
//             mat_A[551] * mat_B[232] +
//             mat_A[552] * mat_B[264] +
//             mat_A[553] * mat_B[296] +
//             mat_A[554] * mat_B[328] +
//             mat_A[555] * mat_B[360] +
//             mat_A[556] * mat_B[392] +
//             mat_A[557] * mat_B[424] +
//             mat_A[558] * mat_B[456] +
//             mat_A[559] * mat_B[488] +
//             mat_A[560] * mat_B[520] +
//             mat_A[561] * mat_B[552] +
//             mat_A[562] * mat_B[584] +
//             mat_A[563] * mat_B[616] +
//             mat_A[564] * mat_B[648] +
//             mat_A[565] * mat_B[680] +
//             mat_A[566] * mat_B[712] +
//             mat_A[567] * mat_B[744] +
//             mat_A[568] * mat_B[776] +
//             mat_A[569] * mat_B[808] +
//             mat_A[570] * mat_B[840] +
//             mat_A[571] * mat_B[872] +
//             mat_A[572] * mat_B[904] +
//             mat_A[573] * mat_B[936] +
//             mat_A[574] * mat_B[968] +
//             mat_A[575] * mat_B[1000];
//  mat_C[553] <= 
//             mat_A[544] * mat_B[9] +
//             mat_A[545] * mat_B[41] +
//             mat_A[546] * mat_B[73] +
//             mat_A[547] * mat_B[105] +
//             mat_A[548] * mat_B[137] +
//             mat_A[549] * mat_B[169] +
//             mat_A[550] * mat_B[201] +
//             mat_A[551] * mat_B[233] +
//             mat_A[552] * mat_B[265] +
//             mat_A[553] * mat_B[297] +
//             mat_A[554] * mat_B[329] +
//             mat_A[555] * mat_B[361] +
//             mat_A[556] * mat_B[393] +
//             mat_A[557] * mat_B[425] +
//             mat_A[558] * mat_B[457] +
//             mat_A[559] * mat_B[489] +
//             mat_A[560] * mat_B[521] +
//             mat_A[561] * mat_B[553] +
//             mat_A[562] * mat_B[585] +
//             mat_A[563] * mat_B[617] +
//             mat_A[564] * mat_B[649] +
//             mat_A[565] * mat_B[681] +
//             mat_A[566] * mat_B[713] +
//             mat_A[567] * mat_B[745] +
//             mat_A[568] * mat_B[777] +
//             mat_A[569] * mat_B[809] +
//             mat_A[570] * mat_B[841] +
//             mat_A[571] * mat_B[873] +
//             mat_A[572] * mat_B[905] +
//             mat_A[573] * mat_B[937] +
//             mat_A[574] * mat_B[969] +
//             mat_A[575] * mat_B[1001];
//  mat_C[554] <= 
//             mat_A[544] * mat_B[10] +
//             mat_A[545] * mat_B[42] +
//             mat_A[546] * mat_B[74] +
//             mat_A[547] * mat_B[106] +
//             mat_A[548] * mat_B[138] +
//             mat_A[549] * mat_B[170] +
//             mat_A[550] * mat_B[202] +
//             mat_A[551] * mat_B[234] +
//             mat_A[552] * mat_B[266] +
//             mat_A[553] * mat_B[298] +
//             mat_A[554] * mat_B[330] +
//             mat_A[555] * mat_B[362] +
//             mat_A[556] * mat_B[394] +
//             mat_A[557] * mat_B[426] +
//             mat_A[558] * mat_B[458] +
//             mat_A[559] * mat_B[490] +
//             mat_A[560] * mat_B[522] +
//             mat_A[561] * mat_B[554] +
//             mat_A[562] * mat_B[586] +
//             mat_A[563] * mat_B[618] +
//             mat_A[564] * mat_B[650] +
//             mat_A[565] * mat_B[682] +
//             mat_A[566] * mat_B[714] +
//             mat_A[567] * mat_B[746] +
//             mat_A[568] * mat_B[778] +
//             mat_A[569] * mat_B[810] +
//             mat_A[570] * mat_B[842] +
//             mat_A[571] * mat_B[874] +
//             mat_A[572] * mat_B[906] +
//             mat_A[573] * mat_B[938] +
//             mat_A[574] * mat_B[970] +
//             mat_A[575] * mat_B[1002];
//  mat_C[555] <= 
//             mat_A[544] * mat_B[11] +
//             mat_A[545] * mat_B[43] +
//             mat_A[546] * mat_B[75] +
//             mat_A[547] * mat_B[107] +
//             mat_A[548] * mat_B[139] +
//             mat_A[549] * mat_B[171] +
//             mat_A[550] * mat_B[203] +
//             mat_A[551] * mat_B[235] +
//             mat_A[552] * mat_B[267] +
//             mat_A[553] * mat_B[299] +
//             mat_A[554] * mat_B[331] +
//             mat_A[555] * mat_B[363] +
//             mat_A[556] * mat_B[395] +
//             mat_A[557] * mat_B[427] +
//             mat_A[558] * mat_B[459] +
//             mat_A[559] * mat_B[491] +
//             mat_A[560] * mat_B[523] +
//             mat_A[561] * mat_B[555] +
//             mat_A[562] * mat_B[587] +
//             mat_A[563] * mat_B[619] +
//             mat_A[564] * mat_B[651] +
//             mat_A[565] * mat_B[683] +
//             mat_A[566] * mat_B[715] +
//             mat_A[567] * mat_B[747] +
//             mat_A[568] * mat_B[779] +
//             mat_A[569] * mat_B[811] +
//             mat_A[570] * mat_B[843] +
//             mat_A[571] * mat_B[875] +
//             mat_A[572] * mat_B[907] +
//             mat_A[573] * mat_B[939] +
//             mat_A[574] * mat_B[971] +
//             mat_A[575] * mat_B[1003];
//  mat_C[556] <= 
//             mat_A[544] * mat_B[12] +
//             mat_A[545] * mat_B[44] +
//             mat_A[546] * mat_B[76] +
//             mat_A[547] * mat_B[108] +
//             mat_A[548] * mat_B[140] +
//             mat_A[549] * mat_B[172] +
//             mat_A[550] * mat_B[204] +
//             mat_A[551] * mat_B[236] +
//             mat_A[552] * mat_B[268] +
//             mat_A[553] * mat_B[300] +
//             mat_A[554] * mat_B[332] +
//             mat_A[555] * mat_B[364] +
//             mat_A[556] * mat_B[396] +
//             mat_A[557] * mat_B[428] +
//             mat_A[558] * mat_B[460] +
//             mat_A[559] * mat_B[492] +
//             mat_A[560] * mat_B[524] +
//             mat_A[561] * mat_B[556] +
//             mat_A[562] * mat_B[588] +
//             mat_A[563] * mat_B[620] +
//             mat_A[564] * mat_B[652] +
//             mat_A[565] * mat_B[684] +
//             mat_A[566] * mat_B[716] +
//             mat_A[567] * mat_B[748] +
//             mat_A[568] * mat_B[780] +
//             mat_A[569] * mat_B[812] +
//             mat_A[570] * mat_B[844] +
//             mat_A[571] * mat_B[876] +
//             mat_A[572] * mat_B[908] +
//             mat_A[573] * mat_B[940] +
//             mat_A[574] * mat_B[972] +
//             mat_A[575] * mat_B[1004];
//  mat_C[557] <= 
//             mat_A[544] * mat_B[13] +
//             mat_A[545] * mat_B[45] +
//             mat_A[546] * mat_B[77] +
//             mat_A[547] * mat_B[109] +
//             mat_A[548] * mat_B[141] +
//             mat_A[549] * mat_B[173] +
//             mat_A[550] * mat_B[205] +
//             mat_A[551] * mat_B[237] +
//             mat_A[552] * mat_B[269] +
//             mat_A[553] * mat_B[301] +
//             mat_A[554] * mat_B[333] +
//             mat_A[555] * mat_B[365] +
//             mat_A[556] * mat_B[397] +
//             mat_A[557] * mat_B[429] +
//             mat_A[558] * mat_B[461] +
//             mat_A[559] * mat_B[493] +
//             mat_A[560] * mat_B[525] +
//             mat_A[561] * mat_B[557] +
//             mat_A[562] * mat_B[589] +
//             mat_A[563] * mat_B[621] +
//             mat_A[564] * mat_B[653] +
//             mat_A[565] * mat_B[685] +
//             mat_A[566] * mat_B[717] +
//             mat_A[567] * mat_B[749] +
//             mat_A[568] * mat_B[781] +
//             mat_A[569] * mat_B[813] +
//             mat_A[570] * mat_B[845] +
//             mat_A[571] * mat_B[877] +
//             mat_A[572] * mat_B[909] +
//             mat_A[573] * mat_B[941] +
//             mat_A[574] * mat_B[973] +
//             mat_A[575] * mat_B[1005];
//  mat_C[558] <= 
//             mat_A[544] * mat_B[14] +
//             mat_A[545] * mat_B[46] +
//             mat_A[546] * mat_B[78] +
//             mat_A[547] * mat_B[110] +
//             mat_A[548] * mat_B[142] +
//             mat_A[549] * mat_B[174] +
//             mat_A[550] * mat_B[206] +
//             mat_A[551] * mat_B[238] +
//             mat_A[552] * mat_B[270] +
//             mat_A[553] * mat_B[302] +
//             mat_A[554] * mat_B[334] +
//             mat_A[555] * mat_B[366] +
//             mat_A[556] * mat_B[398] +
//             mat_A[557] * mat_B[430] +
//             mat_A[558] * mat_B[462] +
//             mat_A[559] * mat_B[494] +
//             mat_A[560] * mat_B[526] +
//             mat_A[561] * mat_B[558] +
//             mat_A[562] * mat_B[590] +
//             mat_A[563] * mat_B[622] +
//             mat_A[564] * mat_B[654] +
//             mat_A[565] * mat_B[686] +
//             mat_A[566] * mat_B[718] +
//             mat_A[567] * mat_B[750] +
//             mat_A[568] * mat_B[782] +
//             mat_A[569] * mat_B[814] +
//             mat_A[570] * mat_B[846] +
//             mat_A[571] * mat_B[878] +
//             mat_A[572] * mat_B[910] +
//             mat_A[573] * mat_B[942] +
//             mat_A[574] * mat_B[974] +
//             mat_A[575] * mat_B[1006];
//  mat_C[559] <= 
//             mat_A[544] * mat_B[15] +
//             mat_A[545] * mat_B[47] +
//             mat_A[546] * mat_B[79] +
//             mat_A[547] * mat_B[111] +
//             mat_A[548] * mat_B[143] +
//             mat_A[549] * mat_B[175] +
//             mat_A[550] * mat_B[207] +
//             mat_A[551] * mat_B[239] +
//             mat_A[552] * mat_B[271] +
//             mat_A[553] * mat_B[303] +
//             mat_A[554] * mat_B[335] +
//             mat_A[555] * mat_B[367] +
//             mat_A[556] * mat_B[399] +
//             mat_A[557] * mat_B[431] +
//             mat_A[558] * mat_B[463] +
//             mat_A[559] * mat_B[495] +
//             mat_A[560] * mat_B[527] +
//             mat_A[561] * mat_B[559] +
//             mat_A[562] * mat_B[591] +
//             mat_A[563] * mat_B[623] +
//             mat_A[564] * mat_B[655] +
//             mat_A[565] * mat_B[687] +
//             mat_A[566] * mat_B[719] +
//             mat_A[567] * mat_B[751] +
//             mat_A[568] * mat_B[783] +
//             mat_A[569] * mat_B[815] +
//             mat_A[570] * mat_B[847] +
//             mat_A[571] * mat_B[879] +
//             mat_A[572] * mat_B[911] +
//             mat_A[573] * mat_B[943] +
//             mat_A[574] * mat_B[975] +
//             mat_A[575] * mat_B[1007];
//  mat_C[560] <= 
//             mat_A[544] * mat_B[16] +
//             mat_A[545] * mat_B[48] +
//             mat_A[546] * mat_B[80] +
//             mat_A[547] * mat_B[112] +
//             mat_A[548] * mat_B[144] +
//             mat_A[549] * mat_B[176] +
//             mat_A[550] * mat_B[208] +
//             mat_A[551] * mat_B[240] +
//             mat_A[552] * mat_B[272] +
//             mat_A[553] * mat_B[304] +
//             mat_A[554] * mat_B[336] +
//             mat_A[555] * mat_B[368] +
//             mat_A[556] * mat_B[400] +
//             mat_A[557] * mat_B[432] +
//             mat_A[558] * mat_B[464] +
//             mat_A[559] * mat_B[496] +
//             mat_A[560] * mat_B[528] +
//             mat_A[561] * mat_B[560] +
//             mat_A[562] * mat_B[592] +
//             mat_A[563] * mat_B[624] +
//             mat_A[564] * mat_B[656] +
//             mat_A[565] * mat_B[688] +
//             mat_A[566] * mat_B[720] +
//             mat_A[567] * mat_B[752] +
//             mat_A[568] * mat_B[784] +
//             mat_A[569] * mat_B[816] +
//             mat_A[570] * mat_B[848] +
//             mat_A[571] * mat_B[880] +
//             mat_A[572] * mat_B[912] +
//             mat_A[573] * mat_B[944] +
//             mat_A[574] * mat_B[976] +
//             mat_A[575] * mat_B[1008];
//  mat_C[561] <= 
//             mat_A[544] * mat_B[17] +
//             mat_A[545] * mat_B[49] +
//             mat_A[546] * mat_B[81] +
//             mat_A[547] * mat_B[113] +
//             mat_A[548] * mat_B[145] +
//             mat_A[549] * mat_B[177] +
//             mat_A[550] * mat_B[209] +
//             mat_A[551] * mat_B[241] +
//             mat_A[552] * mat_B[273] +
//             mat_A[553] * mat_B[305] +
//             mat_A[554] * mat_B[337] +
//             mat_A[555] * mat_B[369] +
//             mat_A[556] * mat_B[401] +
//             mat_A[557] * mat_B[433] +
//             mat_A[558] * mat_B[465] +
//             mat_A[559] * mat_B[497] +
//             mat_A[560] * mat_B[529] +
//             mat_A[561] * mat_B[561] +
//             mat_A[562] * mat_B[593] +
//             mat_A[563] * mat_B[625] +
//             mat_A[564] * mat_B[657] +
//             mat_A[565] * mat_B[689] +
//             mat_A[566] * mat_B[721] +
//             mat_A[567] * mat_B[753] +
//             mat_A[568] * mat_B[785] +
//             mat_A[569] * mat_B[817] +
//             mat_A[570] * mat_B[849] +
//             mat_A[571] * mat_B[881] +
//             mat_A[572] * mat_B[913] +
//             mat_A[573] * mat_B[945] +
//             mat_A[574] * mat_B[977] +
//             mat_A[575] * mat_B[1009];
//  mat_C[562] <= 
//             mat_A[544] * mat_B[18] +
//             mat_A[545] * mat_B[50] +
//             mat_A[546] * mat_B[82] +
//             mat_A[547] * mat_B[114] +
//             mat_A[548] * mat_B[146] +
//             mat_A[549] * mat_B[178] +
//             mat_A[550] * mat_B[210] +
//             mat_A[551] * mat_B[242] +
//             mat_A[552] * mat_B[274] +
//             mat_A[553] * mat_B[306] +
//             mat_A[554] * mat_B[338] +
//             mat_A[555] * mat_B[370] +
//             mat_A[556] * mat_B[402] +
//             mat_A[557] * mat_B[434] +
//             mat_A[558] * mat_B[466] +
//             mat_A[559] * mat_B[498] +
//             mat_A[560] * mat_B[530] +
//             mat_A[561] * mat_B[562] +
//             mat_A[562] * mat_B[594] +
//             mat_A[563] * mat_B[626] +
//             mat_A[564] * mat_B[658] +
//             mat_A[565] * mat_B[690] +
//             mat_A[566] * mat_B[722] +
//             mat_A[567] * mat_B[754] +
//             mat_A[568] * mat_B[786] +
//             mat_A[569] * mat_B[818] +
//             mat_A[570] * mat_B[850] +
//             mat_A[571] * mat_B[882] +
//             mat_A[572] * mat_B[914] +
//             mat_A[573] * mat_B[946] +
//             mat_A[574] * mat_B[978] +
//             mat_A[575] * mat_B[1010];
//  mat_C[563] <= 
//             mat_A[544] * mat_B[19] +
//             mat_A[545] * mat_B[51] +
//             mat_A[546] * mat_B[83] +
//             mat_A[547] * mat_B[115] +
//             mat_A[548] * mat_B[147] +
//             mat_A[549] * mat_B[179] +
//             mat_A[550] * mat_B[211] +
//             mat_A[551] * mat_B[243] +
//             mat_A[552] * mat_B[275] +
//             mat_A[553] * mat_B[307] +
//             mat_A[554] * mat_B[339] +
//             mat_A[555] * mat_B[371] +
//             mat_A[556] * mat_B[403] +
//             mat_A[557] * mat_B[435] +
//             mat_A[558] * mat_B[467] +
//             mat_A[559] * mat_B[499] +
//             mat_A[560] * mat_B[531] +
//             mat_A[561] * mat_B[563] +
//             mat_A[562] * mat_B[595] +
//             mat_A[563] * mat_B[627] +
//             mat_A[564] * mat_B[659] +
//             mat_A[565] * mat_B[691] +
//             mat_A[566] * mat_B[723] +
//             mat_A[567] * mat_B[755] +
//             mat_A[568] * mat_B[787] +
//             mat_A[569] * mat_B[819] +
//             mat_A[570] * mat_B[851] +
//             mat_A[571] * mat_B[883] +
//             mat_A[572] * mat_B[915] +
//             mat_A[573] * mat_B[947] +
//             mat_A[574] * mat_B[979] +
//             mat_A[575] * mat_B[1011];
//  mat_C[564] <= 
//             mat_A[544] * mat_B[20] +
//             mat_A[545] * mat_B[52] +
//             mat_A[546] * mat_B[84] +
//             mat_A[547] * mat_B[116] +
//             mat_A[548] * mat_B[148] +
//             mat_A[549] * mat_B[180] +
//             mat_A[550] * mat_B[212] +
//             mat_A[551] * mat_B[244] +
//             mat_A[552] * mat_B[276] +
//             mat_A[553] * mat_B[308] +
//             mat_A[554] * mat_B[340] +
//             mat_A[555] * mat_B[372] +
//             mat_A[556] * mat_B[404] +
//             mat_A[557] * mat_B[436] +
//             mat_A[558] * mat_B[468] +
//             mat_A[559] * mat_B[500] +
//             mat_A[560] * mat_B[532] +
//             mat_A[561] * mat_B[564] +
//             mat_A[562] * mat_B[596] +
//             mat_A[563] * mat_B[628] +
//             mat_A[564] * mat_B[660] +
//             mat_A[565] * mat_B[692] +
//             mat_A[566] * mat_B[724] +
//             mat_A[567] * mat_B[756] +
//             mat_A[568] * mat_B[788] +
//             mat_A[569] * mat_B[820] +
//             mat_A[570] * mat_B[852] +
//             mat_A[571] * mat_B[884] +
//             mat_A[572] * mat_B[916] +
//             mat_A[573] * mat_B[948] +
//             mat_A[574] * mat_B[980] +
//             mat_A[575] * mat_B[1012];
//  mat_C[565] <= 
//             mat_A[544] * mat_B[21] +
//             mat_A[545] * mat_B[53] +
//             mat_A[546] * mat_B[85] +
//             mat_A[547] * mat_B[117] +
//             mat_A[548] * mat_B[149] +
//             mat_A[549] * mat_B[181] +
//             mat_A[550] * mat_B[213] +
//             mat_A[551] * mat_B[245] +
//             mat_A[552] * mat_B[277] +
//             mat_A[553] * mat_B[309] +
//             mat_A[554] * mat_B[341] +
//             mat_A[555] * mat_B[373] +
//             mat_A[556] * mat_B[405] +
//             mat_A[557] * mat_B[437] +
//             mat_A[558] * mat_B[469] +
//             mat_A[559] * mat_B[501] +
//             mat_A[560] * mat_B[533] +
//             mat_A[561] * mat_B[565] +
//             mat_A[562] * mat_B[597] +
//             mat_A[563] * mat_B[629] +
//             mat_A[564] * mat_B[661] +
//             mat_A[565] * mat_B[693] +
//             mat_A[566] * mat_B[725] +
//             mat_A[567] * mat_B[757] +
//             mat_A[568] * mat_B[789] +
//             mat_A[569] * mat_B[821] +
//             mat_A[570] * mat_B[853] +
//             mat_A[571] * mat_B[885] +
//             mat_A[572] * mat_B[917] +
//             mat_A[573] * mat_B[949] +
//             mat_A[574] * mat_B[981] +
//             mat_A[575] * mat_B[1013];
//  mat_C[566] <= 
//             mat_A[544] * mat_B[22] +
//             mat_A[545] * mat_B[54] +
//             mat_A[546] * mat_B[86] +
//             mat_A[547] * mat_B[118] +
//             mat_A[548] * mat_B[150] +
//             mat_A[549] * mat_B[182] +
//             mat_A[550] * mat_B[214] +
//             mat_A[551] * mat_B[246] +
//             mat_A[552] * mat_B[278] +
//             mat_A[553] * mat_B[310] +
//             mat_A[554] * mat_B[342] +
//             mat_A[555] * mat_B[374] +
//             mat_A[556] * mat_B[406] +
//             mat_A[557] * mat_B[438] +
//             mat_A[558] * mat_B[470] +
//             mat_A[559] * mat_B[502] +
//             mat_A[560] * mat_B[534] +
//             mat_A[561] * mat_B[566] +
//             mat_A[562] * mat_B[598] +
//             mat_A[563] * mat_B[630] +
//             mat_A[564] * mat_B[662] +
//             mat_A[565] * mat_B[694] +
//             mat_A[566] * mat_B[726] +
//             mat_A[567] * mat_B[758] +
//             mat_A[568] * mat_B[790] +
//             mat_A[569] * mat_B[822] +
//             mat_A[570] * mat_B[854] +
//             mat_A[571] * mat_B[886] +
//             mat_A[572] * mat_B[918] +
//             mat_A[573] * mat_B[950] +
//             mat_A[574] * mat_B[982] +
//             mat_A[575] * mat_B[1014];
//  mat_C[567] <= 
//             mat_A[544] * mat_B[23] +
//             mat_A[545] * mat_B[55] +
//             mat_A[546] * mat_B[87] +
//             mat_A[547] * mat_B[119] +
//             mat_A[548] * mat_B[151] +
//             mat_A[549] * mat_B[183] +
//             mat_A[550] * mat_B[215] +
//             mat_A[551] * mat_B[247] +
//             mat_A[552] * mat_B[279] +
//             mat_A[553] * mat_B[311] +
//             mat_A[554] * mat_B[343] +
//             mat_A[555] * mat_B[375] +
//             mat_A[556] * mat_B[407] +
//             mat_A[557] * mat_B[439] +
//             mat_A[558] * mat_B[471] +
//             mat_A[559] * mat_B[503] +
//             mat_A[560] * mat_B[535] +
//             mat_A[561] * mat_B[567] +
//             mat_A[562] * mat_B[599] +
//             mat_A[563] * mat_B[631] +
//             mat_A[564] * mat_B[663] +
//             mat_A[565] * mat_B[695] +
//             mat_A[566] * mat_B[727] +
//             mat_A[567] * mat_B[759] +
//             mat_A[568] * mat_B[791] +
//             mat_A[569] * mat_B[823] +
//             mat_A[570] * mat_B[855] +
//             mat_A[571] * mat_B[887] +
//             mat_A[572] * mat_B[919] +
//             mat_A[573] * mat_B[951] +
//             mat_A[574] * mat_B[983] +
//             mat_A[575] * mat_B[1015];
//  mat_C[568] <= 
//             mat_A[544] * mat_B[24] +
//             mat_A[545] * mat_B[56] +
//             mat_A[546] * mat_B[88] +
//             mat_A[547] * mat_B[120] +
//             mat_A[548] * mat_B[152] +
//             mat_A[549] * mat_B[184] +
//             mat_A[550] * mat_B[216] +
//             mat_A[551] * mat_B[248] +
//             mat_A[552] * mat_B[280] +
//             mat_A[553] * mat_B[312] +
//             mat_A[554] * mat_B[344] +
//             mat_A[555] * mat_B[376] +
//             mat_A[556] * mat_B[408] +
//             mat_A[557] * mat_B[440] +
//             mat_A[558] * mat_B[472] +
//             mat_A[559] * mat_B[504] +
//             mat_A[560] * mat_B[536] +
//             mat_A[561] * mat_B[568] +
//             mat_A[562] * mat_B[600] +
//             mat_A[563] * mat_B[632] +
//             mat_A[564] * mat_B[664] +
//             mat_A[565] * mat_B[696] +
//             mat_A[566] * mat_B[728] +
//             mat_A[567] * mat_B[760] +
//             mat_A[568] * mat_B[792] +
//             mat_A[569] * mat_B[824] +
//             mat_A[570] * mat_B[856] +
//             mat_A[571] * mat_B[888] +
//             mat_A[572] * mat_B[920] +
//             mat_A[573] * mat_B[952] +
//             mat_A[574] * mat_B[984] +
//             mat_A[575] * mat_B[1016];
//  mat_C[569] <= 
//             mat_A[544] * mat_B[25] +
//             mat_A[545] * mat_B[57] +
//             mat_A[546] * mat_B[89] +
//             mat_A[547] * mat_B[121] +
//             mat_A[548] * mat_B[153] +
//             mat_A[549] * mat_B[185] +
//             mat_A[550] * mat_B[217] +
//             mat_A[551] * mat_B[249] +
//             mat_A[552] * mat_B[281] +
//             mat_A[553] * mat_B[313] +
//             mat_A[554] * mat_B[345] +
//             mat_A[555] * mat_B[377] +
//             mat_A[556] * mat_B[409] +
//             mat_A[557] * mat_B[441] +
//             mat_A[558] * mat_B[473] +
//             mat_A[559] * mat_B[505] +
//             mat_A[560] * mat_B[537] +
//             mat_A[561] * mat_B[569] +
//             mat_A[562] * mat_B[601] +
//             mat_A[563] * mat_B[633] +
//             mat_A[564] * mat_B[665] +
//             mat_A[565] * mat_B[697] +
//             mat_A[566] * mat_B[729] +
//             mat_A[567] * mat_B[761] +
//             mat_A[568] * mat_B[793] +
//             mat_A[569] * mat_B[825] +
//             mat_A[570] * mat_B[857] +
//             mat_A[571] * mat_B[889] +
//             mat_A[572] * mat_B[921] +
//             mat_A[573] * mat_B[953] +
//             mat_A[574] * mat_B[985] +
//             mat_A[575] * mat_B[1017];
//  mat_C[570] <= 
//             mat_A[544] * mat_B[26] +
//             mat_A[545] * mat_B[58] +
//             mat_A[546] * mat_B[90] +
//             mat_A[547] * mat_B[122] +
//             mat_A[548] * mat_B[154] +
//             mat_A[549] * mat_B[186] +
//             mat_A[550] * mat_B[218] +
//             mat_A[551] * mat_B[250] +
//             mat_A[552] * mat_B[282] +
//             mat_A[553] * mat_B[314] +
//             mat_A[554] * mat_B[346] +
//             mat_A[555] * mat_B[378] +
//             mat_A[556] * mat_B[410] +
//             mat_A[557] * mat_B[442] +
//             mat_A[558] * mat_B[474] +
//             mat_A[559] * mat_B[506] +
//             mat_A[560] * mat_B[538] +
//             mat_A[561] * mat_B[570] +
//             mat_A[562] * mat_B[602] +
//             mat_A[563] * mat_B[634] +
//             mat_A[564] * mat_B[666] +
//             mat_A[565] * mat_B[698] +
//             mat_A[566] * mat_B[730] +
//             mat_A[567] * mat_B[762] +
//             mat_A[568] * mat_B[794] +
//             mat_A[569] * mat_B[826] +
//             mat_A[570] * mat_B[858] +
//             mat_A[571] * mat_B[890] +
//             mat_A[572] * mat_B[922] +
//             mat_A[573] * mat_B[954] +
//             mat_A[574] * mat_B[986] +
//             mat_A[575] * mat_B[1018];
//  mat_C[571] <= 
//             mat_A[544] * mat_B[27] +
//             mat_A[545] * mat_B[59] +
//             mat_A[546] * mat_B[91] +
//             mat_A[547] * mat_B[123] +
//             mat_A[548] * mat_B[155] +
//             mat_A[549] * mat_B[187] +
//             mat_A[550] * mat_B[219] +
//             mat_A[551] * mat_B[251] +
//             mat_A[552] * mat_B[283] +
//             mat_A[553] * mat_B[315] +
//             mat_A[554] * mat_B[347] +
//             mat_A[555] * mat_B[379] +
//             mat_A[556] * mat_B[411] +
//             mat_A[557] * mat_B[443] +
//             mat_A[558] * mat_B[475] +
//             mat_A[559] * mat_B[507] +
//             mat_A[560] * mat_B[539] +
//             mat_A[561] * mat_B[571] +
//             mat_A[562] * mat_B[603] +
//             mat_A[563] * mat_B[635] +
//             mat_A[564] * mat_B[667] +
//             mat_A[565] * mat_B[699] +
//             mat_A[566] * mat_B[731] +
//             mat_A[567] * mat_B[763] +
//             mat_A[568] * mat_B[795] +
//             mat_A[569] * mat_B[827] +
//             mat_A[570] * mat_B[859] +
//             mat_A[571] * mat_B[891] +
//             mat_A[572] * mat_B[923] +
//             mat_A[573] * mat_B[955] +
//             mat_A[574] * mat_B[987] +
//             mat_A[575] * mat_B[1019];
//  mat_C[572] <= 
//             mat_A[544] * mat_B[28] +
//             mat_A[545] * mat_B[60] +
//             mat_A[546] * mat_B[92] +
//             mat_A[547] * mat_B[124] +
//             mat_A[548] * mat_B[156] +
//             mat_A[549] * mat_B[188] +
//             mat_A[550] * mat_B[220] +
//             mat_A[551] * mat_B[252] +
//             mat_A[552] * mat_B[284] +
//             mat_A[553] * mat_B[316] +
//             mat_A[554] * mat_B[348] +
//             mat_A[555] * mat_B[380] +
//             mat_A[556] * mat_B[412] +
//             mat_A[557] * mat_B[444] +
//             mat_A[558] * mat_B[476] +
//             mat_A[559] * mat_B[508] +
//             mat_A[560] * mat_B[540] +
//             mat_A[561] * mat_B[572] +
//             mat_A[562] * mat_B[604] +
//             mat_A[563] * mat_B[636] +
//             mat_A[564] * mat_B[668] +
//             mat_A[565] * mat_B[700] +
//             mat_A[566] * mat_B[732] +
//             mat_A[567] * mat_B[764] +
//             mat_A[568] * mat_B[796] +
//             mat_A[569] * mat_B[828] +
//             mat_A[570] * mat_B[860] +
//             mat_A[571] * mat_B[892] +
//             mat_A[572] * mat_B[924] +
//             mat_A[573] * mat_B[956] +
//             mat_A[574] * mat_B[988] +
//             mat_A[575] * mat_B[1020];
//  mat_C[573] <= 
//             mat_A[544] * mat_B[29] +
//             mat_A[545] * mat_B[61] +
//             mat_A[546] * mat_B[93] +
//             mat_A[547] * mat_B[125] +
//             mat_A[548] * mat_B[157] +
//             mat_A[549] * mat_B[189] +
//             mat_A[550] * mat_B[221] +
//             mat_A[551] * mat_B[253] +
//             mat_A[552] * mat_B[285] +
//             mat_A[553] * mat_B[317] +
//             mat_A[554] * mat_B[349] +
//             mat_A[555] * mat_B[381] +
//             mat_A[556] * mat_B[413] +
//             mat_A[557] * mat_B[445] +
//             mat_A[558] * mat_B[477] +
//             mat_A[559] * mat_B[509] +
//             mat_A[560] * mat_B[541] +
//             mat_A[561] * mat_B[573] +
//             mat_A[562] * mat_B[605] +
//             mat_A[563] * mat_B[637] +
//             mat_A[564] * mat_B[669] +
//             mat_A[565] * mat_B[701] +
//             mat_A[566] * mat_B[733] +
//             mat_A[567] * mat_B[765] +
//             mat_A[568] * mat_B[797] +
//             mat_A[569] * mat_B[829] +
//             mat_A[570] * mat_B[861] +
//             mat_A[571] * mat_B[893] +
//             mat_A[572] * mat_B[925] +
//             mat_A[573] * mat_B[957] +
//             mat_A[574] * mat_B[989] +
//             mat_A[575] * mat_B[1021];
//  mat_C[574] <= 
//             mat_A[544] * mat_B[30] +
//             mat_A[545] * mat_B[62] +
//             mat_A[546] * mat_B[94] +
//             mat_A[547] * mat_B[126] +
//             mat_A[548] * mat_B[158] +
//             mat_A[549] * mat_B[190] +
//             mat_A[550] * mat_B[222] +
//             mat_A[551] * mat_B[254] +
//             mat_A[552] * mat_B[286] +
//             mat_A[553] * mat_B[318] +
//             mat_A[554] * mat_B[350] +
//             mat_A[555] * mat_B[382] +
//             mat_A[556] * mat_B[414] +
//             mat_A[557] * mat_B[446] +
//             mat_A[558] * mat_B[478] +
//             mat_A[559] * mat_B[510] +
//             mat_A[560] * mat_B[542] +
//             mat_A[561] * mat_B[574] +
//             mat_A[562] * mat_B[606] +
//             mat_A[563] * mat_B[638] +
//             mat_A[564] * mat_B[670] +
//             mat_A[565] * mat_B[702] +
//             mat_A[566] * mat_B[734] +
//             mat_A[567] * mat_B[766] +
//             mat_A[568] * mat_B[798] +
//             mat_A[569] * mat_B[830] +
//             mat_A[570] * mat_B[862] +
//             mat_A[571] * mat_B[894] +
//             mat_A[572] * mat_B[926] +
//             mat_A[573] * mat_B[958] +
//             mat_A[574] * mat_B[990] +
//             mat_A[575] * mat_B[1022];
//  mat_C[575] <= 
//             mat_A[544] * mat_B[31] +
//             mat_A[545] * mat_B[63] +
//             mat_A[546] * mat_B[95] +
//             mat_A[547] * mat_B[127] +
//             mat_A[548] * mat_B[159] +
//             mat_A[549] * mat_B[191] +
//             mat_A[550] * mat_B[223] +
//             mat_A[551] * mat_B[255] +
//             mat_A[552] * mat_B[287] +
//             mat_A[553] * mat_B[319] +
//             mat_A[554] * mat_B[351] +
//             mat_A[555] * mat_B[383] +
//             mat_A[556] * mat_B[415] +
//             mat_A[557] * mat_B[447] +
//             mat_A[558] * mat_B[479] +
//             mat_A[559] * mat_B[511] +
//             mat_A[560] * mat_B[543] +
//             mat_A[561] * mat_B[575] +
//             mat_A[562] * mat_B[607] +
//             mat_A[563] * mat_B[639] +
//             mat_A[564] * mat_B[671] +
//             mat_A[565] * mat_B[703] +
//             mat_A[566] * mat_B[735] +
//             mat_A[567] * mat_B[767] +
//             mat_A[568] * mat_B[799] +
//             mat_A[569] * mat_B[831] +
//             mat_A[570] * mat_B[863] +
//             mat_A[571] * mat_B[895] +
//             mat_A[572] * mat_B[927] +
//             mat_A[573] * mat_B[959] +
//             mat_A[574] * mat_B[991] +
//             mat_A[575] * mat_B[1023];
//  mat_C[576] <= 
//             mat_A[576] * mat_B[0] +
//             mat_A[577] * mat_B[32] +
//             mat_A[578] * mat_B[64] +
//             mat_A[579] * mat_B[96] +
//             mat_A[580] * mat_B[128] +
//             mat_A[581] * mat_B[160] +
//             mat_A[582] * mat_B[192] +
//             mat_A[583] * mat_B[224] +
//             mat_A[584] * mat_B[256] +
//             mat_A[585] * mat_B[288] +
//             mat_A[586] * mat_B[320] +
//             mat_A[587] * mat_B[352] +
//             mat_A[588] * mat_B[384] +
//             mat_A[589] * mat_B[416] +
//             mat_A[590] * mat_B[448] +
//             mat_A[591] * mat_B[480] +
//             mat_A[592] * mat_B[512] +
//             mat_A[593] * mat_B[544] +
//             mat_A[594] * mat_B[576] +
//             mat_A[595] * mat_B[608] +
//             mat_A[596] * mat_B[640] +
//             mat_A[597] * mat_B[672] +
//             mat_A[598] * mat_B[704] +
//             mat_A[599] * mat_B[736] +
//             mat_A[600] * mat_B[768] +
//             mat_A[601] * mat_B[800] +
//             mat_A[602] * mat_B[832] +
//             mat_A[603] * mat_B[864] +
//             mat_A[604] * mat_B[896] +
//             mat_A[605] * mat_B[928] +
//             mat_A[606] * mat_B[960] +
//             mat_A[607] * mat_B[992];
//  mat_C[577] <= 
//             mat_A[576] * mat_B[1] +
//             mat_A[577] * mat_B[33] +
//             mat_A[578] * mat_B[65] +
//             mat_A[579] * mat_B[97] +
//             mat_A[580] * mat_B[129] +
//             mat_A[581] * mat_B[161] +
//             mat_A[582] * mat_B[193] +
//             mat_A[583] * mat_B[225] +
//             mat_A[584] * mat_B[257] +
//             mat_A[585] * mat_B[289] +
//             mat_A[586] * mat_B[321] +
//             mat_A[587] * mat_B[353] +
//             mat_A[588] * mat_B[385] +
//             mat_A[589] * mat_B[417] +
//             mat_A[590] * mat_B[449] +
//             mat_A[591] * mat_B[481] +
//             mat_A[592] * mat_B[513] +
//             mat_A[593] * mat_B[545] +
//             mat_A[594] * mat_B[577] +
//             mat_A[595] * mat_B[609] +
//             mat_A[596] * mat_B[641] +
//             mat_A[597] * mat_B[673] +
//             mat_A[598] * mat_B[705] +
//             mat_A[599] * mat_B[737] +
//             mat_A[600] * mat_B[769] +
//             mat_A[601] * mat_B[801] +
//             mat_A[602] * mat_B[833] +
//             mat_A[603] * mat_B[865] +
//             mat_A[604] * mat_B[897] +
//             mat_A[605] * mat_B[929] +
//             mat_A[606] * mat_B[961] +
//             mat_A[607] * mat_B[993];
//  mat_C[578] <= 
//             mat_A[576] * mat_B[2] +
//             mat_A[577] * mat_B[34] +
//             mat_A[578] * mat_B[66] +
//             mat_A[579] * mat_B[98] +
//             mat_A[580] * mat_B[130] +
//             mat_A[581] * mat_B[162] +
//             mat_A[582] * mat_B[194] +
//             mat_A[583] * mat_B[226] +
//             mat_A[584] * mat_B[258] +
//             mat_A[585] * mat_B[290] +
//             mat_A[586] * mat_B[322] +
//             mat_A[587] * mat_B[354] +
//             mat_A[588] * mat_B[386] +
//             mat_A[589] * mat_B[418] +
//             mat_A[590] * mat_B[450] +
//             mat_A[591] * mat_B[482] +
//             mat_A[592] * mat_B[514] +
//             mat_A[593] * mat_B[546] +
//             mat_A[594] * mat_B[578] +
//             mat_A[595] * mat_B[610] +
//             mat_A[596] * mat_B[642] +
//             mat_A[597] * mat_B[674] +
//             mat_A[598] * mat_B[706] +
//             mat_A[599] * mat_B[738] +
//             mat_A[600] * mat_B[770] +
//             mat_A[601] * mat_B[802] +
//             mat_A[602] * mat_B[834] +
//             mat_A[603] * mat_B[866] +
//             mat_A[604] * mat_B[898] +
//             mat_A[605] * mat_B[930] +
//             mat_A[606] * mat_B[962] +
//             mat_A[607] * mat_B[994];
//  mat_C[579] <= 
//             mat_A[576] * mat_B[3] +
//             mat_A[577] * mat_B[35] +
//             mat_A[578] * mat_B[67] +
//             mat_A[579] * mat_B[99] +
//             mat_A[580] * mat_B[131] +
//             mat_A[581] * mat_B[163] +
//             mat_A[582] * mat_B[195] +
//             mat_A[583] * mat_B[227] +
//             mat_A[584] * mat_B[259] +
//             mat_A[585] * mat_B[291] +
//             mat_A[586] * mat_B[323] +
//             mat_A[587] * mat_B[355] +
//             mat_A[588] * mat_B[387] +
//             mat_A[589] * mat_B[419] +
//             mat_A[590] * mat_B[451] +
//             mat_A[591] * mat_B[483] +
//             mat_A[592] * mat_B[515] +
//             mat_A[593] * mat_B[547] +
//             mat_A[594] * mat_B[579] +
//             mat_A[595] * mat_B[611] +
//             mat_A[596] * mat_B[643] +
//             mat_A[597] * mat_B[675] +
//             mat_A[598] * mat_B[707] +
//             mat_A[599] * mat_B[739] +
//             mat_A[600] * mat_B[771] +
//             mat_A[601] * mat_B[803] +
//             mat_A[602] * mat_B[835] +
//             mat_A[603] * mat_B[867] +
//             mat_A[604] * mat_B[899] +
//             mat_A[605] * mat_B[931] +
//             mat_A[606] * mat_B[963] +
//             mat_A[607] * mat_B[995];
//  mat_C[580] <= 
//             mat_A[576] * mat_B[4] +
//             mat_A[577] * mat_B[36] +
//             mat_A[578] * mat_B[68] +
//             mat_A[579] * mat_B[100] +
//             mat_A[580] * mat_B[132] +
//             mat_A[581] * mat_B[164] +
//             mat_A[582] * mat_B[196] +
//             mat_A[583] * mat_B[228] +
//             mat_A[584] * mat_B[260] +
//             mat_A[585] * mat_B[292] +
//             mat_A[586] * mat_B[324] +
//             mat_A[587] * mat_B[356] +
//             mat_A[588] * mat_B[388] +
//             mat_A[589] * mat_B[420] +
//             mat_A[590] * mat_B[452] +
//             mat_A[591] * mat_B[484] +
//             mat_A[592] * mat_B[516] +
//             mat_A[593] * mat_B[548] +
//             mat_A[594] * mat_B[580] +
//             mat_A[595] * mat_B[612] +
//             mat_A[596] * mat_B[644] +
//             mat_A[597] * mat_B[676] +
//             mat_A[598] * mat_B[708] +
//             mat_A[599] * mat_B[740] +
//             mat_A[600] * mat_B[772] +
//             mat_A[601] * mat_B[804] +
//             mat_A[602] * mat_B[836] +
//             mat_A[603] * mat_B[868] +
//             mat_A[604] * mat_B[900] +
//             mat_A[605] * mat_B[932] +
//             mat_A[606] * mat_B[964] +
//             mat_A[607] * mat_B[996];
//  mat_C[581] <= 
//             mat_A[576] * mat_B[5] +
//             mat_A[577] * mat_B[37] +
//             mat_A[578] * mat_B[69] +
//             mat_A[579] * mat_B[101] +
//             mat_A[580] * mat_B[133] +
//             mat_A[581] * mat_B[165] +
//             mat_A[582] * mat_B[197] +
//             mat_A[583] * mat_B[229] +
//             mat_A[584] * mat_B[261] +
//             mat_A[585] * mat_B[293] +
//             mat_A[586] * mat_B[325] +
//             mat_A[587] * mat_B[357] +
//             mat_A[588] * mat_B[389] +
//             mat_A[589] * mat_B[421] +
//             mat_A[590] * mat_B[453] +
//             mat_A[591] * mat_B[485] +
//             mat_A[592] * mat_B[517] +
//             mat_A[593] * mat_B[549] +
//             mat_A[594] * mat_B[581] +
//             mat_A[595] * mat_B[613] +
//             mat_A[596] * mat_B[645] +
//             mat_A[597] * mat_B[677] +
//             mat_A[598] * mat_B[709] +
//             mat_A[599] * mat_B[741] +
//             mat_A[600] * mat_B[773] +
//             mat_A[601] * mat_B[805] +
//             mat_A[602] * mat_B[837] +
//             mat_A[603] * mat_B[869] +
//             mat_A[604] * mat_B[901] +
//             mat_A[605] * mat_B[933] +
//             mat_A[606] * mat_B[965] +
//             mat_A[607] * mat_B[997];
//  mat_C[582] <= 
//             mat_A[576] * mat_B[6] +
//             mat_A[577] * mat_B[38] +
//             mat_A[578] * mat_B[70] +
//             mat_A[579] * mat_B[102] +
//             mat_A[580] * mat_B[134] +
//             mat_A[581] * mat_B[166] +
//             mat_A[582] * mat_B[198] +
//             mat_A[583] * mat_B[230] +
//             mat_A[584] * mat_B[262] +
//             mat_A[585] * mat_B[294] +
//             mat_A[586] * mat_B[326] +
//             mat_A[587] * mat_B[358] +
//             mat_A[588] * mat_B[390] +
//             mat_A[589] * mat_B[422] +
//             mat_A[590] * mat_B[454] +
//             mat_A[591] * mat_B[486] +
//             mat_A[592] * mat_B[518] +
//             mat_A[593] * mat_B[550] +
//             mat_A[594] * mat_B[582] +
//             mat_A[595] * mat_B[614] +
//             mat_A[596] * mat_B[646] +
//             mat_A[597] * mat_B[678] +
//             mat_A[598] * mat_B[710] +
//             mat_A[599] * mat_B[742] +
//             mat_A[600] * mat_B[774] +
//             mat_A[601] * mat_B[806] +
//             mat_A[602] * mat_B[838] +
//             mat_A[603] * mat_B[870] +
//             mat_A[604] * mat_B[902] +
//             mat_A[605] * mat_B[934] +
//             mat_A[606] * mat_B[966] +
//             mat_A[607] * mat_B[998];
//  mat_C[583] <= 
//             mat_A[576] * mat_B[7] +
//             mat_A[577] * mat_B[39] +
//             mat_A[578] * mat_B[71] +
//             mat_A[579] * mat_B[103] +
//             mat_A[580] * mat_B[135] +
//             mat_A[581] * mat_B[167] +
//             mat_A[582] * mat_B[199] +
//             mat_A[583] * mat_B[231] +
//             mat_A[584] * mat_B[263] +
//             mat_A[585] * mat_B[295] +
//             mat_A[586] * mat_B[327] +
//             mat_A[587] * mat_B[359] +
//             mat_A[588] * mat_B[391] +
//             mat_A[589] * mat_B[423] +
//             mat_A[590] * mat_B[455] +
//             mat_A[591] * mat_B[487] +
//             mat_A[592] * mat_B[519] +
//             mat_A[593] * mat_B[551] +
//             mat_A[594] * mat_B[583] +
//             mat_A[595] * mat_B[615] +
//             mat_A[596] * mat_B[647] +
//             mat_A[597] * mat_B[679] +
//             mat_A[598] * mat_B[711] +
//             mat_A[599] * mat_B[743] +
//             mat_A[600] * mat_B[775] +
//             mat_A[601] * mat_B[807] +
//             mat_A[602] * mat_B[839] +
//             mat_A[603] * mat_B[871] +
//             mat_A[604] * mat_B[903] +
//             mat_A[605] * mat_B[935] +
//             mat_A[606] * mat_B[967] +
//             mat_A[607] * mat_B[999];
//  mat_C[584] <= 
//             mat_A[576] * mat_B[8] +
//             mat_A[577] * mat_B[40] +
//             mat_A[578] * mat_B[72] +
//             mat_A[579] * mat_B[104] +
//             mat_A[580] * mat_B[136] +
//             mat_A[581] * mat_B[168] +
//             mat_A[582] * mat_B[200] +
//             mat_A[583] * mat_B[232] +
//             mat_A[584] * mat_B[264] +
//             mat_A[585] * mat_B[296] +
//             mat_A[586] * mat_B[328] +
//             mat_A[587] * mat_B[360] +
//             mat_A[588] * mat_B[392] +
//             mat_A[589] * mat_B[424] +
//             mat_A[590] * mat_B[456] +
//             mat_A[591] * mat_B[488] +
//             mat_A[592] * mat_B[520] +
//             mat_A[593] * mat_B[552] +
//             mat_A[594] * mat_B[584] +
//             mat_A[595] * mat_B[616] +
//             mat_A[596] * mat_B[648] +
//             mat_A[597] * mat_B[680] +
//             mat_A[598] * mat_B[712] +
//             mat_A[599] * mat_B[744] +
//             mat_A[600] * mat_B[776] +
//             mat_A[601] * mat_B[808] +
//             mat_A[602] * mat_B[840] +
//             mat_A[603] * mat_B[872] +
//             mat_A[604] * mat_B[904] +
//             mat_A[605] * mat_B[936] +
//             mat_A[606] * mat_B[968] +
//             mat_A[607] * mat_B[1000];
//  mat_C[585] <= 
//             mat_A[576] * mat_B[9] +
//             mat_A[577] * mat_B[41] +
//             mat_A[578] * mat_B[73] +
//             mat_A[579] * mat_B[105] +
//             mat_A[580] * mat_B[137] +
//             mat_A[581] * mat_B[169] +
//             mat_A[582] * mat_B[201] +
//             mat_A[583] * mat_B[233] +
//             mat_A[584] * mat_B[265] +
//             mat_A[585] * mat_B[297] +
//             mat_A[586] * mat_B[329] +
//             mat_A[587] * mat_B[361] +
//             mat_A[588] * mat_B[393] +
//             mat_A[589] * mat_B[425] +
//             mat_A[590] * mat_B[457] +
//             mat_A[591] * mat_B[489] +
//             mat_A[592] * mat_B[521] +
//             mat_A[593] * mat_B[553] +
//             mat_A[594] * mat_B[585] +
//             mat_A[595] * mat_B[617] +
//             mat_A[596] * mat_B[649] +
//             mat_A[597] * mat_B[681] +
//             mat_A[598] * mat_B[713] +
//             mat_A[599] * mat_B[745] +
//             mat_A[600] * mat_B[777] +
//             mat_A[601] * mat_B[809] +
//             mat_A[602] * mat_B[841] +
//             mat_A[603] * mat_B[873] +
//             mat_A[604] * mat_B[905] +
//             mat_A[605] * mat_B[937] +
//             mat_A[606] * mat_B[969] +
//             mat_A[607] * mat_B[1001];
//  mat_C[586] <= 
//             mat_A[576] * mat_B[10] +
//             mat_A[577] * mat_B[42] +
//             mat_A[578] * mat_B[74] +
//             mat_A[579] * mat_B[106] +
//             mat_A[580] * mat_B[138] +
//             mat_A[581] * mat_B[170] +
//             mat_A[582] * mat_B[202] +
//             mat_A[583] * mat_B[234] +
//             mat_A[584] * mat_B[266] +
//             mat_A[585] * mat_B[298] +
//             mat_A[586] * mat_B[330] +
//             mat_A[587] * mat_B[362] +
//             mat_A[588] * mat_B[394] +
//             mat_A[589] * mat_B[426] +
//             mat_A[590] * mat_B[458] +
//             mat_A[591] * mat_B[490] +
//             mat_A[592] * mat_B[522] +
//             mat_A[593] * mat_B[554] +
//             mat_A[594] * mat_B[586] +
//             mat_A[595] * mat_B[618] +
//             mat_A[596] * mat_B[650] +
//             mat_A[597] * mat_B[682] +
//             mat_A[598] * mat_B[714] +
//             mat_A[599] * mat_B[746] +
//             mat_A[600] * mat_B[778] +
//             mat_A[601] * mat_B[810] +
//             mat_A[602] * mat_B[842] +
//             mat_A[603] * mat_B[874] +
//             mat_A[604] * mat_B[906] +
//             mat_A[605] * mat_B[938] +
//             mat_A[606] * mat_B[970] +
//             mat_A[607] * mat_B[1002];
//  mat_C[587] <= 
//             mat_A[576] * mat_B[11] +
//             mat_A[577] * mat_B[43] +
//             mat_A[578] * mat_B[75] +
//             mat_A[579] * mat_B[107] +
//             mat_A[580] * mat_B[139] +
//             mat_A[581] * mat_B[171] +
//             mat_A[582] * mat_B[203] +
//             mat_A[583] * mat_B[235] +
//             mat_A[584] * mat_B[267] +
//             mat_A[585] * mat_B[299] +
//             mat_A[586] * mat_B[331] +
//             mat_A[587] * mat_B[363] +
//             mat_A[588] * mat_B[395] +
//             mat_A[589] * mat_B[427] +
//             mat_A[590] * mat_B[459] +
//             mat_A[591] * mat_B[491] +
//             mat_A[592] * mat_B[523] +
//             mat_A[593] * mat_B[555] +
//             mat_A[594] * mat_B[587] +
//             mat_A[595] * mat_B[619] +
//             mat_A[596] * mat_B[651] +
//             mat_A[597] * mat_B[683] +
//             mat_A[598] * mat_B[715] +
//             mat_A[599] * mat_B[747] +
//             mat_A[600] * mat_B[779] +
//             mat_A[601] * mat_B[811] +
//             mat_A[602] * mat_B[843] +
//             mat_A[603] * mat_B[875] +
//             mat_A[604] * mat_B[907] +
//             mat_A[605] * mat_B[939] +
//             mat_A[606] * mat_B[971] +
//             mat_A[607] * mat_B[1003];
//  mat_C[588] <= 
//             mat_A[576] * mat_B[12] +
//             mat_A[577] * mat_B[44] +
//             mat_A[578] * mat_B[76] +
//             mat_A[579] * mat_B[108] +
//             mat_A[580] * mat_B[140] +
//             mat_A[581] * mat_B[172] +
//             mat_A[582] * mat_B[204] +
//             mat_A[583] * mat_B[236] +
//             mat_A[584] * mat_B[268] +
//             mat_A[585] * mat_B[300] +
//             mat_A[586] * mat_B[332] +
//             mat_A[587] * mat_B[364] +
//             mat_A[588] * mat_B[396] +
//             mat_A[589] * mat_B[428] +
//             mat_A[590] * mat_B[460] +
//             mat_A[591] * mat_B[492] +
//             mat_A[592] * mat_B[524] +
//             mat_A[593] * mat_B[556] +
//             mat_A[594] * mat_B[588] +
//             mat_A[595] * mat_B[620] +
//             mat_A[596] * mat_B[652] +
//             mat_A[597] * mat_B[684] +
//             mat_A[598] * mat_B[716] +
//             mat_A[599] * mat_B[748] +
//             mat_A[600] * mat_B[780] +
//             mat_A[601] * mat_B[812] +
//             mat_A[602] * mat_B[844] +
//             mat_A[603] * mat_B[876] +
//             mat_A[604] * mat_B[908] +
//             mat_A[605] * mat_B[940] +
//             mat_A[606] * mat_B[972] +
//             mat_A[607] * mat_B[1004];
//  mat_C[589] <= 
//             mat_A[576] * mat_B[13] +
//             mat_A[577] * mat_B[45] +
//             mat_A[578] * mat_B[77] +
//             mat_A[579] * mat_B[109] +
//             mat_A[580] * mat_B[141] +
//             mat_A[581] * mat_B[173] +
//             mat_A[582] * mat_B[205] +
//             mat_A[583] * mat_B[237] +
//             mat_A[584] * mat_B[269] +
//             mat_A[585] * mat_B[301] +
//             mat_A[586] * mat_B[333] +
//             mat_A[587] * mat_B[365] +
//             mat_A[588] * mat_B[397] +
//             mat_A[589] * mat_B[429] +
//             mat_A[590] * mat_B[461] +
//             mat_A[591] * mat_B[493] +
//             mat_A[592] * mat_B[525] +
//             mat_A[593] * mat_B[557] +
//             mat_A[594] * mat_B[589] +
//             mat_A[595] * mat_B[621] +
//             mat_A[596] * mat_B[653] +
//             mat_A[597] * mat_B[685] +
//             mat_A[598] * mat_B[717] +
//             mat_A[599] * mat_B[749] +
//             mat_A[600] * mat_B[781] +
//             mat_A[601] * mat_B[813] +
//             mat_A[602] * mat_B[845] +
//             mat_A[603] * mat_B[877] +
//             mat_A[604] * mat_B[909] +
//             mat_A[605] * mat_B[941] +
//             mat_A[606] * mat_B[973] +
//             mat_A[607] * mat_B[1005];
//  mat_C[590] <= 
//             mat_A[576] * mat_B[14] +
//             mat_A[577] * mat_B[46] +
//             mat_A[578] * mat_B[78] +
//             mat_A[579] * mat_B[110] +
//             mat_A[580] * mat_B[142] +
//             mat_A[581] * mat_B[174] +
//             mat_A[582] * mat_B[206] +
//             mat_A[583] * mat_B[238] +
//             mat_A[584] * mat_B[270] +
//             mat_A[585] * mat_B[302] +
//             mat_A[586] * mat_B[334] +
//             mat_A[587] * mat_B[366] +
//             mat_A[588] * mat_B[398] +
//             mat_A[589] * mat_B[430] +
//             mat_A[590] * mat_B[462] +
//             mat_A[591] * mat_B[494] +
//             mat_A[592] * mat_B[526] +
//             mat_A[593] * mat_B[558] +
//             mat_A[594] * mat_B[590] +
//             mat_A[595] * mat_B[622] +
//             mat_A[596] * mat_B[654] +
//             mat_A[597] * mat_B[686] +
//             mat_A[598] * mat_B[718] +
//             mat_A[599] * mat_B[750] +
//             mat_A[600] * mat_B[782] +
//             mat_A[601] * mat_B[814] +
//             mat_A[602] * mat_B[846] +
//             mat_A[603] * mat_B[878] +
//             mat_A[604] * mat_B[910] +
//             mat_A[605] * mat_B[942] +
//             mat_A[606] * mat_B[974] +
//             mat_A[607] * mat_B[1006];
//  mat_C[591] <= 
//             mat_A[576] * mat_B[15] +
//             mat_A[577] * mat_B[47] +
//             mat_A[578] * mat_B[79] +
//             mat_A[579] * mat_B[111] +
//             mat_A[580] * mat_B[143] +
//             mat_A[581] * mat_B[175] +
//             mat_A[582] * mat_B[207] +
//             mat_A[583] * mat_B[239] +
//             mat_A[584] * mat_B[271] +
//             mat_A[585] * mat_B[303] +
//             mat_A[586] * mat_B[335] +
//             mat_A[587] * mat_B[367] +
//             mat_A[588] * mat_B[399] +
//             mat_A[589] * mat_B[431] +
//             mat_A[590] * mat_B[463] +
//             mat_A[591] * mat_B[495] +
//             mat_A[592] * mat_B[527] +
//             mat_A[593] * mat_B[559] +
//             mat_A[594] * mat_B[591] +
//             mat_A[595] * mat_B[623] +
//             mat_A[596] * mat_B[655] +
//             mat_A[597] * mat_B[687] +
//             mat_A[598] * mat_B[719] +
//             mat_A[599] * mat_B[751] +
//             mat_A[600] * mat_B[783] +
//             mat_A[601] * mat_B[815] +
//             mat_A[602] * mat_B[847] +
//             mat_A[603] * mat_B[879] +
//             mat_A[604] * mat_B[911] +
//             mat_A[605] * mat_B[943] +
//             mat_A[606] * mat_B[975] +
//             mat_A[607] * mat_B[1007];
//  mat_C[592] <= 
//             mat_A[576] * mat_B[16] +
//             mat_A[577] * mat_B[48] +
//             mat_A[578] * mat_B[80] +
//             mat_A[579] * mat_B[112] +
//             mat_A[580] * mat_B[144] +
//             mat_A[581] * mat_B[176] +
//             mat_A[582] * mat_B[208] +
//             mat_A[583] * mat_B[240] +
//             mat_A[584] * mat_B[272] +
//             mat_A[585] * mat_B[304] +
//             mat_A[586] * mat_B[336] +
//             mat_A[587] * mat_B[368] +
//             mat_A[588] * mat_B[400] +
//             mat_A[589] * mat_B[432] +
//             mat_A[590] * mat_B[464] +
//             mat_A[591] * mat_B[496] +
//             mat_A[592] * mat_B[528] +
//             mat_A[593] * mat_B[560] +
//             mat_A[594] * mat_B[592] +
//             mat_A[595] * mat_B[624] +
//             mat_A[596] * mat_B[656] +
//             mat_A[597] * mat_B[688] +
//             mat_A[598] * mat_B[720] +
//             mat_A[599] * mat_B[752] +
//             mat_A[600] * mat_B[784] +
//             mat_A[601] * mat_B[816] +
//             mat_A[602] * mat_B[848] +
//             mat_A[603] * mat_B[880] +
//             mat_A[604] * mat_B[912] +
//             mat_A[605] * mat_B[944] +
//             mat_A[606] * mat_B[976] +
//             mat_A[607] * mat_B[1008];
//  mat_C[593] <= 
//             mat_A[576] * mat_B[17] +
//             mat_A[577] * mat_B[49] +
//             mat_A[578] * mat_B[81] +
//             mat_A[579] * mat_B[113] +
//             mat_A[580] * mat_B[145] +
//             mat_A[581] * mat_B[177] +
//             mat_A[582] * mat_B[209] +
//             mat_A[583] * mat_B[241] +
//             mat_A[584] * mat_B[273] +
//             mat_A[585] * mat_B[305] +
//             mat_A[586] * mat_B[337] +
//             mat_A[587] * mat_B[369] +
//             mat_A[588] * mat_B[401] +
//             mat_A[589] * mat_B[433] +
//             mat_A[590] * mat_B[465] +
//             mat_A[591] * mat_B[497] +
//             mat_A[592] * mat_B[529] +
//             mat_A[593] * mat_B[561] +
//             mat_A[594] * mat_B[593] +
//             mat_A[595] * mat_B[625] +
//             mat_A[596] * mat_B[657] +
//             mat_A[597] * mat_B[689] +
//             mat_A[598] * mat_B[721] +
//             mat_A[599] * mat_B[753] +
//             mat_A[600] * mat_B[785] +
//             mat_A[601] * mat_B[817] +
//             mat_A[602] * mat_B[849] +
//             mat_A[603] * mat_B[881] +
//             mat_A[604] * mat_B[913] +
//             mat_A[605] * mat_B[945] +
//             mat_A[606] * mat_B[977] +
//             mat_A[607] * mat_B[1009];
//  mat_C[594] <= 
//             mat_A[576] * mat_B[18] +
//             mat_A[577] * mat_B[50] +
//             mat_A[578] * mat_B[82] +
//             mat_A[579] * mat_B[114] +
//             mat_A[580] * mat_B[146] +
//             mat_A[581] * mat_B[178] +
//             mat_A[582] * mat_B[210] +
//             mat_A[583] * mat_B[242] +
//             mat_A[584] * mat_B[274] +
//             mat_A[585] * mat_B[306] +
//             mat_A[586] * mat_B[338] +
//             mat_A[587] * mat_B[370] +
//             mat_A[588] * mat_B[402] +
//             mat_A[589] * mat_B[434] +
//             mat_A[590] * mat_B[466] +
//             mat_A[591] * mat_B[498] +
//             mat_A[592] * mat_B[530] +
//             mat_A[593] * mat_B[562] +
//             mat_A[594] * mat_B[594] +
//             mat_A[595] * mat_B[626] +
//             mat_A[596] * mat_B[658] +
//             mat_A[597] * mat_B[690] +
//             mat_A[598] * mat_B[722] +
//             mat_A[599] * mat_B[754] +
//             mat_A[600] * mat_B[786] +
//             mat_A[601] * mat_B[818] +
//             mat_A[602] * mat_B[850] +
//             mat_A[603] * mat_B[882] +
//             mat_A[604] * mat_B[914] +
//             mat_A[605] * mat_B[946] +
//             mat_A[606] * mat_B[978] +
//             mat_A[607] * mat_B[1010];
//  mat_C[595] <= 
//             mat_A[576] * mat_B[19] +
//             mat_A[577] * mat_B[51] +
//             mat_A[578] * mat_B[83] +
//             mat_A[579] * mat_B[115] +
//             mat_A[580] * mat_B[147] +
//             mat_A[581] * mat_B[179] +
//             mat_A[582] * mat_B[211] +
//             mat_A[583] * mat_B[243] +
//             mat_A[584] * mat_B[275] +
//             mat_A[585] * mat_B[307] +
//             mat_A[586] * mat_B[339] +
//             mat_A[587] * mat_B[371] +
//             mat_A[588] * mat_B[403] +
//             mat_A[589] * mat_B[435] +
//             mat_A[590] * mat_B[467] +
//             mat_A[591] * mat_B[499] +
//             mat_A[592] * mat_B[531] +
//             mat_A[593] * mat_B[563] +
//             mat_A[594] * mat_B[595] +
//             mat_A[595] * mat_B[627] +
//             mat_A[596] * mat_B[659] +
//             mat_A[597] * mat_B[691] +
//             mat_A[598] * mat_B[723] +
//             mat_A[599] * mat_B[755] +
//             mat_A[600] * mat_B[787] +
//             mat_A[601] * mat_B[819] +
//             mat_A[602] * mat_B[851] +
//             mat_A[603] * mat_B[883] +
//             mat_A[604] * mat_B[915] +
//             mat_A[605] * mat_B[947] +
//             mat_A[606] * mat_B[979] +
//             mat_A[607] * mat_B[1011];
//  mat_C[596] <= 
//             mat_A[576] * mat_B[20] +
//             mat_A[577] * mat_B[52] +
//             mat_A[578] * mat_B[84] +
//             mat_A[579] * mat_B[116] +
//             mat_A[580] * mat_B[148] +
//             mat_A[581] * mat_B[180] +
//             mat_A[582] * mat_B[212] +
//             mat_A[583] * mat_B[244] +
//             mat_A[584] * mat_B[276] +
//             mat_A[585] * mat_B[308] +
//             mat_A[586] * mat_B[340] +
//             mat_A[587] * mat_B[372] +
//             mat_A[588] * mat_B[404] +
//             mat_A[589] * mat_B[436] +
//             mat_A[590] * mat_B[468] +
//             mat_A[591] * mat_B[500] +
//             mat_A[592] * mat_B[532] +
//             mat_A[593] * mat_B[564] +
//             mat_A[594] * mat_B[596] +
//             mat_A[595] * mat_B[628] +
//             mat_A[596] * mat_B[660] +
//             mat_A[597] * mat_B[692] +
//             mat_A[598] * mat_B[724] +
//             mat_A[599] * mat_B[756] +
//             mat_A[600] * mat_B[788] +
//             mat_A[601] * mat_B[820] +
//             mat_A[602] * mat_B[852] +
//             mat_A[603] * mat_B[884] +
//             mat_A[604] * mat_B[916] +
//             mat_A[605] * mat_B[948] +
//             mat_A[606] * mat_B[980] +
//             mat_A[607] * mat_B[1012];
//  mat_C[597] <= 
//             mat_A[576] * mat_B[21] +
//             mat_A[577] * mat_B[53] +
//             mat_A[578] * mat_B[85] +
//             mat_A[579] * mat_B[117] +
//             mat_A[580] * mat_B[149] +
//             mat_A[581] * mat_B[181] +
//             mat_A[582] * mat_B[213] +
//             mat_A[583] * mat_B[245] +
//             mat_A[584] * mat_B[277] +
//             mat_A[585] * mat_B[309] +
//             mat_A[586] * mat_B[341] +
//             mat_A[587] * mat_B[373] +
//             mat_A[588] * mat_B[405] +
//             mat_A[589] * mat_B[437] +
//             mat_A[590] * mat_B[469] +
//             mat_A[591] * mat_B[501] +
//             mat_A[592] * mat_B[533] +
//             mat_A[593] * mat_B[565] +
//             mat_A[594] * mat_B[597] +
//             mat_A[595] * mat_B[629] +
//             mat_A[596] * mat_B[661] +
//             mat_A[597] * mat_B[693] +
//             mat_A[598] * mat_B[725] +
//             mat_A[599] * mat_B[757] +
//             mat_A[600] * mat_B[789] +
//             mat_A[601] * mat_B[821] +
//             mat_A[602] * mat_B[853] +
//             mat_A[603] * mat_B[885] +
//             mat_A[604] * mat_B[917] +
//             mat_A[605] * mat_B[949] +
//             mat_A[606] * mat_B[981] +
//             mat_A[607] * mat_B[1013];
//  mat_C[598] <= 
//             mat_A[576] * mat_B[22] +
//             mat_A[577] * mat_B[54] +
//             mat_A[578] * mat_B[86] +
//             mat_A[579] * mat_B[118] +
//             mat_A[580] * mat_B[150] +
//             mat_A[581] * mat_B[182] +
//             mat_A[582] * mat_B[214] +
//             mat_A[583] * mat_B[246] +
//             mat_A[584] * mat_B[278] +
//             mat_A[585] * mat_B[310] +
//             mat_A[586] * mat_B[342] +
//             mat_A[587] * mat_B[374] +
//             mat_A[588] * mat_B[406] +
//             mat_A[589] * mat_B[438] +
//             mat_A[590] * mat_B[470] +
//             mat_A[591] * mat_B[502] +
//             mat_A[592] * mat_B[534] +
//             mat_A[593] * mat_B[566] +
//             mat_A[594] * mat_B[598] +
//             mat_A[595] * mat_B[630] +
//             mat_A[596] * mat_B[662] +
//             mat_A[597] * mat_B[694] +
//             mat_A[598] * mat_B[726] +
//             mat_A[599] * mat_B[758] +
//             mat_A[600] * mat_B[790] +
//             mat_A[601] * mat_B[822] +
//             mat_A[602] * mat_B[854] +
//             mat_A[603] * mat_B[886] +
//             mat_A[604] * mat_B[918] +
//             mat_A[605] * mat_B[950] +
//             mat_A[606] * mat_B[982] +
//             mat_A[607] * mat_B[1014];
//  mat_C[599] <= 
//             mat_A[576] * mat_B[23] +
//             mat_A[577] * mat_B[55] +
//             mat_A[578] * mat_B[87] +
//             mat_A[579] * mat_B[119] +
//             mat_A[580] * mat_B[151] +
//             mat_A[581] * mat_B[183] +
//             mat_A[582] * mat_B[215] +
//             mat_A[583] * mat_B[247] +
//             mat_A[584] * mat_B[279] +
//             mat_A[585] * mat_B[311] +
//             mat_A[586] * mat_B[343] +
//             mat_A[587] * mat_B[375] +
//             mat_A[588] * mat_B[407] +
//             mat_A[589] * mat_B[439] +
//             mat_A[590] * mat_B[471] +
//             mat_A[591] * mat_B[503] +
//             mat_A[592] * mat_B[535] +
//             mat_A[593] * mat_B[567] +
//             mat_A[594] * mat_B[599] +
//             mat_A[595] * mat_B[631] +
//             mat_A[596] * mat_B[663] +
//             mat_A[597] * mat_B[695] +
//             mat_A[598] * mat_B[727] +
//             mat_A[599] * mat_B[759] +
//             mat_A[600] * mat_B[791] +
//             mat_A[601] * mat_B[823] +
//             mat_A[602] * mat_B[855] +
//             mat_A[603] * mat_B[887] +
//             mat_A[604] * mat_B[919] +
//             mat_A[605] * mat_B[951] +
//             mat_A[606] * mat_B[983] +
//             mat_A[607] * mat_B[1015];
//  mat_C[600] <= 
//             mat_A[576] * mat_B[24] +
//             mat_A[577] * mat_B[56] +
//             mat_A[578] * mat_B[88] +
//             mat_A[579] * mat_B[120] +
//             mat_A[580] * mat_B[152] +
//             mat_A[581] * mat_B[184] +
//             mat_A[582] * mat_B[216] +
//             mat_A[583] * mat_B[248] +
//             mat_A[584] * mat_B[280] +
//             mat_A[585] * mat_B[312] +
//             mat_A[586] * mat_B[344] +
//             mat_A[587] * mat_B[376] +
//             mat_A[588] * mat_B[408] +
//             mat_A[589] * mat_B[440] +
//             mat_A[590] * mat_B[472] +
//             mat_A[591] * mat_B[504] +
//             mat_A[592] * mat_B[536] +
//             mat_A[593] * mat_B[568] +
//             mat_A[594] * mat_B[600] +
//             mat_A[595] * mat_B[632] +
//             mat_A[596] * mat_B[664] +
//             mat_A[597] * mat_B[696] +
//             mat_A[598] * mat_B[728] +
//             mat_A[599] * mat_B[760] +
//             mat_A[600] * mat_B[792] +
//             mat_A[601] * mat_B[824] +
//             mat_A[602] * mat_B[856] +
//             mat_A[603] * mat_B[888] +
//             mat_A[604] * mat_B[920] +
//             mat_A[605] * mat_B[952] +
//             mat_A[606] * mat_B[984] +
//             mat_A[607] * mat_B[1016];
//  mat_C[601] <= 
//             mat_A[576] * mat_B[25] +
//             mat_A[577] * mat_B[57] +
//             mat_A[578] * mat_B[89] +
//             mat_A[579] * mat_B[121] +
//             mat_A[580] * mat_B[153] +
//             mat_A[581] * mat_B[185] +
//             mat_A[582] * mat_B[217] +
//             mat_A[583] * mat_B[249] +
//             mat_A[584] * mat_B[281] +
//             mat_A[585] * mat_B[313] +
//             mat_A[586] * mat_B[345] +
//             mat_A[587] * mat_B[377] +
//             mat_A[588] * mat_B[409] +
//             mat_A[589] * mat_B[441] +
//             mat_A[590] * mat_B[473] +
//             mat_A[591] * mat_B[505] +
//             mat_A[592] * mat_B[537] +
//             mat_A[593] * mat_B[569] +
//             mat_A[594] * mat_B[601] +
//             mat_A[595] * mat_B[633] +
//             mat_A[596] * mat_B[665] +
//             mat_A[597] * mat_B[697] +
//             mat_A[598] * mat_B[729] +
//             mat_A[599] * mat_B[761] +
//             mat_A[600] * mat_B[793] +
//             mat_A[601] * mat_B[825] +
//             mat_A[602] * mat_B[857] +
//             mat_A[603] * mat_B[889] +
//             mat_A[604] * mat_B[921] +
//             mat_A[605] * mat_B[953] +
//             mat_A[606] * mat_B[985] +
//             mat_A[607] * mat_B[1017];
//  mat_C[602] <= 
//             mat_A[576] * mat_B[26] +
//             mat_A[577] * mat_B[58] +
//             mat_A[578] * mat_B[90] +
//             mat_A[579] * mat_B[122] +
//             mat_A[580] * mat_B[154] +
//             mat_A[581] * mat_B[186] +
//             mat_A[582] * mat_B[218] +
//             mat_A[583] * mat_B[250] +
//             mat_A[584] * mat_B[282] +
//             mat_A[585] * mat_B[314] +
//             mat_A[586] * mat_B[346] +
//             mat_A[587] * mat_B[378] +
//             mat_A[588] * mat_B[410] +
//             mat_A[589] * mat_B[442] +
//             mat_A[590] * mat_B[474] +
//             mat_A[591] * mat_B[506] +
//             mat_A[592] * mat_B[538] +
//             mat_A[593] * mat_B[570] +
//             mat_A[594] * mat_B[602] +
//             mat_A[595] * mat_B[634] +
//             mat_A[596] * mat_B[666] +
//             mat_A[597] * mat_B[698] +
//             mat_A[598] * mat_B[730] +
//             mat_A[599] * mat_B[762] +
//             mat_A[600] * mat_B[794] +
//             mat_A[601] * mat_B[826] +
//             mat_A[602] * mat_B[858] +
//             mat_A[603] * mat_B[890] +
//             mat_A[604] * mat_B[922] +
//             mat_A[605] * mat_B[954] +
//             mat_A[606] * mat_B[986] +
//             mat_A[607] * mat_B[1018];
//  mat_C[603] <= 
//             mat_A[576] * mat_B[27] +
//             mat_A[577] * mat_B[59] +
//             mat_A[578] * mat_B[91] +
//             mat_A[579] * mat_B[123] +
//             mat_A[580] * mat_B[155] +
//             mat_A[581] * mat_B[187] +
//             mat_A[582] * mat_B[219] +
//             mat_A[583] * mat_B[251] +
//             mat_A[584] * mat_B[283] +
//             mat_A[585] * mat_B[315] +
//             mat_A[586] * mat_B[347] +
//             mat_A[587] * mat_B[379] +
//             mat_A[588] * mat_B[411] +
//             mat_A[589] * mat_B[443] +
//             mat_A[590] * mat_B[475] +
//             mat_A[591] * mat_B[507] +
//             mat_A[592] * mat_B[539] +
//             mat_A[593] * mat_B[571] +
//             mat_A[594] * mat_B[603] +
//             mat_A[595] * mat_B[635] +
//             mat_A[596] * mat_B[667] +
//             mat_A[597] * mat_B[699] +
//             mat_A[598] * mat_B[731] +
//             mat_A[599] * mat_B[763] +
//             mat_A[600] * mat_B[795] +
//             mat_A[601] * mat_B[827] +
//             mat_A[602] * mat_B[859] +
//             mat_A[603] * mat_B[891] +
//             mat_A[604] * mat_B[923] +
//             mat_A[605] * mat_B[955] +
//             mat_A[606] * mat_B[987] +
//             mat_A[607] * mat_B[1019];
//  mat_C[604] <= 
//             mat_A[576] * mat_B[28] +
//             mat_A[577] * mat_B[60] +
//             mat_A[578] * mat_B[92] +
//             mat_A[579] * mat_B[124] +
//             mat_A[580] * mat_B[156] +
//             mat_A[581] * mat_B[188] +
//             mat_A[582] * mat_B[220] +
//             mat_A[583] * mat_B[252] +
//             mat_A[584] * mat_B[284] +
//             mat_A[585] * mat_B[316] +
//             mat_A[586] * mat_B[348] +
//             mat_A[587] * mat_B[380] +
//             mat_A[588] * mat_B[412] +
//             mat_A[589] * mat_B[444] +
//             mat_A[590] * mat_B[476] +
//             mat_A[591] * mat_B[508] +
//             mat_A[592] * mat_B[540] +
//             mat_A[593] * mat_B[572] +
//             mat_A[594] * mat_B[604] +
//             mat_A[595] * mat_B[636] +
//             mat_A[596] * mat_B[668] +
//             mat_A[597] * mat_B[700] +
//             mat_A[598] * mat_B[732] +
//             mat_A[599] * mat_B[764] +
//             mat_A[600] * mat_B[796] +
//             mat_A[601] * mat_B[828] +
//             mat_A[602] * mat_B[860] +
//             mat_A[603] * mat_B[892] +
//             mat_A[604] * mat_B[924] +
//             mat_A[605] * mat_B[956] +
//             mat_A[606] * mat_B[988] +
//             mat_A[607] * mat_B[1020];
//  mat_C[605] <= 
//             mat_A[576] * mat_B[29] +
//             mat_A[577] * mat_B[61] +
//             mat_A[578] * mat_B[93] +
//             mat_A[579] * mat_B[125] +
//             mat_A[580] * mat_B[157] +
//             mat_A[581] * mat_B[189] +
//             mat_A[582] * mat_B[221] +
//             mat_A[583] * mat_B[253] +
//             mat_A[584] * mat_B[285] +
//             mat_A[585] * mat_B[317] +
//             mat_A[586] * mat_B[349] +
//             mat_A[587] * mat_B[381] +
//             mat_A[588] * mat_B[413] +
//             mat_A[589] * mat_B[445] +
//             mat_A[590] * mat_B[477] +
//             mat_A[591] * mat_B[509] +
//             mat_A[592] * mat_B[541] +
//             mat_A[593] * mat_B[573] +
//             mat_A[594] * mat_B[605] +
//             mat_A[595] * mat_B[637] +
//             mat_A[596] * mat_B[669] +
//             mat_A[597] * mat_B[701] +
//             mat_A[598] * mat_B[733] +
//             mat_A[599] * mat_B[765] +
//             mat_A[600] * mat_B[797] +
//             mat_A[601] * mat_B[829] +
//             mat_A[602] * mat_B[861] +
//             mat_A[603] * mat_B[893] +
//             mat_A[604] * mat_B[925] +
//             mat_A[605] * mat_B[957] +
//             mat_A[606] * mat_B[989] +
//             mat_A[607] * mat_B[1021];
//  mat_C[606] <= 
//             mat_A[576] * mat_B[30] +
//             mat_A[577] * mat_B[62] +
//             mat_A[578] * mat_B[94] +
//             mat_A[579] * mat_B[126] +
//             mat_A[580] * mat_B[158] +
//             mat_A[581] * mat_B[190] +
//             mat_A[582] * mat_B[222] +
//             mat_A[583] * mat_B[254] +
//             mat_A[584] * mat_B[286] +
//             mat_A[585] * mat_B[318] +
//             mat_A[586] * mat_B[350] +
//             mat_A[587] * mat_B[382] +
//             mat_A[588] * mat_B[414] +
//             mat_A[589] * mat_B[446] +
//             mat_A[590] * mat_B[478] +
//             mat_A[591] * mat_B[510] +
//             mat_A[592] * mat_B[542] +
//             mat_A[593] * mat_B[574] +
//             mat_A[594] * mat_B[606] +
//             mat_A[595] * mat_B[638] +
//             mat_A[596] * mat_B[670] +
//             mat_A[597] * mat_B[702] +
//             mat_A[598] * mat_B[734] +
//             mat_A[599] * mat_B[766] +
//             mat_A[600] * mat_B[798] +
//             mat_A[601] * mat_B[830] +
//             mat_A[602] * mat_B[862] +
//             mat_A[603] * mat_B[894] +
//             mat_A[604] * mat_B[926] +
//             mat_A[605] * mat_B[958] +
//             mat_A[606] * mat_B[990] +
//             mat_A[607] * mat_B[1022];
//  mat_C[607] <= 
//             mat_A[576] * mat_B[31] +
//             mat_A[577] * mat_B[63] +
//             mat_A[578] * mat_B[95] +
//             mat_A[579] * mat_B[127] +
//             mat_A[580] * mat_B[159] +
//             mat_A[581] * mat_B[191] +
//             mat_A[582] * mat_B[223] +
//             mat_A[583] * mat_B[255] +
//             mat_A[584] * mat_B[287] +
//             mat_A[585] * mat_B[319] +
//             mat_A[586] * mat_B[351] +
//             mat_A[587] * mat_B[383] +
//             mat_A[588] * mat_B[415] +
//             mat_A[589] * mat_B[447] +
//             mat_A[590] * mat_B[479] +
//             mat_A[591] * mat_B[511] +
//             mat_A[592] * mat_B[543] +
//             mat_A[593] * mat_B[575] +
//             mat_A[594] * mat_B[607] +
//             mat_A[595] * mat_B[639] +
//             mat_A[596] * mat_B[671] +
//             mat_A[597] * mat_B[703] +
//             mat_A[598] * mat_B[735] +
//             mat_A[599] * mat_B[767] +
//             mat_A[600] * mat_B[799] +
//             mat_A[601] * mat_B[831] +
//             mat_A[602] * mat_B[863] +
//             mat_A[603] * mat_B[895] +
//             mat_A[604] * mat_B[927] +
//             mat_A[605] * mat_B[959] +
//             mat_A[606] * mat_B[991] +
//             mat_A[607] * mat_B[1023];
//  mat_C[608] <= 
//             mat_A[608] * mat_B[0] +
//             mat_A[609] * mat_B[32] +
//             mat_A[610] * mat_B[64] +
//             mat_A[611] * mat_B[96] +
//             mat_A[612] * mat_B[128] +
//             mat_A[613] * mat_B[160] +
//             mat_A[614] * mat_B[192] +
//             mat_A[615] * mat_B[224] +
//             mat_A[616] * mat_B[256] +
//             mat_A[617] * mat_B[288] +
//             mat_A[618] * mat_B[320] +
//             mat_A[619] * mat_B[352] +
//             mat_A[620] * mat_B[384] +
//             mat_A[621] * mat_B[416] +
//             mat_A[622] * mat_B[448] +
//             mat_A[623] * mat_B[480] +
//             mat_A[624] * mat_B[512] +
//             mat_A[625] * mat_B[544] +
//             mat_A[626] * mat_B[576] +
//             mat_A[627] * mat_B[608] +
//             mat_A[628] * mat_B[640] +
//             mat_A[629] * mat_B[672] +
//             mat_A[630] * mat_B[704] +
//             mat_A[631] * mat_B[736] +
//             mat_A[632] * mat_B[768] +
//             mat_A[633] * mat_B[800] +
//             mat_A[634] * mat_B[832] +
//             mat_A[635] * mat_B[864] +
//             mat_A[636] * mat_B[896] +
//             mat_A[637] * mat_B[928] +
//             mat_A[638] * mat_B[960] +
//             mat_A[639] * mat_B[992];
//  mat_C[609] <= 
//             mat_A[608] * mat_B[1] +
//             mat_A[609] * mat_B[33] +
//             mat_A[610] * mat_B[65] +
//             mat_A[611] * mat_B[97] +
//             mat_A[612] * mat_B[129] +
//             mat_A[613] * mat_B[161] +
//             mat_A[614] * mat_B[193] +
//             mat_A[615] * mat_B[225] +
//             mat_A[616] * mat_B[257] +
//             mat_A[617] * mat_B[289] +
//             mat_A[618] * mat_B[321] +
//             mat_A[619] * mat_B[353] +
//             mat_A[620] * mat_B[385] +
//             mat_A[621] * mat_B[417] +
//             mat_A[622] * mat_B[449] +
//             mat_A[623] * mat_B[481] +
//             mat_A[624] * mat_B[513] +
//             mat_A[625] * mat_B[545] +
//             mat_A[626] * mat_B[577] +
//             mat_A[627] * mat_B[609] +
//             mat_A[628] * mat_B[641] +
//             mat_A[629] * mat_B[673] +
//             mat_A[630] * mat_B[705] +
//             mat_A[631] * mat_B[737] +
//             mat_A[632] * mat_B[769] +
//             mat_A[633] * mat_B[801] +
//             mat_A[634] * mat_B[833] +
//             mat_A[635] * mat_B[865] +
//             mat_A[636] * mat_B[897] +
//             mat_A[637] * mat_B[929] +
//             mat_A[638] * mat_B[961] +
//             mat_A[639] * mat_B[993];
//  mat_C[610] <= 
//             mat_A[608] * mat_B[2] +
//             mat_A[609] * mat_B[34] +
//             mat_A[610] * mat_B[66] +
//             mat_A[611] * mat_B[98] +
//             mat_A[612] * mat_B[130] +
//             mat_A[613] * mat_B[162] +
//             mat_A[614] * mat_B[194] +
//             mat_A[615] * mat_B[226] +
//             mat_A[616] * mat_B[258] +
//             mat_A[617] * mat_B[290] +
//             mat_A[618] * mat_B[322] +
//             mat_A[619] * mat_B[354] +
//             mat_A[620] * mat_B[386] +
//             mat_A[621] * mat_B[418] +
//             mat_A[622] * mat_B[450] +
//             mat_A[623] * mat_B[482] +
//             mat_A[624] * mat_B[514] +
//             mat_A[625] * mat_B[546] +
//             mat_A[626] * mat_B[578] +
//             mat_A[627] * mat_B[610] +
//             mat_A[628] * mat_B[642] +
//             mat_A[629] * mat_B[674] +
//             mat_A[630] * mat_B[706] +
//             mat_A[631] * mat_B[738] +
//             mat_A[632] * mat_B[770] +
//             mat_A[633] * mat_B[802] +
//             mat_A[634] * mat_B[834] +
//             mat_A[635] * mat_B[866] +
//             mat_A[636] * mat_B[898] +
//             mat_A[637] * mat_B[930] +
//             mat_A[638] * mat_B[962] +
//             mat_A[639] * mat_B[994];
//  mat_C[611] <= 
//             mat_A[608] * mat_B[3] +
//             mat_A[609] * mat_B[35] +
//             mat_A[610] * mat_B[67] +
//             mat_A[611] * mat_B[99] +
//             mat_A[612] * mat_B[131] +
//             mat_A[613] * mat_B[163] +
//             mat_A[614] * mat_B[195] +
//             mat_A[615] * mat_B[227] +
//             mat_A[616] * mat_B[259] +
//             mat_A[617] * mat_B[291] +
//             mat_A[618] * mat_B[323] +
//             mat_A[619] * mat_B[355] +
//             mat_A[620] * mat_B[387] +
//             mat_A[621] * mat_B[419] +
//             mat_A[622] * mat_B[451] +
//             mat_A[623] * mat_B[483] +
//             mat_A[624] * mat_B[515] +
//             mat_A[625] * mat_B[547] +
//             mat_A[626] * mat_B[579] +
//             mat_A[627] * mat_B[611] +
//             mat_A[628] * mat_B[643] +
//             mat_A[629] * mat_B[675] +
//             mat_A[630] * mat_B[707] +
//             mat_A[631] * mat_B[739] +
//             mat_A[632] * mat_B[771] +
//             mat_A[633] * mat_B[803] +
//             mat_A[634] * mat_B[835] +
//             mat_A[635] * mat_B[867] +
//             mat_A[636] * mat_B[899] +
//             mat_A[637] * mat_B[931] +
//             mat_A[638] * mat_B[963] +
//             mat_A[639] * mat_B[995];
//  mat_C[612] <= 
//             mat_A[608] * mat_B[4] +
//             mat_A[609] * mat_B[36] +
//             mat_A[610] * mat_B[68] +
//             mat_A[611] * mat_B[100] +
//             mat_A[612] * mat_B[132] +
//             mat_A[613] * mat_B[164] +
//             mat_A[614] * mat_B[196] +
//             mat_A[615] * mat_B[228] +
//             mat_A[616] * mat_B[260] +
//             mat_A[617] * mat_B[292] +
//             mat_A[618] * mat_B[324] +
//             mat_A[619] * mat_B[356] +
//             mat_A[620] * mat_B[388] +
//             mat_A[621] * mat_B[420] +
//             mat_A[622] * mat_B[452] +
//             mat_A[623] * mat_B[484] +
//             mat_A[624] * mat_B[516] +
//             mat_A[625] * mat_B[548] +
//             mat_A[626] * mat_B[580] +
//             mat_A[627] * mat_B[612] +
//             mat_A[628] * mat_B[644] +
//             mat_A[629] * mat_B[676] +
//             mat_A[630] * mat_B[708] +
//             mat_A[631] * mat_B[740] +
//             mat_A[632] * mat_B[772] +
//             mat_A[633] * mat_B[804] +
//             mat_A[634] * mat_B[836] +
//             mat_A[635] * mat_B[868] +
//             mat_A[636] * mat_B[900] +
//             mat_A[637] * mat_B[932] +
//             mat_A[638] * mat_B[964] +
//             mat_A[639] * mat_B[996];
//  mat_C[613] <= 
//             mat_A[608] * mat_B[5] +
//             mat_A[609] * mat_B[37] +
//             mat_A[610] * mat_B[69] +
//             mat_A[611] * mat_B[101] +
//             mat_A[612] * mat_B[133] +
//             mat_A[613] * mat_B[165] +
//             mat_A[614] * mat_B[197] +
//             mat_A[615] * mat_B[229] +
//             mat_A[616] * mat_B[261] +
//             mat_A[617] * mat_B[293] +
//             mat_A[618] * mat_B[325] +
//             mat_A[619] * mat_B[357] +
//             mat_A[620] * mat_B[389] +
//             mat_A[621] * mat_B[421] +
//             mat_A[622] * mat_B[453] +
//             mat_A[623] * mat_B[485] +
//             mat_A[624] * mat_B[517] +
//             mat_A[625] * mat_B[549] +
//             mat_A[626] * mat_B[581] +
//             mat_A[627] * mat_B[613] +
//             mat_A[628] * mat_B[645] +
//             mat_A[629] * mat_B[677] +
//             mat_A[630] * mat_B[709] +
//             mat_A[631] * mat_B[741] +
//             mat_A[632] * mat_B[773] +
//             mat_A[633] * mat_B[805] +
//             mat_A[634] * mat_B[837] +
//             mat_A[635] * mat_B[869] +
//             mat_A[636] * mat_B[901] +
//             mat_A[637] * mat_B[933] +
//             mat_A[638] * mat_B[965] +
//             mat_A[639] * mat_B[997];
//  mat_C[614] <= 
//             mat_A[608] * mat_B[6] +
//             mat_A[609] * mat_B[38] +
//             mat_A[610] * mat_B[70] +
//             mat_A[611] * mat_B[102] +
//             mat_A[612] * mat_B[134] +
//             mat_A[613] * mat_B[166] +
//             mat_A[614] * mat_B[198] +
//             mat_A[615] * mat_B[230] +
//             mat_A[616] * mat_B[262] +
//             mat_A[617] * mat_B[294] +
//             mat_A[618] * mat_B[326] +
//             mat_A[619] * mat_B[358] +
//             mat_A[620] * mat_B[390] +
//             mat_A[621] * mat_B[422] +
//             mat_A[622] * mat_B[454] +
//             mat_A[623] * mat_B[486] +
//             mat_A[624] * mat_B[518] +
//             mat_A[625] * mat_B[550] +
//             mat_A[626] * mat_B[582] +
//             mat_A[627] * mat_B[614] +
//             mat_A[628] * mat_B[646] +
//             mat_A[629] * mat_B[678] +
//             mat_A[630] * mat_B[710] +
//             mat_A[631] * mat_B[742] +
//             mat_A[632] * mat_B[774] +
//             mat_A[633] * mat_B[806] +
//             mat_A[634] * mat_B[838] +
//             mat_A[635] * mat_B[870] +
//             mat_A[636] * mat_B[902] +
//             mat_A[637] * mat_B[934] +
//             mat_A[638] * mat_B[966] +
//             mat_A[639] * mat_B[998];
//  mat_C[615] <= 
//             mat_A[608] * mat_B[7] +
//             mat_A[609] * mat_B[39] +
//             mat_A[610] * mat_B[71] +
//             mat_A[611] * mat_B[103] +
//             mat_A[612] * mat_B[135] +
//             mat_A[613] * mat_B[167] +
//             mat_A[614] * mat_B[199] +
//             mat_A[615] * mat_B[231] +
//             mat_A[616] * mat_B[263] +
//             mat_A[617] * mat_B[295] +
//             mat_A[618] * mat_B[327] +
//             mat_A[619] * mat_B[359] +
//             mat_A[620] * mat_B[391] +
//             mat_A[621] * mat_B[423] +
//             mat_A[622] * mat_B[455] +
//             mat_A[623] * mat_B[487] +
//             mat_A[624] * mat_B[519] +
//             mat_A[625] * mat_B[551] +
//             mat_A[626] * mat_B[583] +
//             mat_A[627] * mat_B[615] +
//             mat_A[628] * mat_B[647] +
//             mat_A[629] * mat_B[679] +
//             mat_A[630] * mat_B[711] +
//             mat_A[631] * mat_B[743] +
//             mat_A[632] * mat_B[775] +
//             mat_A[633] * mat_B[807] +
//             mat_A[634] * mat_B[839] +
//             mat_A[635] * mat_B[871] +
//             mat_A[636] * mat_B[903] +
//             mat_A[637] * mat_B[935] +
//             mat_A[638] * mat_B[967] +
//             mat_A[639] * mat_B[999];
//  mat_C[616] <= 
//             mat_A[608] * mat_B[8] +
//             mat_A[609] * mat_B[40] +
//             mat_A[610] * mat_B[72] +
//             mat_A[611] * mat_B[104] +
//             mat_A[612] * mat_B[136] +
//             mat_A[613] * mat_B[168] +
//             mat_A[614] * mat_B[200] +
//             mat_A[615] * mat_B[232] +
//             mat_A[616] * mat_B[264] +
//             mat_A[617] * mat_B[296] +
//             mat_A[618] * mat_B[328] +
//             mat_A[619] * mat_B[360] +
//             mat_A[620] * mat_B[392] +
//             mat_A[621] * mat_B[424] +
//             mat_A[622] * mat_B[456] +
//             mat_A[623] * mat_B[488] +
//             mat_A[624] * mat_B[520] +
//             mat_A[625] * mat_B[552] +
//             mat_A[626] * mat_B[584] +
//             mat_A[627] * mat_B[616] +
//             mat_A[628] * mat_B[648] +
//             mat_A[629] * mat_B[680] +
//             mat_A[630] * mat_B[712] +
//             mat_A[631] * mat_B[744] +
//             mat_A[632] * mat_B[776] +
//             mat_A[633] * mat_B[808] +
//             mat_A[634] * mat_B[840] +
//             mat_A[635] * mat_B[872] +
//             mat_A[636] * mat_B[904] +
//             mat_A[637] * mat_B[936] +
//             mat_A[638] * mat_B[968] +
//             mat_A[639] * mat_B[1000];
//  mat_C[617] <= 
//             mat_A[608] * mat_B[9] +
//             mat_A[609] * mat_B[41] +
//             mat_A[610] * mat_B[73] +
//             mat_A[611] * mat_B[105] +
//             mat_A[612] * mat_B[137] +
//             mat_A[613] * mat_B[169] +
//             mat_A[614] * mat_B[201] +
//             mat_A[615] * mat_B[233] +
//             mat_A[616] * mat_B[265] +
//             mat_A[617] * mat_B[297] +
//             mat_A[618] * mat_B[329] +
//             mat_A[619] * mat_B[361] +
//             mat_A[620] * mat_B[393] +
//             mat_A[621] * mat_B[425] +
//             mat_A[622] * mat_B[457] +
//             mat_A[623] * mat_B[489] +
//             mat_A[624] * mat_B[521] +
//             mat_A[625] * mat_B[553] +
//             mat_A[626] * mat_B[585] +
//             mat_A[627] * mat_B[617] +
//             mat_A[628] * mat_B[649] +
//             mat_A[629] * mat_B[681] +
//             mat_A[630] * mat_B[713] +
//             mat_A[631] * mat_B[745] +
//             mat_A[632] * mat_B[777] +
//             mat_A[633] * mat_B[809] +
//             mat_A[634] * mat_B[841] +
//             mat_A[635] * mat_B[873] +
//             mat_A[636] * mat_B[905] +
//             mat_A[637] * mat_B[937] +
//             mat_A[638] * mat_B[969] +
//             mat_A[639] * mat_B[1001];
//  mat_C[618] <= 
//             mat_A[608] * mat_B[10] +
//             mat_A[609] * mat_B[42] +
//             mat_A[610] * mat_B[74] +
//             mat_A[611] * mat_B[106] +
//             mat_A[612] * mat_B[138] +
//             mat_A[613] * mat_B[170] +
//             mat_A[614] * mat_B[202] +
//             mat_A[615] * mat_B[234] +
//             mat_A[616] * mat_B[266] +
//             mat_A[617] * mat_B[298] +
//             mat_A[618] * mat_B[330] +
//             mat_A[619] * mat_B[362] +
//             mat_A[620] * mat_B[394] +
//             mat_A[621] * mat_B[426] +
//             mat_A[622] * mat_B[458] +
//             mat_A[623] * mat_B[490] +
//             mat_A[624] * mat_B[522] +
//             mat_A[625] * mat_B[554] +
//             mat_A[626] * mat_B[586] +
//             mat_A[627] * mat_B[618] +
//             mat_A[628] * mat_B[650] +
//             mat_A[629] * mat_B[682] +
//             mat_A[630] * mat_B[714] +
//             mat_A[631] * mat_B[746] +
//             mat_A[632] * mat_B[778] +
//             mat_A[633] * mat_B[810] +
//             mat_A[634] * mat_B[842] +
//             mat_A[635] * mat_B[874] +
//             mat_A[636] * mat_B[906] +
//             mat_A[637] * mat_B[938] +
//             mat_A[638] * mat_B[970] +
//             mat_A[639] * mat_B[1002];
//  mat_C[619] <= 
//             mat_A[608] * mat_B[11] +
//             mat_A[609] * mat_B[43] +
//             mat_A[610] * mat_B[75] +
//             mat_A[611] * mat_B[107] +
//             mat_A[612] * mat_B[139] +
//             mat_A[613] * mat_B[171] +
//             mat_A[614] * mat_B[203] +
//             mat_A[615] * mat_B[235] +
//             mat_A[616] * mat_B[267] +
//             mat_A[617] * mat_B[299] +
//             mat_A[618] * mat_B[331] +
//             mat_A[619] * mat_B[363] +
//             mat_A[620] * mat_B[395] +
//             mat_A[621] * mat_B[427] +
//             mat_A[622] * mat_B[459] +
//             mat_A[623] * mat_B[491] +
//             mat_A[624] * mat_B[523] +
//             mat_A[625] * mat_B[555] +
//             mat_A[626] * mat_B[587] +
//             mat_A[627] * mat_B[619] +
//             mat_A[628] * mat_B[651] +
//             mat_A[629] * mat_B[683] +
//             mat_A[630] * mat_B[715] +
//             mat_A[631] * mat_B[747] +
//             mat_A[632] * mat_B[779] +
//             mat_A[633] * mat_B[811] +
//             mat_A[634] * mat_B[843] +
//             mat_A[635] * mat_B[875] +
//             mat_A[636] * mat_B[907] +
//             mat_A[637] * mat_B[939] +
//             mat_A[638] * mat_B[971] +
//             mat_A[639] * mat_B[1003];
//  mat_C[620] <= 
//             mat_A[608] * mat_B[12] +
//             mat_A[609] * mat_B[44] +
//             mat_A[610] * mat_B[76] +
//             mat_A[611] * mat_B[108] +
//             mat_A[612] * mat_B[140] +
//             mat_A[613] * mat_B[172] +
//             mat_A[614] * mat_B[204] +
//             mat_A[615] * mat_B[236] +
//             mat_A[616] * mat_B[268] +
//             mat_A[617] * mat_B[300] +
//             mat_A[618] * mat_B[332] +
//             mat_A[619] * mat_B[364] +
//             mat_A[620] * mat_B[396] +
//             mat_A[621] * mat_B[428] +
//             mat_A[622] * mat_B[460] +
//             mat_A[623] * mat_B[492] +
//             mat_A[624] * mat_B[524] +
//             mat_A[625] * mat_B[556] +
//             mat_A[626] * mat_B[588] +
//             mat_A[627] * mat_B[620] +
//             mat_A[628] * mat_B[652] +
//             mat_A[629] * mat_B[684] +
//             mat_A[630] * mat_B[716] +
//             mat_A[631] * mat_B[748] +
//             mat_A[632] * mat_B[780] +
//             mat_A[633] * mat_B[812] +
//             mat_A[634] * mat_B[844] +
//             mat_A[635] * mat_B[876] +
//             mat_A[636] * mat_B[908] +
//             mat_A[637] * mat_B[940] +
//             mat_A[638] * mat_B[972] +
//             mat_A[639] * mat_B[1004];
//  mat_C[621] <= 
//             mat_A[608] * mat_B[13] +
//             mat_A[609] * mat_B[45] +
//             mat_A[610] * mat_B[77] +
//             mat_A[611] * mat_B[109] +
//             mat_A[612] * mat_B[141] +
//             mat_A[613] * mat_B[173] +
//             mat_A[614] * mat_B[205] +
//             mat_A[615] * mat_B[237] +
//             mat_A[616] * mat_B[269] +
//             mat_A[617] * mat_B[301] +
//             mat_A[618] * mat_B[333] +
//             mat_A[619] * mat_B[365] +
//             mat_A[620] * mat_B[397] +
//             mat_A[621] * mat_B[429] +
//             mat_A[622] * mat_B[461] +
//             mat_A[623] * mat_B[493] +
//             mat_A[624] * mat_B[525] +
//             mat_A[625] * mat_B[557] +
//             mat_A[626] * mat_B[589] +
//             mat_A[627] * mat_B[621] +
//             mat_A[628] * mat_B[653] +
//             mat_A[629] * mat_B[685] +
//             mat_A[630] * mat_B[717] +
//             mat_A[631] * mat_B[749] +
//             mat_A[632] * mat_B[781] +
//             mat_A[633] * mat_B[813] +
//             mat_A[634] * mat_B[845] +
//             mat_A[635] * mat_B[877] +
//             mat_A[636] * mat_B[909] +
//             mat_A[637] * mat_B[941] +
//             mat_A[638] * mat_B[973] +
//             mat_A[639] * mat_B[1005];
//  mat_C[622] <= 
//             mat_A[608] * mat_B[14] +
//             mat_A[609] * mat_B[46] +
//             mat_A[610] * mat_B[78] +
//             mat_A[611] * mat_B[110] +
//             mat_A[612] * mat_B[142] +
//             mat_A[613] * mat_B[174] +
//             mat_A[614] * mat_B[206] +
//             mat_A[615] * mat_B[238] +
//             mat_A[616] * mat_B[270] +
//             mat_A[617] * mat_B[302] +
//             mat_A[618] * mat_B[334] +
//             mat_A[619] * mat_B[366] +
//             mat_A[620] * mat_B[398] +
//             mat_A[621] * mat_B[430] +
//             mat_A[622] * mat_B[462] +
//             mat_A[623] * mat_B[494] +
//             mat_A[624] * mat_B[526] +
//             mat_A[625] * mat_B[558] +
//             mat_A[626] * mat_B[590] +
//             mat_A[627] * mat_B[622] +
//             mat_A[628] * mat_B[654] +
//             mat_A[629] * mat_B[686] +
//             mat_A[630] * mat_B[718] +
//             mat_A[631] * mat_B[750] +
//             mat_A[632] * mat_B[782] +
//             mat_A[633] * mat_B[814] +
//             mat_A[634] * mat_B[846] +
//             mat_A[635] * mat_B[878] +
//             mat_A[636] * mat_B[910] +
//             mat_A[637] * mat_B[942] +
//             mat_A[638] * mat_B[974] +
//             mat_A[639] * mat_B[1006];
//  mat_C[623] <= 
//             mat_A[608] * mat_B[15] +
//             mat_A[609] * mat_B[47] +
//             mat_A[610] * mat_B[79] +
//             mat_A[611] * mat_B[111] +
//             mat_A[612] * mat_B[143] +
//             mat_A[613] * mat_B[175] +
//             mat_A[614] * mat_B[207] +
//             mat_A[615] * mat_B[239] +
//             mat_A[616] * mat_B[271] +
//             mat_A[617] * mat_B[303] +
//             mat_A[618] * mat_B[335] +
//             mat_A[619] * mat_B[367] +
//             mat_A[620] * mat_B[399] +
//             mat_A[621] * mat_B[431] +
//             mat_A[622] * mat_B[463] +
//             mat_A[623] * mat_B[495] +
//             mat_A[624] * mat_B[527] +
//             mat_A[625] * mat_B[559] +
//             mat_A[626] * mat_B[591] +
//             mat_A[627] * mat_B[623] +
//             mat_A[628] * mat_B[655] +
//             mat_A[629] * mat_B[687] +
//             mat_A[630] * mat_B[719] +
//             mat_A[631] * mat_B[751] +
//             mat_A[632] * mat_B[783] +
//             mat_A[633] * mat_B[815] +
//             mat_A[634] * mat_B[847] +
//             mat_A[635] * mat_B[879] +
//             mat_A[636] * mat_B[911] +
//             mat_A[637] * mat_B[943] +
//             mat_A[638] * mat_B[975] +
//             mat_A[639] * mat_B[1007];
//  mat_C[624] <= 
//             mat_A[608] * mat_B[16] +
//             mat_A[609] * mat_B[48] +
//             mat_A[610] * mat_B[80] +
//             mat_A[611] * mat_B[112] +
//             mat_A[612] * mat_B[144] +
//             mat_A[613] * mat_B[176] +
//             mat_A[614] * mat_B[208] +
//             mat_A[615] * mat_B[240] +
//             mat_A[616] * mat_B[272] +
//             mat_A[617] * mat_B[304] +
//             mat_A[618] * mat_B[336] +
//             mat_A[619] * mat_B[368] +
//             mat_A[620] * mat_B[400] +
//             mat_A[621] * mat_B[432] +
//             mat_A[622] * mat_B[464] +
//             mat_A[623] * mat_B[496] +
//             mat_A[624] * mat_B[528] +
//             mat_A[625] * mat_B[560] +
//             mat_A[626] * mat_B[592] +
//             mat_A[627] * mat_B[624] +
//             mat_A[628] * mat_B[656] +
//             mat_A[629] * mat_B[688] +
//             mat_A[630] * mat_B[720] +
//             mat_A[631] * mat_B[752] +
//             mat_A[632] * mat_B[784] +
//             mat_A[633] * mat_B[816] +
//             mat_A[634] * mat_B[848] +
//             mat_A[635] * mat_B[880] +
//             mat_A[636] * mat_B[912] +
//             mat_A[637] * mat_B[944] +
//             mat_A[638] * mat_B[976] +
//             mat_A[639] * mat_B[1008];
//  mat_C[625] <= 
//             mat_A[608] * mat_B[17] +
//             mat_A[609] * mat_B[49] +
//             mat_A[610] * mat_B[81] +
//             mat_A[611] * mat_B[113] +
//             mat_A[612] * mat_B[145] +
//             mat_A[613] * mat_B[177] +
//             mat_A[614] * mat_B[209] +
//             mat_A[615] * mat_B[241] +
//             mat_A[616] * mat_B[273] +
//             mat_A[617] * mat_B[305] +
//             mat_A[618] * mat_B[337] +
//             mat_A[619] * mat_B[369] +
//             mat_A[620] * mat_B[401] +
//             mat_A[621] * mat_B[433] +
//             mat_A[622] * mat_B[465] +
//             mat_A[623] * mat_B[497] +
//             mat_A[624] * mat_B[529] +
//             mat_A[625] * mat_B[561] +
//             mat_A[626] * mat_B[593] +
//             mat_A[627] * mat_B[625] +
//             mat_A[628] * mat_B[657] +
//             mat_A[629] * mat_B[689] +
//             mat_A[630] * mat_B[721] +
//             mat_A[631] * mat_B[753] +
//             mat_A[632] * mat_B[785] +
//             mat_A[633] * mat_B[817] +
//             mat_A[634] * mat_B[849] +
//             mat_A[635] * mat_B[881] +
//             mat_A[636] * mat_B[913] +
//             mat_A[637] * mat_B[945] +
//             mat_A[638] * mat_B[977] +
//             mat_A[639] * mat_B[1009];
//  mat_C[626] <= 
//             mat_A[608] * mat_B[18] +
//             mat_A[609] * mat_B[50] +
//             mat_A[610] * mat_B[82] +
//             mat_A[611] * mat_B[114] +
//             mat_A[612] * mat_B[146] +
//             mat_A[613] * mat_B[178] +
//             mat_A[614] * mat_B[210] +
//             mat_A[615] * mat_B[242] +
//             mat_A[616] * mat_B[274] +
//             mat_A[617] * mat_B[306] +
//             mat_A[618] * mat_B[338] +
//             mat_A[619] * mat_B[370] +
//             mat_A[620] * mat_B[402] +
//             mat_A[621] * mat_B[434] +
//             mat_A[622] * mat_B[466] +
//             mat_A[623] * mat_B[498] +
//             mat_A[624] * mat_B[530] +
//             mat_A[625] * mat_B[562] +
//             mat_A[626] * mat_B[594] +
//             mat_A[627] * mat_B[626] +
//             mat_A[628] * mat_B[658] +
//             mat_A[629] * mat_B[690] +
//             mat_A[630] * mat_B[722] +
//             mat_A[631] * mat_B[754] +
//             mat_A[632] * mat_B[786] +
//             mat_A[633] * mat_B[818] +
//             mat_A[634] * mat_B[850] +
//             mat_A[635] * mat_B[882] +
//             mat_A[636] * mat_B[914] +
//             mat_A[637] * mat_B[946] +
//             mat_A[638] * mat_B[978] +
//             mat_A[639] * mat_B[1010];
//  mat_C[627] <= 
//             mat_A[608] * mat_B[19] +
//             mat_A[609] * mat_B[51] +
//             mat_A[610] * mat_B[83] +
//             mat_A[611] * mat_B[115] +
//             mat_A[612] * mat_B[147] +
//             mat_A[613] * mat_B[179] +
//             mat_A[614] * mat_B[211] +
//             mat_A[615] * mat_B[243] +
//             mat_A[616] * mat_B[275] +
//             mat_A[617] * mat_B[307] +
//             mat_A[618] * mat_B[339] +
//             mat_A[619] * mat_B[371] +
//             mat_A[620] * mat_B[403] +
//             mat_A[621] * mat_B[435] +
//             mat_A[622] * mat_B[467] +
//             mat_A[623] * mat_B[499] +
//             mat_A[624] * mat_B[531] +
//             mat_A[625] * mat_B[563] +
//             mat_A[626] * mat_B[595] +
//             mat_A[627] * mat_B[627] +
//             mat_A[628] * mat_B[659] +
//             mat_A[629] * mat_B[691] +
//             mat_A[630] * mat_B[723] +
//             mat_A[631] * mat_B[755] +
//             mat_A[632] * mat_B[787] +
//             mat_A[633] * mat_B[819] +
//             mat_A[634] * mat_B[851] +
//             mat_A[635] * mat_B[883] +
//             mat_A[636] * mat_B[915] +
//             mat_A[637] * mat_B[947] +
//             mat_A[638] * mat_B[979] +
//             mat_A[639] * mat_B[1011];
//  mat_C[628] <= 
//             mat_A[608] * mat_B[20] +
//             mat_A[609] * mat_B[52] +
//             mat_A[610] * mat_B[84] +
//             mat_A[611] * mat_B[116] +
//             mat_A[612] * mat_B[148] +
//             mat_A[613] * mat_B[180] +
//             mat_A[614] * mat_B[212] +
//             mat_A[615] * mat_B[244] +
//             mat_A[616] * mat_B[276] +
//             mat_A[617] * mat_B[308] +
//             mat_A[618] * mat_B[340] +
//             mat_A[619] * mat_B[372] +
//             mat_A[620] * mat_B[404] +
//             mat_A[621] * mat_B[436] +
//             mat_A[622] * mat_B[468] +
//             mat_A[623] * mat_B[500] +
//             mat_A[624] * mat_B[532] +
//             mat_A[625] * mat_B[564] +
//             mat_A[626] * mat_B[596] +
//             mat_A[627] * mat_B[628] +
//             mat_A[628] * mat_B[660] +
//             mat_A[629] * mat_B[692] +
//             mat_A[630] * mat_B[724] +
//             mat_A[631] * mat_B[756] +
//             mat_A[632] * mat_B[788] +
//             mat_A[633] * mat_B[820] +
//             mat_A[634] * mat_B[852] +
//             mat_A[635] * mat_B[884] +
//             mat_A[636] * mat_B[916] +
//             mat_A[637] * mat_B[948] +
//             mat_A[638] * mat_B[980] +
//             mat_A[639] * mat_B[1012];
//  mat_C[629] <= 
//             mat_A[608] * mat_B[21] +
//             mat_A[609] * mat_B[53] +
//             mat_A[610] * mat_B[85] +
//             mat_A[611] * mat_B[117] +
//             mat_A[612] * mat_B[149] +
//             mat_A[613] * mat_B[181] +
//             mat_A[614] * mat_B[213] +
//             mat_A[615] * mat_B[245] +
//             mat_A[616] * mat_B[277] +
//             mat_A[617] * mat_B[309] +
//             mat_A[618] * mat_B[341] +
//             mat_A[619] * mat_B[373] +
//             mat_A[620] * mat_B[405] +
//             mat_A[621] * mat_B[437] +
//             mat_A[622] * mat_B[469] +
//             mat_A[623] * mat_B[501] +
//             mat_A[624] * mat_B[533] +
//             mat_A[625] * mat_B[565] +
//             mat_A[626] * mat_B[597] +
//             mat_A[627] * mat_B[629] +
//             mat_A[628] * mat_B[661] +
//             mat_A[629] * mat_B[693] +
//             mat_A[630] * mat_B[725] +
//             mat_A[631] * mat_B[757] +
//             mat_A[632] * mat_B[789] +
//             mat_A[633] * mat_B[821] +
//             mat_A[634] * mat_B[853] +
//             mat_A[635] * mat_B[885] +
//             mat_A[636] * mat_B[917] +
//             mat_A[637] * mat_B[949] +
//             mat_A[638] * mat_B[981] +
//             mat_A[639] * mat_B[1013];
//  mat_C[630] <= 
//             mat_A[608] * mat_B[22] +
//             mat_A[609] * mat_B[54] +
//             mat_A[610] * mat_B[86] +
//             mat_A[611] * mat_B[118] +
//             mat_A[612] * mat_B[150] +
//             mat_A[613] * mat_B[182] +
//             mat_A[614] * mat_B[214] +
//             mat_A[615] * mat_B[246] +
//             mat_A[616] * mat_B[278] +
//             mat_A[617] * mat_B[310] +
//             mat_A[618] * mat_B[342] +
//             mat_A[619] * mat_B[374] +
//             mat_A[620] * mat_B[406] +
//             mat_A[621] * mat_B[438] +
//             mat_A[622] * mat_B[470] +
//             mat_A[623] * mat_B[502] +
//             mat_A[624] * mat_B[534] +
//             mat_A[625] * mat_B[566] +
//             mat_A[626] * mat_B[598] +
//             mat_A[627] * mat_B[630] +
//             mat_A[628] * mat_B[662] +
//             mat_A[629] * mat_B[694] +
//             mat_A[630] * mat_B[726] +
//             mat_A[631] * mat_B[758] +
//             mat_A[632] * mat_B[790] +
//             mat_A[633] * mat_B[822] +
//             mat_A[634] * mat_B[854] +
//             mat_A[635] * mat_B[886] +
//             mat_A[636] * mat_B[918] +
//             mat_A[637] * mat_B[950] +
//             mat_A[638] * mat_B[982] +
//             mat_A[639] * mat_B[1014];
//  mat_C[631] <= 
//             mat_A[608] * mat_B[23] +
//             mat_A[609] * mat_B[55] +
//             mat_A[610] * mat_B[87] +
//             mat_A[611] * mat_B[119] +
//             mat_A[612] * mat_B[151] +
//             mat_A[613] * mat_B[183] +
//             mat_A[614] * mat_B[215] +
//             mat_A[615] * mat_B[247] +
//             mat_A[616] * mat_B[279] +
//             mat_A[617] * mat_B[311] +
//             mat_A[618] * mat_B[343] +
//             mat_A[619] * mat_B[375] +
//             mat_A[620] * mat_B[407] +
//             mat_A[621] * mat_B[439] +
//             mat_A[622] * mat_B[471] +
//             mat_A[623] * mat_B[503] +
//             mat_A[624] * mat_B[535] +
//             mat_A[625] * mat_B[567] +
//             mat_A[626] * mat_B[599] +
//             mat_A[627] * mat_B[631] +
//             mat_A[628] * mat_B[663] +
//             mat_A[629] * mat_B[695] +
//             mat_A[630] * mat_B[727] +
//             mat_A[631] * mat_B[759] +
//             mat_A[632] * mat_B[791] +
//             mat_A[633] * mat_B[823] +
//             mat_A[634] * mat_B[855] +
//             mat_A[635] * mat_B[887] +
//             mat_A[636] * mat_B[919] +
//             mat_A[637] * mat_B[951] +
//             mat_A[638] * mat_B[983] +
//             mat_A[639] * mat_B[1015];
//  mat_C[632] <= 
//             mat_A[608] * mat_B[24] +
//             mat_A[609] * mat_B[56] +
//             mat_A[610] * mat_B[88] +
//             mat_A[611] * mat_B[120] +
//             mat_A[612] * mat_B[152] +
//             mat_A[613] * mat_B[184] +
//             mat_A[614] * mat_B[216] +
//             mat_A[615] * mat_B[248] +
//             mat_A[616] * mat_B[280] +
//             mat_A[617] * mat_B[312] +
//             mat_A[618] * mat_B[344] +
//             mat_A[619] * mat_B[376] +
//             mat_A[620] * mat_B[408] +
//             mat_A[621] * mat_B[440] +
//             mat_A[622] * mat_B[472] +
//             mat_A[623] * mat_B[504] +
//             mat_A[624] * mat_B[536] +
//             mat_A[625] * mat_B[568] +
//             mat_A[626] * mat_B[600] +
//             mat_A[627] * mat_B[632] +
//             mat_A[628] * mat_B[664] +
//             mat_A[629] * mat_B[696] +
//             mat_A[630] * mat_B[728] +
//             mat_A[631] * mat_B[760] +
//             mat_A[632] * mat_B[792] +
//             mat_A[633] * mat_B[824] +
//             mat_A[634] * mat_B[856] +
//             mat_A[635] * mat_B[888] +
//             mat_A[636] * mat_B[920] +
//             mat_A[637] * mat_B[952] +
//             mat_A[638] * mat_B[984] +
//             mat_A[639] * mat_B[1016];
//  mat_C[633] <= 
//             mat_A[608] * mat_B[25] +
//             mat_A[609] * mat_B[57] +
//             mat_A[610] * mat_B[89] +
//             mat_A[611] * mat_B[121] +
//             mat_A[612] * mat_B[153] +
//             mat_A[613] * mat_B[185] +
//             mat_A[614] * mat_B[217] +
//             mat_A[615] * mat_B[249] +
//             mat_A[616] * mat_B[281] +
//             mat_A[617] * mat_B[313] +
//             mat_A[618] * mat_B[345] +
//             mat_A[619] * mat_B[377] +
//             mat_A[620] * mat_B[409] +
//             mat_A[621] * mat_B[441] +
//             mat_A[622] * mat_B[473] +
//             mat_A[623] * mat_B[505] +
//             mat_A[624] * mat_B[537] +
//             mat_A[625] * mat_B[569] +
//             mat_A[626] * mat_B[601] +
//             mat_A[627] * mat_B[633] +
//             mat_A[628] * mat_B[665] +
//             mat_A[629] * mat_B[697] +
//             mat_A[630] * mat_B[729] +
//             mat_A[631] * mat_B[761] +
//             mat_A[632] * mat_B[793] +
//             mat_A[633] * mat_B[825] +
//             mat_A[634] * mat_B[857] +
//             mat_A[635] * mat_B[889] +
//             mat_A[636] * mat_B[921] +
//             mat_A[637] * mat_B[953] +
//             mat_A[638] * mat_B[985] +
//             mat_A[639] * mat_B[1017];
//  mat_C[634] <= 
//             mat_A[608] * mat_B[26] +
//             mat_A[609] * mat_B[58] +
//             mat_A[610] * mat_B[90] +
//             mat_A[611] * mat_B[122] +
//             mat_A[612] * mat_B[154] +
//             mat_A[613] * mat_B[186] +
//             mat_A[614] * mat_B[218] +
//             mat_A[615] * mat_B[250] +
//             mat_A[616] * mat_B[282] +
//             mat_A[617] * mat_B[314] +
//             mat_A[618] * mat_B[346] +
//             mat_A[619] * mat_B[378] +
//             mat_A[620] * mat_B[410] +
//             mat_A[621] * mat_B[442] +
//             mat_A[622] * mat_B[474] +
//             mat_A[623] * mat_B[506] +
//             mat_A[624] * mat_B[538] +
//             mat_A[625] * mat_B[570] +
//             mat_A[626] * mat_B[602] +
//             mat_A[627] * mat_B[634] +
//             mat_A[628] * mat_B[666] +
//             mat_A[629] * mat_B[698] +
//             mat_A[630] * mat_B[730] +
//             mat_A[631] * mat_B[762] +
//             mat_A[632] * mat_B[794] +
//             mat_A[633] * mat_B[826] +
//             mat_A[634] * mat_B[858] +
//             mat_A[635] * mat_B[890] +
//             mat_A[636] * mat_B[922] +
//             mat_A[637] * mat_B[954] +
//             mat_A[638] * mat_B[986] +
//             mat_A[639] * mat_B[1018];
//  mat_C[635] <= 
//             mat_A[608] * mat_B[27] +
//             mat_A[609] * mat_B[59] +
//             mat_A[610] * mat_B[91] +
//             mat_A[611] * mat_B[123] +
//             mat_A[612] * mat_B[155] +
//             mat_A[613] * mat_B[187] +
//             mat_A[614] * mat_B[219] +
//             mat_A[615] * mat_B[251] +
//             mat_A[616] * mat_B[283] +
//             mat_A[617] * mat_B[315] +
//             mat_A[618] * mat_B[347] +
//             mat_A[619] * mat_B[379] +
//             mat_A[620] * mat_B[411] +
//             mat_A[621] * mat_B[443] +
//             mat_A[622] * mat_B[475] +
//             mat_A[623] * mat_B[507] +
//             mat_A[624] * mat_B[539] +
//             mat_A[625] * mat_B[571] +
//             mat_A[626] * mat_B[603] +
//             mat_A[627] * mat_B[635] +
//             mat_A[628] * mat_B[667] +
//             mat_A[629] * mat_B[699] +
//             mat_A[630] * mat_B[731] +
//             mat_A[631] * mat_B[763] +
//             mat_A[632] * mat_B[795] +
//             mat_A[633] * mat_B[827] +
//             mat_A[634] * mat_B[859] +
//             mat_A[635] * mat_B[891] +
//             mat_A[636] * mat_B[923] +
//             mat_A[637] * mat_B[955] +
//             mat_A[638] * mat_B[987] +
//             mat_A[639] * mat_B[1019];
//  mat_C[636] <= 
//             mat_A[608] * mat_B[28] +
//             mat_A[609] * mat_B[60] +
//             mat_A[610] * mat_B[92] +
//             mat_A[611] * mat_B[124] +
//             mat_A[612] * mat_B[156] +
//             mat_A[613] * mat_B[188] +
//             mat_A[614] * mat_B[220] +
//             mat_A[615] * mat_B[252] +
//             mat_A[616] * mat_B[284] +
//             mat_A[617] * mat_B[316] +
//             mat_A[618] * mat_B[348] +
//             mat_A[619] * mat_B[380] +
//             mat_A[620] * mat_B[412] +
//             mat_A[621] * mat_B[444] +
//             mat_A[622] * mat_B[476] +
//             mat_A[623] * mat_B[508] +
//             mat_A[624] * mat_B[540] +
//             mat_A[625] * mat_B[572] +
//             mat_A[626] * mat_B[604] +
//             mat_A[627] * mat_B[636] +
//             mat_A[628] * mat_B[668] +
//             mat_A[629] * mat_B[700] +
//             mat_A[630] * mat_B[732] +
//             mat_A[631] * mat_B[764] +
//             mat_A[632] * mat_B[796] +
//             mat_A[633] * mat_B[828] +
//             mat_A[634] * mat_B[860] +
//             mat_A[635] * mat_B[892] +
//             mat_A[636] * mat_B[924] +
//             mat_A[637] * mat_B[956] +
//             mat_A[638] * mat_B[988] +
//             mat_A[639] * mat_B[1020];
//  mat_C[637] <= 
//             mat_A[608] * mat_B[29] +
//             mat_A[609] * mat_B[61] +
//             mat_A[610] * mat_B[93] +
//             mat_A[611] * mat_B[125] +
//             mat_A[612] * mat_B[157] +
//             mat_A[613] * mat_B[189] +
//             mat_A[614] * mat_B[221] +
//             mat_A[615] * mat_B[253] +
//             mat_A[616] * mat_B[285] +
//             mat_A[617] * mat_B[317] +
//             mat_A[618] * mat_B[349] +
//             mat_A[619] * mat_B[381] +
//             mat_A[620] * mat_B[413] +
//             mat_A[621] * mat_B[445] +
//             mat_A[622] * mat_B[477] +
//             mat_A[623] * mat_B[509] +
//             mat_A[624] * mat_B[541] +
//             mat_A[625] * mat_B[573] +
//             mat_A[626] * mat_B[605] +
//             mat_A[627] * mat_B[637] +
//             mat_A[628] * mat_B[669] +
//             mat_A[629] * mat_B[701] +
//             mat_A[630] * mat_B[733] +
//             mat_A[631] * mat_B[765] +
//             mat_A[632] * mat_B[797] +
//             mat_A[633] * mat_B[829] +
//             mat_A[634] * mat_B[861] +
//             mat_A[635] * mat_B[893] +
//             mat_A[636] * mat_B[925] +
//             mat_A[637] * mat_B[957] +
//             mat_A[638] * mat_B[989] +
//             mat_A[639] * mat_B[1021];
//  mat_C[638] <= 
//             mat_A[608] * mat_B[30] +
//             mat_A[609] * mat_B[62] +
//             mat_A[610] * mat_B[94] +
//             mat_A[611] * mat_B[126] +
//             mat_A[612] * mat_B[158] +
//             mat_A[613] * mat_B[190] +
//             mat_A[614] * mat_B[222] +
//             mat_A[615] * mat_B[254] +
//             mat_A[616] * mat_B[286] +
//             mat_A[617] * mat_B[318] +
//             mat_A[618] * mat_B[350] +
//             mat_A[619] * mat_B[382] +
//             mat_A[620] * mat_B[414] +
//             mat_A[621] * mat_B[446] +
//             mat_A[622] * mat_B[478] +
//             mat_A[623] * mat_B[510] +
//             mat_A[624] * mat_B[542] +
//             mat_A[625] * mat_B[574] +
//             mat_A[626] * mat_B[606] +
//             mat_A[627] * mat_B[638] +
//             mat_A[628] * mat_B[670] +
//             mat_A[629] * mat_B[702] +
//             mat_A[630] * mat_B[734] +
//             mat_A[631] * mat_B[766] +
//             mat_A[632] * mat_B[798] +
//             mat_A[633] * mat_B[830] +
//             mat_A[634] * mat_B[862] +
//             mat_A[635] * mat_B[894] +
//             mat_A[636] * mat_B[926] +
//             mat_A[637] * mat_B[958] +
//             mat_A[638] * mat_B[990] +
//             mat_A[639] * mat_B[1022];
//  mat_C[639] <= 
//             mat_A[608] * mat_B[31] +
//             mat_A[609] * mat_B[63] +
//             mat_A[610] * mat_B[95] +
//             mat_A[611] * mat_B[127] +
//             mat_A[612] * mat_B[159] +
//             mat_A[613] * mat_B[191] +
//             mat_A[614] * mat_B[223] +
//             mat_A[615] * mat_B[255] +
//             mat_A[616] * mat_B[287] +
//             mat_A[617] * mat_B[319] +
//             mat_A[618] * mat_B[351] +
//             mat_A[619] * mat_B[383] +
//             mat_A[620] * mat_B[415] +
//             mat_A[621] * mat_B[447] +
//             mat_A[622] * mat_B[479] +
//             mat_A[623] * mat_B[511] +
//             mat_A[624] * mat_B[543] +
//             mat_A[625] * mat_B[575] +
//             mat_A[626] * mat_B[607] +
//             mat_A[627] * mat_B[639] +
//             mat_A[628] * mat_B[671] +
//             mat_A[629] * mat_B[703] +
//             mat_A[630] * mat_B[735] +
//             mat_A[631] * mat_B[767] +
//             mat_A[632] * mat_B[799] +
//             mat_A[633] * mat_B[831] +
//             mat_A[634] * mat_B[863] +
//             mat_A[635] * mat_B[895] +
//             mat_A[636] * mat_B[927] +
//             mat_A[637] * mat_B[959] +
//             mat_A[638] * mat_B[991] +
//             mat_A[639] * mat_B[1023];
//  mat_C[640] <= 
//             mat_A[640] * mat_B[0] +
//             mat_A[641] * mat_B[32] +
//             mat_A[642] * mat_B[64] +
//             mat_A[643] * mat_B[96] +
//             mat_A[644] * mat_B[128] +
//             mat_A[645] * mat_B[160] +
//             mat_A[646] * mat_B[192] +
//             mat_A[647] * mat_B[224] +
//             mat_A[648] * mat_B[256] +
//             mat_A[649] * mat_B[288] +
//             mat_A[650] * mat_B[320] +
//             mat_A[651] * mat_B[352] +
//             mat_A[652] * mat_B[384] +
//             mat_A[653] * mat_B[416] +
//             mat_A[654] * mat_B[448] +
//             mat_A[655] * mat_B[480] +
//             mat_A[656] * mat_B[512] +
//             mat_A[657] * mat_B[544] +
//             mat_A[658] * mat_B[576] +
//             mat_A[659] * mat_B[608] +
//             mat_A[660] * mat_B[640] +
//             mat_A[661] * mat_B[672] +
//             mat_A[662] * mat_B[704] +
//             mat_A[663] * mat_B[736] +
//             mat_A[664] * mat_B[768] +
//             mat_A[665] * mat_B[800] +
//             mat_A[666] * mat_B[832] +
//             mat_A[667] * mat_B[864] +
//             mat_A[668] * mat_B[896] +
//             mat_A[669] * mat_B[928] +
//             mat_A[670] * mat_B[960] +
//             mat_A[671] * mat_B[992];
//  mat_C[641] <= 
//             mat_A[640] * mat_B[1] +
//             mat_A[641] * mat_B[33] +
//             mat_A[642] * mat_B[65] +
//             mat_A[643] * mat_B[97] +
//             mat_A[644] * mat_B[129] +
//             mat_A[645] * mat_B[161] +
//             mat_A[646] * mat_B[193] +
//             mat_A[647] * mat_B[225] +
//             mat_A[648] * mat_B[257] +
//             mat_A[649] * mat_B[289] +
//             mat_A[650] * mat_B[321] +
//             mat_A[651] * mat_B[353] +
//             mat_A[652] * mat_B[385] +
//             mat_A[653] * mat_B[417] +
//             mat_A[654] * mat_B[449] +
//             mat_A[655] * mat_B[481] +
//             mat_A[656] * mat_B[513] +
//             mat_A[657] * mat_B[545] +
//             mat_A[658] * mat_B[577] +
//             mat_A[659] * mat_B[609] +
//             mat_A[660] * mat_B[641] +
//             mat_A[661] * mat_B[673] +
//             mat_A[662] * mat_B[705] +
//             mat_A[663] * mat_B[737] +
//             mat_A[664] * mat_B[769] +
//             mat_A[665] * mat_B[801] +
//             mat_A[666] * mat_B[833] +
//             mat_A[667] * mat_B[865] +
//             mat_A[668] * mat_B[897] +
//             mat_A[669] * mat_B[929] +
//             mat_A[670] * mat_B[961] +
//             mat_A[671] * mat_B[993];
//  mat_C[642] <= 
//             mat_A[640] * mat_B[2] +
//             mat_A[641] * mat_B[34] +
//             mat_A[642] * mat_B[66] +
//             mat_A[643] * mat_B[98] +
//             mat_A[644] * mat_B[130] +
//             mat_A[645] * mat_B[162] +
//             mat_A[646] * mat_B[194] +
//             mat_A[647] * mat_B[226] +
//             mat_A[648] * mat_B[258] +
//             mat_A[649] * mat_B[290] +
//             mat_A[650] * mat_B[322] +
//             mat_A[651] * mat_B[354] +
//             mat_A[652] * mat_B[386] +
//             mat_A[653] * mat_B[418] +
//             mat_A[654] * mat_B[450] +
//             mat_A[655] * mat_B[482] +
//             mat_A[656] * mat_B[514] +
//             mat_A[657] * mat_B[546] +
//             mat_A[658] * mat_B[578] +
//             mat_A[659] * mat_B[610] +
//             mat_A[660] * mat_B[642] +
//             mat_A[661] * mat_B[674] +
//             mat_A[662] * mat_B[706] +
//             mat_A[663] * mat_B[738] +
//             mat_A[664] * mat_B[770] +
//             mat_A[665] * mat_B[802] +
//             mat_A[666] * mat_B[834] +
//             mat_A[667] * mat_B[866] +
//             mat_A[668] * mat_B[898] +
//             mat_A[669] * mat_B[930] +
//             mat_A[670] * mat_B[962] +
//             mat_A[671] * mat_B[994];
//  mat_C[643] <= 
//             mat_A[640] * mat_B[3] +
//             mat_A[641] * mat_B[35] +
//             mat_A[642] * mat_B[67] +
//             mat_A[643] * mat_B[99] +
//             mat_A[644] * mat_B[131] +
//             mat_A[645] * mat_B[163] +
//             mat_A[646] * mat_B[195] +
//             mat_A[647] * mat_B[227] +
//             mat_A[648] * mat_B[259] +
//             mat_A[649] * mat_B[291] +
//             mat_A[650] * mat_B[323] +
//             mat_A[651] * mat_B[355] +
//             mat_A[652] * mat_B[387] +
//             mat_A[653] * mat_B[419] +
//             mat_A[654] * mat_B[451] +
//             mat_A[655] * mat_B[483] +
//             mat_A[656] * mat_B[515] +
//             mat_A[657] * mat_B[547] +
//             mat_A[658] * mat_B[579] +
//             mat_A[659] * mat_B[611] +
//             mat_A[660] * mat_B[643] +
//             mat_A[661] * mat_B[675] +
//             mat_A[662] * mat_B[707] +
//             mat_A[663] * mat_B[739] +
//             mat_A[664] * mat_B[771] +
//             mat_A[665] * mat_B[803] +
//             mat_A[666] * mat_B[835] +
//             mat_A[667] * mat_B[867] +
//             mat_A[668] * mat_B[899] +
//             mat_A[669] * mat_B[931] +
//             mat_A[670] * mat_B[963] +
//             mat_A[671] * mat_B[995];
//  mat_C[644] <= 
//             mat_A[640] * mat_B[4] +
//             mat_A[641] * mat_B[36] +
//             mat_A[642] * mat_B[68] +
//             mat_A[643] * mat_B[100] +
//             mat_A[644] * mat_B[132] +
//             mat_A[645] * mat_B[164] +
//             mat_A[646] * mat_B[196] +
//             mat_A[647] * mat_B[228] +
//             mat_A[648] * mat_B[260] +
//             mat_A[649] * mat_B[292] +
//             mat_A[650] * mat_B[324] +
//             mat_A[651] * mat_B[356] +
//             mat_A[652] * mat_B[388] +
//             mat_A[653] * mat_B[420] +
//             mat_A[654] * mat_B[452] +
//             mat_A[655] * mat_B[484] +
//             mat_A[656] * mat_B[516] +
//             mat_A[657] * mat_B[548] +
//             mat_A[658] * mat_B[580] +
//             mat_A[659] * mat_B[612] +
//             mat_A[660] * mat_B[644] +
//             mat_A[661] * mat_B[676] +
//             mat_A[662] * mat_B[708] +
//             mat_A[663] * mat_B[740] +
//             mat_A[664] * mat_B[772] +
//             mat_A[665] * mat_B[804] +
//             mat_A[666] * mat_B[836] +
//             mat_A[667] * mat_B[868] +
//             mat_A[668] * mat_B[900] +
//             mat_A[669] * mat_B[932] +
//             mat_A[670] * mat_B[964] +
//             mat_A[671] * mat_B[996];
//  mat_C[645] <= 
//             mat_A[640] * mat_B[5] +
//             mat_A[641] * mat_B[37] +
//             mat_A[642] * mat_B[69] +
//             mat_A[643] * mat_B[101] +
//             mat_A[644] * mat_B[133] +
//             mat_A[645] * mat_B[165] +
//             mat_A[646] * mat_B[197] +
//             mat_A[647] * mat_B[229] +
//             mat_A[648] * mat_B[261] +
//             mat_A[649] * mat_B[293] +
//             mat_A[650] * mat_B[325] +
//             mat_A[651] * mat_B[357] +
//             mat_A[652] * mat_B[389] +
//             mat_A[653] * mat_B[421] +
//             mat_A[654] * mat_B[453] +
//             mat_A[655] * mat_B[485] +
//             mat_A[656] * mat_B[517] +
//             mat_A[657] * mat_B[549] +
//             mat_A[658] * mat_B[581] +
//             mat_A[659] * mat_B[613] +
//             mat_A[660] * mat_B[645] +
//             mat_A[661] * mat_B[677] +
//             mat_A[662] * mat_B[709] +
//             mat_A[663] * mat_B[741] +
//             mat_A[664] * mat_B[773] +
//             mat_A[665] * mat_B[805] +
//             mat_A[666] * mat_B[837] +
//             mat_A[667] * mat_B[869] +
//             mat_A[668] * mat_B[901] +
//             mat_A[669] * mat_B[933] +
//             mat_A[670] * mat_B[965] +
//             mat_A[671] * mat_B[997];
//  mat_C[646] <= 
//             mat_A[640] * mat_B[6] +
//             mat_A[641] * mat_B[38] +
//             mat_A[642] * mat_B[70] +
//             mat_A[643] * mat_B[102] +
//             mat_A[644] * mat_B[134] +
//             mat_A[645] * mat_B[166] +
//             mat_A[646] * mat_B[198] +
//             mat_A[647] * mat_B[230] +
//             mat_A[648] * mat_B[262] +
//             mat_A[649] * mat_B[294] +
//             mat_A[650] * mat_B[326] +
//             mat_A[651] * mat_B[358] +
//             mat_A[652] * mat_B[390] +
//             mat_A[653] * mat_B[422] +
//             mat_A[654] * mat_B[454] +
//             mat_A[655] * mat_B[486] +
//             mat_A[656] * mat_B[518] +
//             mat_A[657] * mat_B[550] +
//             mat_A[658] * mat_B[582] +
//             mat_A[659] * mat_B[614] +
//             mat_A[660] * mat_B[646] +
//             mat_A[661] * mat_B[678] +
//             mat_A[662] * mat_B[710] +
//             mat_A[663] * mat_B[742] +
//             mat_A[664] * mat_B[774] +
//             mat_A[665] * mat_B[806] +
//             mat_A[666] * mat_B[838] +
//             mat_A[667] * mat_B[870] +
//             mat_A[668] * mat_B[902] +
//             mat_A[669] * mat_B[934] +
//             mat_A[670] * mat_B[966] +
//             mat_A[671] * mat_B[998];
//  mat_C[647] <= 
//             mat_A[640] * mat_B[7] +
//             mat_A[641] * mat_B[39] +
//             mat_A[642] * mat_B[71] +
//             mat_A[643] * mat_B[103] +
//             mat_A[644] * mat_B[135] +
//             mat_A[645] * mat_B[167] +
//             mat_A[646] * mat_B[199] +
//             mat_A[647] * mat_B[231] +
//             mat_A[648] * mat_B[263] +
//             mat_A[649] * mat_B[295] +
//             mat_A[650] * mat_B[327] +
//             mat_A[651] * mat_B[359] +
//             mat_A[652] * mat_B[391] +
//             mat_A[653] * mat_B[423] +
//             mat_A[654] * mat_B[455] +
//             mat_A[655] * mat_B[487] +
//             mat_A[656] * mat_B[519] +
//             mat_A[657] * mat_B[551] +
//             mat_A[658] * mat_B[583] +
//             mat_A[659] * mat_B[615] +
//             mat_A[660] * mat_B[647] +
//             mat_A[661] * mat_B[679] +
//             mat_A[662] * mat_B[711] +
//             mat_A[663] * mat_B[743] +
//             mat_A[664] * mat_B[775] +
//             mat_A[665] * mat_B[807] +
//             mat_A[666] * mat_B[839] +
//             mat_A[667] * mat_B[871] +
//             mat_A[668] * mat_B[903] +
//             mat_A[669] * mat_B[935] +
//             mat_A[670] * mat_B[967] +
//             mat_A[671] * mat_B[999];
//  mat_C[648] <= 
//             mat_A[640] * mat_B[8] +
//             mat_A[641] * mat_B[40] +
//             mat_A[642] * mat_B[72] +
//             mat_A[643] * mat_B[104] +
//             mat_A[644] * mat_B[136] +
//             mat_A[645] * mat_B[168] +
//             mat_A[646] * mat_B[200] +
//             mat_A[647] * mat_B[232] +
//             mat_A[648] * mat_B[264] +
//             mat_A[649] * mat_B[296] +
//             mat_A[650] * mat_B[328] +
//             mat_A[651] * mat_B[360] +
//             mat_A[652] * mat_B[392] +
//             mat_A[653] * mat_B[424] +
//             mat_A[654] * mat_B[456] +
//             mat_A[655] * mat_B[488] +
//             mat_A[656] * mat_B[520] +
//             mat_A[657] * mat_B[552] +
//             mat_A[658] * mat_B[584] +
//             mat_A[659] * mat_B[616] +
//             mat_A[660] * mat_B[648] +
//             mat_A[661] * mat_B[680] +
//             mat_A[662] * mat_B[712] +
//             mat_A[663] * mat_B[744] +
//             mat_A[664] * mat_B[776] +
//             mat_A[665] * mat_B[808] +
//             mat_A[666] * mat_B[840] +
//             mat_A[667] * mat_B[872] +
//             mat_A[668] * mat_B[904] +
//             mat_A[669] * mat_B[936] +
//             mat_A[670] * mat_B[968] +
//             mat_A[671] * mat_B[1000];
//  mat_C[649] <= 
//             mat_A[640] * mat_B[9] +
//             mat_A[641] * mat_B[41] +
//             mat_A[642] * mat_B[73] +
//             mat_A[643] * mat_B[105] +
//             mat_A[644] * mat_B[137] +
//             mat_A[645] * mat_B[169] +
//             mat_A[646] * mat_B[201] +
//             mat_A[647] * mat_B[233] +
//             mat_A[648] * mat_B[265] +
//             mat_A[649] * mat_B[297] +
//             mat_A[650] * mat_B[329] +
//             mat_A[651] * mat_B[361] +
//             mat_A[652] * mat_B[393] +
//             mat_A[653] * mat_B[425] +
//             mat_A[654] * mat_B[457] +
//             mat_A[655] * mat_B[489] +
//             mat_A[656] * mat_B[521] +
//             mat_A[657] * mat_B[553] +
//             mat_A[658] * mat_B[585] +
//             mat_A[659] * mat_B[617] +
//             mat_A[660] * mat_B[649] +
//             mat_A[661] * mat_B[681] +
//             mat_A[662] * mat_B[713] +
//             mat_A[663] * mat_B[745] +
//             mat_A[664] * mat_B[777] +
//             mat_A[665] * mat_B[809] +
//             mat_A[666] * mat_B[841] +
//             mat_A[667] * mat_B[873] +
//             mat_A[668] * mat_B[905] +
//             mat_A[669] * mat_B[937] +
//             mat_A[670] * mat_B[969] +
//             mat_A[671] * mat_B[1001];
//  mat_C[650] <= 
//             mat_A[640] * mat_B[10] +
//             mat_A[641] * mat_B[42] +
//             mat_A[642] * mat_B[74] +
//             mat_A[643] * mat_B[106] +
//             mat_A[644] * mat_B[138] +
//             mat_A[645] * mat_B[170] +
//             mat_A[646] * mat_B[202] +
//             mat_A[647] * mat_B[234] +
//             mat_A[648] * mat_B[266] +
//             mat_A[649] * mat_B[298] +
//             mat_A[650] * mat_B[330] +
//             mat_A[651] * mat_B[362] +
//             mat_A[652] * mat_B[394] +
//             mat_A[653] * mat_B[426] +
//             mat_A[654] * mat_B[458] +
//             mat_A[655] * mat_B[490] +
//             mat_A[656] * mat_B[522] +
//             mat_A[657] * mat_B[554] +
//             mat_A[658] * mat_B[586] +
//             mat_A[659] * mat_B[618] +
//             mat_A[660] * mat_B[650] +
//             mat_A[661] * mat_B[682] +
//             mat_A[662] * mat_B[714] +
//             mat_A[663] * mat_B[746] +
//             mat_A[664] * mat_B[778] +
//             mat_A[665] * mat_B[810] +
//             mat_A[666] * mat_B[842] +
//             mat_A[667] * mat_B[874] +
//             mat_A[668] * mat_B[906] +
//             mat_A[669] * mat_B[938] +
//             mat_A[670] * mat_B[970] +
//             mat_A[671] * mat_B[1002];
//  mat_C[651] <= 
//             mat_A[640] * mat_B[11] +
//             mat_A[641] * mat_B[43] +
//             mat_A[642] * mat_B[75] +
//             mat_A[643] * mat_B[107] +
//             mat_A[644] * mat_B[139] +
//             mat_A[645] * mat_B[171] +
//             mat_A[646] * mat_B[203] +
//             mat_A[647] * mat_B[235] +
//             mat_A[648] * mat_B[267] +
//             mat_A[649] * mat_B[299] +
//             mat_A[650] * mat_B[331] +
//             mat_A[651] * mat_B[363] +
//             mat_A[652] * mat_B[395] +
//             mat_A[653] * mat_B[427] +
//             mat_A[654] * mat_B[459] +
//             mat_A[655] * mat_B[491] +
//             mat_A[656] * mat_B[523] +
//             mat_A[657] * mat_B[555] +
//             mat_A[658] * mat_B[587] +
//             mat_A[659] * mat_B[619] +
//             mat_A[660] * mat_B[651] +
//             mat_A[661] * mat_B[683] +
//             mat_A[662] * mat_B[715] +
//             mat_A[663] * mat_B[747] +
//             mat_A[664] * mat_B[779] +
//             mat_A[665] * mat_B[811] +
//             mat_A[666] * mat_B[843] +
//             mat_A[667] * mat_B[875] +
//             mat_A[668] * mat_B[907] +
//             mat_A[669] * mat_B[939] +
//             mat_A[670] * mat_B[971] +
//             mat_A[671] * mat_B[1003];
//  mat_C[652] <= 
//             mat_A[640] * mat_B[12] +
//             mat_A[641] * mat_B[44] +
//             mat_A[642] * mat_B[76] +
//             mat_A[643] * mat_B[108] +
//             mat_A[644] * mat_B[140] +
//             mat_A[645] * mat_B[172] +
//             mat_A[646] * mat_B[204] +
//             mat_A[647] * mat_B[236] +
//             mat_A[648] * mat_B[268] +
//             mat_A[649] * mat_B[300] +
//             mat_A[650] * mat_B[332] +
//             mat_A[651] * mat_B[364] +
//             mat_A[652] * mat_B[396] +
//             mat_A[653] * mat_B[428] +
//             mat_A[654] * mat_B[460] +
//             mat_A[655] * mat_B[492] +
//             mat_A[656] * mat_B[524] +
//             mat_A[657] * mat_B[556] +
//             mat_A[658] * mat_B[588] +
//             mat_A[659] * mat_B[620] +
//             mat_A[660] * mat_B[652] +
//             mat_A[661] * mat_B[684] +
//             mat_A[662] * mat_B[716] +
//             mat_A[663] * mat_B[748] +
//             mat_A[664] * mat_B[780] +
//             mat_A[665] * mat_B[812] +
//             mat_A[666] * mat_B[844] +
//             mat_A[667] * mat_B[876] +
//             mat_A[668] * mat_B[908] +
//             mat_A[669] * mat_B[940] +
//             mat_A[670] * mat_B[972] +
//             mat_A[671] * mat_B[1004];
//  mat_C[653] <= 
//             mat_A[640] * mat_B[13] +
//             mat_A[641] * mat_B[45] +
//             mat_A[642] * mat_B[77] +
//             mat_A[643] * mat_B[109] +
//             mat_A[644] * mat_B[141] +
//             mat_A[645] * mat_B[173] +
//             mat_A[646] * mat_B[205] +
//             mat_A[647] * mat_B[237] +
//             mat_A[648] * mat_B[269] +
//             mat_A[649] * mat_B[301] +
//             mat_A[650] * mat_B[333] +
//             mat_A[651] * mat_B[365] +
//             mat_A[652] * mat_B[397] +
//             mat_A[653] * mat_B[429] +
//             mat_A[654] * mat_B[461] +
//             mat_A[655] * mat_B[493] +
//             mat_A[656] * mat_B[525] +
//             mat_A[657] * mat_B[557] +
//             mat_A[658] * mat_B[589] +
//             mat_A[659] * mat_B[621] +
//             mat_A[660] * mat_B[653] +
//             mat_A[661] * mat_B[685] +
//             mat_A[662] * mat_B[717] +
//             mat_A[663] * mat_B[749] +
//             mat_A[664] * mat_B[781] +
//             mat_A[665] * mat_B[813] +
//             mat_A[666] * mat_B[845] +
//             mat_A[667] * mat_B[877] +
//             mat_A[668] * mat_B[909] +
//             mat_A[669] * mat_B[941] +
//             mat_A[670] * mat_B[973] +
//             mat_A[671] * mat_B[1005];
//  mat_C[654] <= 
//             mat_A[640] * mat_B[14] +
//             mat_A[641] * mat_B[46] +
//             mat_A[642] * mat_B[78] +
//             mat_A[643] * mat_B[110] +
//             mat_A[644] * mat_B[142] +
//             mat_A[645] * mat_B[174] +
//             mat_A[646] * mat_B[206] +
//             mat_A[647] * mat_B[238] +
//             mat_A[648] * mat_B[270] +
//             mat_A[649] * mat_B[302] +
//             mat_A[650] * mat_B[334] +
//             mat_A[651] * mat_B[366] +
//             mat_A[652] * mat_B[398] +
//             mat_A[653] * mat_B[430] +
//             mat_A[654] * mat_B[462] +
//             mat_A[655] * mat_B[494] +
//             mat_A[656] * mat_B[526] +
//             mat_A[657] * mat_B[558] +
//             mat_A[658] * mat_B[590] +
//             mat_A[659] * mat_B[622] +
//             mat_A[660] * mat_B[654] +
//             mat_A[661] * mat_B[686] +
//             mat_A[662] * mat_B[718] +
//             mat_A[663] * mat_B[750] +
//             mat_A[664] * mat_B[782] +
//             mat_A[665] * mat_B[814] +
//             mat_A[666] * mat_B[846] +
//             mat_A[667] * mat_B[878] +
//             mat_A[668] * mat_B[910] +
//             mat_A[669] * mat_B[942] +
//             mat_A[670] * mat_B[974] +
//             mat_A[671] * mat_B[1006];
//  mat_C[655] <= 
//             mat_A[640] * mat_B[15] +
//             mat_A[641] * mat_B[47] +
//             mat_A[642] * mat_B[79] +
//             mat_A[643] * mat_B[111] +
//             mat_A[644] * mat_B[143] +
//             mat_A[645] * mat_B[175] +
//             mat_A[646] * mat_B[207] +
//             mat_A[647] * mat_B[239] +
//             mat_A[648] * mat_B[271] +
//             mat_A[649] * mat_B[303] +
//             mat_A[650] * mat_B[335] +
//             mat_A[651] * mat_B[367] +
//             mat_A[652] * mat_B[399] +
//             mat_A[653] * mat_B[431] +
//             mat_A[654] * mat_B[463] +
//             mat_A[655] * mat_B[495] +
//             mat_A[656] * mat_B[527] +
//             mat_A[657] * mat_B[559] +
//             mat_A[658] * mat_B[591] +
//             mat_A[659] * mat_B[623] +
//             mat_A[660] * mat_B[655] +
//             mat_A[661] * mat_B[687] +
//             mat_A[662] * mat_B[719] +
//             mat_A[663] * mat_B[751] +
//             mat_A[664] * mat_B[783] +
//             mat_A[665] * mat_B[815] +
//             mat_A[666] * mat_B[847] +
//             mat_A[667] * mat_B[879] +
//             mat_A[668] * mat_B[911] +
//             mat_A[669] * mat_B[943] +
//             mat_A[670] * mat_B[975] +
//             mat_A[671] * mat_B[1007];
//  mat_C[656] <= 
//             mat_A[640] * mat_B[16] +
//             mat_A[641] * mat_B[48] +
//             mat_A[642] * mat_B[80] +
//             mat_A[643] * mat_B[112] +
//             mat_A[644] * mat_B[144] +
//             mat_A[645] * mat_B[176] +
//             mat_A[646] * mat_B[208] +
//             mat_A[647] * mat_B[240] +
//             mat_A[648] * mat_B[272] +
//             mat_A[649] * mat_B[304] +
//             mat_A[650] * mat_B[336] +
//             mat_A[651] * mat_B[368] +
//             mat_A[652] * mat_B[400] +
//             mat_A[653] * mat_B[432] +
//             mat_A[654] * mat_B[464] +
//             mat_A[655] * mat_B[496] +
//             mat_A[656] * mat_B[528] +
//             mat_A[657] * mat_B[560] +
//             mat_A[658] * mat_B[592] +
//             mat_A[659] * mat_B[624] +
//             mat_A[660] * mat_B[656] +
//             mat_A[661] * mat_B[688] +
//             mat_A[662] * mat_B[720] +
//             mat_A[663] * mat_B[752] +
//             mat_A[664] * mat_B[784] +
//             mat_A[665] * mat_B[816] +
//             mat_A[666] * mat_B[848] +
//             mat_A[667] * mat_B[880] +
//             mat_A[668] * mat_B[912] +
//             mat_A[669] * mat_B[944] +
//             mat_A[670] * mat_B[976] +
//             mat_A[671] * mat_B[1008];
//  mat_C[657] <= 
//             mat_A[640] * mat_B[17] +
//             mat_A[641] * mat_B[49] +
//             mat_A[642] * mat_B[81] +
//             mat_A[643] * mat_B[113] +
//             mat_A[644] * mat_B[145] +
//             mat_A[645] * mat_B[177] +
//             mat_A[646] * mat_B[209] +
//             mat_A[647] * mat_B[241] +
//             mat_A[648] * mat_B[273] +
//             mat_A[649] * mat_B[305] +
//             mat_A[650] * mat_B[337] +
//             mat_A[651] * mat_B[369] +
//             mat_A[652] * mat_B[401] +
//             mat_A[653] * mat_B[433] +
//             mat_A[654] * mat_B[465] +
//             mat_A[655] * mat_B[497] +
//             mat_A[656] * mat_B[529] +
//             mat_A[657] * mat_B[561] +
//             mat_A[658] * mat_B[593] +
//             mat_A[659] * mat_B[625] +
//             mat_A[660] * mat_B[657] +
//             mat_A[661] * mat_B[689] +
//             mat_A[662] * mat_B[721] +
//             mat_A[663] * mat_B[753] +
//             mat_A[664] * mat_B[785] +
//             mat_A[665] * mat_B[817] +
//             mat_A[666] * mat_B[849] +
//             mat_A[667] * mat_B[881] +
//             mat_A[668] * mat_B[913] +
//             mat_A[669] * mat_B[945] +
//             mat_A[670] * mat_B[977] +
//             mat_A[671] * mat_B[1009];
//  mat_C[658] <= 
//             mat_A[640] * mat_B[18] +
//             mat_A[641] * mat_B[50] +
//             mat_A[642] * mat_B[82] +
//             mat_A[643] * mat_B[114] +
//             mat_A[644] * mat_B[146] +
//             mat_A[645] * mat_B[178] +
//             mat_A[646] * mat_B[210] +
//             mat_A[647] * mat_B[242] +
//             mat_A[648] * mat_B[274] +
//             mat_A[649] * mat_B[306] +
//             mat_A[650] * mat_B[338] +
//             mat_A[651] * mat_B[370] +
//             mat_A[652] * mat_B[402] +
//             mat_A[653] * mat_B[434] +
//             mat_A[654] * mat_B[466] +
//             mat_A[655] * mat_B[498] +
//             mat_A[656] * mat_B[530] +
//             mat_A[657] * mat_B[562] +
//             mat_A[658] * mat_B[594] +
//             mat_A[659] * mat_B[626] +
//             mat_A[660] * mat_B[658] +
//             mat_A[661] * mat_B[690] +
//             mat_A[662] * mat_B[722] +
//             mat_A[663] * mat_B[754] +
//             mat_A[664] * mat_B[786] +
//             mat_A[665] * mat_B[818] +
//             mat_A[666] * mat_B[850] +
//             mat_A[667] * mat_B[882] +
//             mat_A[668] * mat_B[914] +
//             mat_A[669] * mat_B[946] +
//             mat_A[670] * mat_B[978] +
//             mat_A[671] * mat_B[1010];
//  mat_C[659] <= 
//             mat_A[640] * mat_B[19] +
//             mat_A[641] * mat_B[51] +
//             mat_A[642] * mat_B[83] +
//             mat_A[643] * mat_B[115] +
//             mat_A[644] * mat_B[147] +
//             mat_A[645] * mat_B[179] +
//             mat_A[646] * mat_B[211] +
//             mat_A[647] * mat_B[243] +
//             mat_A[648] * mat_B[275] +
//             mat_A[649] * mat_B[307] +
//             mat_A[650] * mat_B[339] +
//             mat_A[651] * mat_B[371] +
//             mat_A[652] * mat_B[403] +
//             mat_A[653] * mat_B[435] +
//             mat_A[654] * mat_B[467] +
//             mat_A[655] * mat_B[499] +
//             mat_A[656] * mat_B[531] +
//             mat_A[657] * mat_B[563] +
//             mat_A[658] * mat_B[595] +
//             mat_A[659] * mat_B[627] +
//             mat_A[660] * mat_B[659] +
//             mat_A[661] * mat_B[691] +
//             mat_A[662] * mat_B[723] +
//             mat_A[663] * mat_B[755] +
//             mat_A[664] * mat_B[787] +
//             mat_A[665] * mat_B[819] +
//             mat_A[666] * mat_B[851] +
//             mat_A[667] * mat_B[883] +
//             mat_A[668] * mat_B[915] +
//             mat_A[669] * mat_B[947] +
//             mat_A[670] * mat_B[979] +
//             mat_A[671] * mat_B[1011];
//  mat_C[660] <= 
//             mat_A[640] * mat_B[20] +
//             mat_A[641] * mat_B[52] +
//             mat_A[642] * mat_B[84] +
//             mat_A[643] * mat_B[116] +
//             mat_A[644] * mat_B[148] +
//             mat_A[645] * mat_B[180] +
//             mat_A[646] * mat_B[212] +
//             mat_A[647] * mat_B[244] +
//             mat_A[648] * mat_B[276] +
//             mat_A[649] * mat_B[308] +
//             mat_A[650] * mat_B[340] +
//             mat_A[651] * mat_B[372] +
//             mat_A[652] * mat_B[404] +
//             mat_A[653] * mat_B[436] +
//             mat_A[654] * mat_B[468] +
//             mat_A[655] * mat_B[500] +
//             mat_A[656] * mat_B[532] +
//             mat_A[657] * mat_B[564] +
//             mat_A[658] * mat_B[596] +
//             mat_A[659] * mat_B[628] +
//             mat_A[660] * mat_B[660] +
//             mat_A[661] * mat_B[692] +
//             mat_A[662] * mat_B[724] +
//             mat_A[663] * mat_B[756] +
//             mat_A[664] * mat_B[788] +
//             mat_A[665] * mat_B[820] +
//             mat_A[666] * mat_B[852] +
//             mat_A[667] * mat_B[884] +
//             mat_A[668] * mat_B[916] +
//             mat_A[669] * mat_B[948] +
//             mat_A[670] * mat_B[980] +
//             mat_A[671] * mat_B[1012];
//  mat_C[661] <= 
//             mat_A[640] * mat_B[21] +
//             mat_A[641] * mat_B[53] +
//             mat_A[642] * mat_B[85] +
//             mat_A[643] * mat_B[117] +
//             mat_A[644] * mat_B[149] +
//             mat_A[645] * mat_B[181] +
//             mat_A[646] * mat_B[213] +
//             mat_A[647] * mat_B[245] +
//             mat_A[648] * mat_B[277] +
//             mat_A[649] * mat_B[309] +
//             mat_A[650] * mat_B[341] +
//             mat_A[651] * mat_B[373] +
//             mat_A[652] * mat_B[405] +
//             mat_A[653] * mat_B[437] +
//             mat_A[654] * mat_B[469] +
//             mat_A[655] * mat_B[501] +
//             mat_A[656] * mat_B[533] +
//             mat_A[657] * mat_B[565] +
//             mat_A[658] * mat_B[597] +
//             mat_A[659] * mat_B[629] +
//             mat_A[660] * mat_B[661] +
//             mat_A[661] * mat_B[693] +
//             mat_A[662] * mat_B[725] +
//             mat_A[663] * mat_B[757] +
//             mat_A[664] * mat_B[789] +
//             mat_A[665] * mat_B[821] +
//             mat_A[666] * mat_B[853] +
//             mat_A[667] * mat_B[885] +
//             mat_A[668] * mat_B[917] +
//             mat_A[669] * mat_B[949] +
//             mat_A[670] * mat_B[981] +
//             mat_A[671] * mat_B[1013];
//  mat_C[662] <= 
//             mat_A[640] * mat_B[22] +
//             mat_A[641] * mat_B[54] +
//             mat_A[642] * mat_B[86] +
//             mat_A[643] * mat_B[118] +
//             mat_A[644] * mat_B[150] +
//             mat_A[645] * mat_B[182] +
//             mat_A[646] * mat_B[214] +
//             mat_A[647] * mat_B[246] +
//             mat_A[648] * mat_B[278] +
//             mat_A[649] * mat_B[310] +
//             mat_A[650] * mat_B[342] +
//             mat_A[651] * mat_B[374] +
//             mat_A[652] * mat_B[406] +
//             mat_A[653] * mat_B[438] +
//             mat_A[654] * mat_B[470] +
//             mat_A[655] * mat_B[502] +
//             mat_A[656] * mat_B[534] +
//             mat_A[657] * mat_B[566] +
//             mat_A[658] * mat_B[598] +
//             mat_A[659] * mat_B[630] +
//             mat_A[660] * mat_B[662] +
//             mat_A[661] * mat_B[694] +
//             mat_A[662] * mat_B[726] +
//             mat_A[663] * mat_B[758] +
//             mat_A[664] * mat_B[790] +
//             mat_A[665] * mat_B[822] +
//             mat_A[666] * mat_B[854] +
//             mat_A[667] * mat_B[886] +
//             mat_A[668] * mat_B[918] +
//             mat_A[669] * mat_B[950] +
//             mat_A[670] * mat_B[982] +
//             mat_A[671] * mat_B[1014];
//  mat_C[663] <= 
//             mat_A[640] * mat_B[23] +
//             mat_A[641] * mat_B[55] +
//             mat_A[642] * mat_B[87] +
//             mat_A[643] * mat_B[119] +
//             mat_A[644] * mat_B[151] +
//             mat_A[645] * mat_B[183] +
//             mat_A[646] * mat_B[215] +
//             mat_A[647] * mat_B[247] +
//             mat_A[648] * mat_B[279] +
//             mat_A[649] * mat_B[311] +
//             mat_A[650] * mat_B[343] +
//             mat_A[651] * mat_B[375] +
//             mat_A[652] * mat_B[407] +
//             mat_A[653] * mat_B[439] +
//             mat_A[654] * mat_B[471] +
//             mat_A[655] * mat_B[503] +
//             mat_A[656] * mat_B[535] +
//             mat_A[657] * mat_B[567] +
//             mat_A[658] * mat_B[599] +
//             mat_A[659] * mat_B[631] +
//             mat_A[660] * mat_B[663] +
//             mat_A[661] * mat_B[695] +
//             mat_A[662] * mat_B[727] +
//             mat_A[663] * mat_B[759] +
//             mat_A[664] * mat_B[791] +
//             mat_A[665] * mat_B[823] +
//             mat_A[666] * mat_B[855] +
//             mat_A[667] * mat_B[887] +
//             mat_A[668] * mat_B[919] +
//             mat_A[669] * mat_B[951] +
//             mat_A[670] * mat_B[983] +
//             mat_A[671] * mat_B[1015];
//  mat_C[664] <= 
//             mat_A[640] * mat_B[24] +
//             mat_A[641] * mat_B[56] +
//             mat_A[642] * mat_B[88] +
//             mat_A[643] * mat_B[120] +
//             mat_A[644] * mat_B[152] +
//             mat_A[645] * mat_B[184] +
//             mat_A[646] * mat_B[216] +
//             mat_A[647] * mat_B[248] +
//             mat_A[648] * mat_B[280] +
//             mat_A[649] * mat_B[312] +
//             mat_A[650] * mat_B[344] +
//             mat_A[651] * mat_B[376] +
//             mat_A[652] * mat_B[408] +
//             mat_A[653] * mat_B[440] +
//             mat_A[654] * mat_B[472] +
//             mat_A[655] * mat_B[504] +
//             mat_A[656] * mat_B[536] +
//             mat_A[657] * mat_B[568] +
//             mat_A[658] * mat_B[600] +
//             mat_A[659] * mat_B[632] +
//             mat_A[660] * mat_B[664] +
//             mat_A[661] * mat_B[696] +
//             mat_A[662] * mat_B[728] +
//             mat_A[663] * mat_B[760] +
//             mat_A[664] * mat_B[792] +
//             mat_A[665] * mat_B[824] +
//             mat_A[666] * mat_B[856] +
//             mat_A[667] * mat_B[888] +
//             mat_A[668] * mat_B[920] +
//             mat_A[669] * mat_B[952] +
//             mat_A[670] * mat_B[984] +
//             mat_A[671] * mat_B[1016];
//  mat_C[665] <= 
//             mat_A[640] * mat_B[25] +
//             mat_A[641] * mat_B[57] +
//             mat_A[642] * mat_B[89] +
//             mat_A[643] * mat_B[121] +
//             mat_A[644] * mat_B[153] +
//             mat_A[645] * mat_B[185] +
//             mat_A[646] * mat_B[217] +
//             mat_A[647] * mat_B[249] +
//             mat_A[648] * mat_B[281] +
//             mat_A[649] * mat_B[313] +
//             mat_A[650] * mat_B[345] +
//             mat_A[651] * mat_B[377] +
//             mat_A[652] * mat_B[409] +
//             mat_A[653] * mat_B[441] +
//             mat_A[654] * mat_B[473] +
//             mat_A[655] * mat_B[505] +
//             mat_A[656] * mat_B[537] +
//             mat_A[657] * mat_B[569] +
//             mat_A[658] * mat_B[601] +
//             mat_A[659] * mat_B[633] +
//             mat_A[660] * mat_B[665] +
//             mat_A[661] * mat_B[697] +
//             mat_A[662] * mat_B[729] +
//             mat_A[663] * mat_B[761] +
//             mat_A[664] * mat_B[793] +
//             mat_A[665] * mat_B[825] +
//             mat_A[666] * mat_B[857] +
//             mat_A[667] * mat_B[889] +
//             mat_A[668] * mat_B[921] +
//             mat_A[669] * mat_B[953] +
//             mat_A[670] * mat_B[985] +
//             mat_A[671] * mat_B[1017];
//  mat_C[666] <= 
//             mat_A[640] * mat_B[26] +
//             mat_A[641] * mat_B[58] +
//             mat_A[642] * mat_B[90] +
//             mat_A[643] * mat_B[122] +
//             mat_A[644] * mat_B[154] +
//             mat_A[645] * mat_B[186] +
//             mat_A[646] * mat_B[218] +
//             mat_A[647] * mat_B[250] +
//             mat_A[648] * mat_B[282] +
//             mat_A[649] * mat_B[314] +
//             mat_A[650] * mat_B[346] +
//             mat_A[651] * mat_B[378] +
//             mat_A[652] * mat_B[410] +
//             mat_A[653] * mat_B[442] +
//             mat_A[654] * mat_B[474] +
//             mat_A[655] * mat_B[506] +
//             mat_A[656] * mat_B[538] +
//             mat_A[657] * mat_B[570] +
//             mat_A[658] * mat_B[602] +
//             mat_A[659] * mat_B[634] +
//             mat_A[660] * mat_B[666] +
//             mat_A[661] * mat_B[698] +
//             mat_A[662] * mat_B[730] +
//             mat_A[663] * mat_B[762] +
//             mat_A[664] * mat_B[794] +
//             mat_A[665] * mat_B[826] +
//             mat_A[666] * mat_B[858] +
//             mat_A[667] * mat_B[890] +
//             mat_A[668] * mat_B[922] +
//             mat_A[669] * mat_B[954] +
//             mat_A[670] * mat_B[986] +
//             mat_A[671] * mat_B[1018];
//  mat_C[667] <= 
//             mat_A[640] * mat_B[27] +
//             mat_A[641] * mat_B[59] +
//             mat_A[642] * mat_B[91] +
//             mat_A[643] * mat_B[123] +
//             mat_A[644] * mat_B[155] +
//             mat_A[645] * mat_B[187] +
//             mat_A[646] * mat_B[219] +
//             mat_A[647] * mat_B[251] +
//             mat_A[648] * mat_B[283] +
//             mat_A[649] * mat_B[315] +
//             mat_A[650] * mat_B[347] +
//             mat_A[651] * mat_B[379] +
//             mat_A[652] * mat_B[411] +
//             mat_A[653] * mat_B[443] +
//             mat_A[654] * mat_B[475] +
//             mat_A[655] * mat_B[507] +
//             mat_A[656] * mat_B[539] +
//             mat_A[657] * mat_B[571] +
//             mat_A[658] * mat_B[603] +
//             mat_A[659] * mat_B[635] +
//             mat_A[660] * mat_B[667] +
//             mat_A[661] * mat_B[699] +
//             mat_A[662] * mat_B[731] +
//             mat_A[663] * mat_B[763] +
//             mat_A[664] * mat_B[795] +
//             mat_A[665] * mat_B[827] +
//             mat_A[666] * mat_B[859] +
//             mat_A[667] * mat_B[891] +
//             mat_A[668] * mat_B[923] +
//             mat_A[669] * mat_B[955] +
//             mat_A[670] * mat_B[987] +
//             mat_A[671] * mat_B[1019];
//  mat_C[668] <= 
//             mat_A[640] * mat_B[28] +
//             mat_A[641] * mat_B[60] +
//             mat_A[642] * mat_B[92] +
//             mat_A[643] * mat_B[124] +
//             mat_A[644] * mat_B[156] +
//             mat_A[645] * mat_B[188] +
//             mat_A[646] * mat_B[220] +
//             mat_A[647] * mat_B[252] +
//             mat_A[648] * mat_B[284] +
//             mat_A[649] * mat_B[316] +
//             mat_A[650] * mat_B[348] +
//             mat_A[651] * mat_B[380] +
//             mat_A[652] * mat_B[412] +
//             mat_A[653] * mat_B[444] +
//             mat_A[654] * mat_B[476] +
//             mat_A[655] * mat_B[508] +
//             mat_A[656] * mat_B[540] +
//             mat_A[657] * mat_B[572] +
//             mat_A[658] * mat_B[604] +
//             mat_A[659] * mat_B[636] +
//             mat_A[660] * mat_B[668] +
//             mat_A[661] * mat_B[700] +
//             mat_A[662] * mat_B[732] +
//             mat_A[663] * mat_B[764] +
//             mat_A[664] * mat_B[796] +
//             mat_A[665] * mat_B[828] +
//             mat_A[666] * mat_B[860] +
//             mat_A[667] * mat_B[892] +
//             mat_A[668] * mat_B[924] +
//             mat_A[669] * mat_B[956] +
//             mat_A[670] * mat_B[988] +
//             mat_A[671] * mat_B[1020];
//  mat_C[669] <= 
//             mat_A[640] * mat_B[29] +
//             mat_A[641] * mat_B[61] +
//             mat_A[642] * mat_B[93] +
//             mat_A[643] * mat_B[125] +
//             mat_A[644] * mat_B[157] +
//             mat_A[645] * mat_B[189] +
//             mat_A[646] * mat_B[221] +
//             mat_A[647] * mat_B[253] +
//             mat_A[648] * mat_B[285] +
//             mat_A[649] * mat_B[317] +
//             mat_A[650] * mat_B[349] +
//             mat_A[651] * mat_B[381] +
//             mat_A[652] * mat_B[413] +
//             mat_A[653] * mat_B[445] +
//             mat_A[654] * mat_B[477] +
//             mat_A[655] * mat_B[509] +
//             mat_A[656] * mat_B[541] +
//             mat_A[657] * mat_B[573] +
//             mat_A[658] * mat_B[605] +
//             mat_A[659] * mat_B[637] +
//             mat_A[660] * mat_B[669] +
//             mat_A[661] * mat_B[701] +
//             mat_A[662] * mat_B[733] +
//             mat_A[663] * mat_B[765] +
//             mat_A[664] * mat_B[797] +
//             mat_A[665] * mat_B[829] +
//             mat_A[666] * mat_B[861] +
//             mat_A[667] * mat_B[893] +
//             mat_A[668] * mat_B[925] +
//             mat_A[669] * mat_B[957] +
//             mat_A[670] * mat_B[989] +
//             mat_A[671] * mat_B[1021];
//  mat_C[670] <= 
//             mat_A[640] * mat_B[30] +
//             mat_A[641] * mat_B[62] +
//             mat_A[642] * mat_B[94] +
//             mat_A[643] * mat_B[126] +
//             mat_A[644] * mat_B[158] +
//             mat_A[645] * mat_B[190] +
//             mat_A[646] * mat_B[222] +
//             mat_A[647] * mat_B[254] +
//             mat_A[648] * mat_B[286] +
//             mat_A[649] * mat_B[318] +
//             mat_A[650] * mat_B[350] +
//             mat_A[651] * mat_B[382] +
//             mat_A[652] * mat_B[414] +
//             mat_A[653] * mat_B[446] +
//             mat_A[654] * mat_B[478] +
//             mat_A[655] * mat_B[510] +
//             mat_A[656] * mat_B[542] +
//             mat_A[657] * mat_B[574] +
//             mat_A[658] * mat_B[606] +
//             mat_A[659] * mat_B[638] +
//             mat_A[660] * mat_B[670] +
//             mat_A[661] * mat_B[702] +
//             mat_A[662] * mat_B[734] +
//             mat_A[663] * mat_B[766] +
//             mat_A[664] * mat_B[798] +
//             mat_A[665] * mat_B[830] +
//             mat_A[666] * mat_B[862] +
//             mat_A[667] * mat_B[894] +
//             mat_A[668] * mat_B[926] +
//             mat_A[669] * mat_B[958] +
//             mat_A[670] * mat_B[990] +
//             mat_A[671] * mat_B[1022];
//  mat_C[671] <= 
//             mat_A[640] * mat_B[31] +
//             mat_A[641] * mat_B[63] +
//             mat_A[642] * mat_B[95] +
//             mat_A[643] * mat_B[127] +
//             mat_A[644] * mat_B[159] +
//             mat_A[645] * mat_B[191] +
//             mat_A[646] * mat_B[223] +
//             mat_A[647] * mat_B[255] +
//             mat_A[648] * mat_B[287] +
//             mat_A[649] * mat_B[319] +
//             mat_A[650] * mat_B[351] +
//             mat_A[651] * mat_B[383] +
//             mat_A[652] * mat_B[415] +
//             mat_A[653] * mat_B[447] +
//             mat_A[654] * mat_B[479] +
//             mat_A[655] * mat_B[511] +
//             mat_A[656] * mat_B[543] +
//             mat_A[657] * mat_B[575] +
//             mat_A[658] * mat_B[607] +
//             mat_A[659] * mat_B[639] +
//             mat_A[660] * mat_B[671] +
//             mat_A[661] * mat_B[703] +
//             mat_A[662] * mat_B[735] +
//             mat_A[663] * mat_B[767] +
//             mat_A[664] * mat_B[799] +
//             mat_A[665] * mat_B[831] +
//             mat_A[666] * mat_B[863] +
//             mat_A[667] * mat_B[895] +
//             mat_A[668] * mat_B[927] +
//             mat_A[669] * mat_B[959] +
//             mat_A[670] * mat_B[991] +
//             mat_A[671] * mat_B[1023];
//  mat_C[672] <= 
//             mat_A[672] * mat_B[0] +
//             mat_A[673] * mat_B[32] +
//             mat_A[674] * mat_B[64] +
//             mat_A[675] * mat_B[96] +
//             mat_A[676] * mat_B[128] +
//             mat_A[677] * mat_B[160] +
//             mat_A[678] * mat_B[192] +
//             mat_A[679] * mat_B[224] +
//             mat_A[680] * mat_B[256] +
//             mat_A[681] * mat_B[288] +
//             mat_A[682] * mat_B[320] +
//             mat_A[683] * mat_B[352] +
//             mat_A[684] * mat_B[384] +
//             mat_A[685] * mat_B[416] +
//             mat_A[686] * mat_B[448] +
//             mat_A[687] * mat_B[480] +
//             mat_A[688] * mat_B[512] +
//             mat_A[689] * mat_B[544] +
//             mat_A[690] * mat_B[576] +
//             mat_A[691] * mat_B[608] +
//             mat_A[692] * mat_B[640] +
//             mat_A[693] * mat_B[672] +
//             mat_A[694] * mat_B[704] +
//             mat_A[695] * mat_B[736] +
//             mat_A[696] * mat_B[768] +
//             mat_A[697] * mat_B[800] +
//             mat_A[698] * mat_B[832] +
//             mat_A[699] * mat_B[864] +
//             mat_A[700] * mat_B[896] +
//             mat_A[701] * mat_B[928] +
//             mat_A[702] * mat_B[960] +
//             mat_A[703] * mat_B[992];
//  mat_C[673] <= 
//             mat_A[672] * mat_B[1] +
//             mat_A[673] * mat_B[33] +
//             mat_A[674] * mat_B[65] +
//             mat_A[675] * mat_B[97] +
//             mat_A[676] * mat_B[129] +
//             mat_A[677] * mat_B[161] +
//             mat_A[678] * mat_B[193] +
//             mat_A[679] * mat_B[225] +
//             mat_A[680] * mat_B[257] +
//             mat_A[681] * mat_B[289] +
//             mat_A[682] * mat_B[321] +
//             mat_A[683] * mat_B[353] +
//             mat_A[684] * mat_B[385] +
//             mat_A[685] * mat_B[417] +
//             mat_A[686] * mat_B[449] +
//             mat_A[687] * mat_B[481] +
//             mat_A[688] * mat_B[513] +
//             mat_A[689] * mat_B[545] +
//             mat_A[690] * mat_B[577] +
//             mat_A[691] * mat_B[609] +
//             mat_A[692] * mat_B[641] +
//             mat_A[693] * mat_B[673] +
//             mat_A[694] * mat_B[705] +
//             mat_A[695] * mat_B[737] +
//             mat_A[696] * mat_B[769] +
//             mat_A[697] * mat_B[801] +
//             mat_A[698] * mat_B[833] +
//             mat_A[699] * mat_B[865] +
//             mat_A[700] * mat_B[897] +
//             mat_A[701] * mat_B[929] +
//             mat_A[702] * mat_B[961] +
//             mat_A[703] * mat_B[993];
//  mat_C[674] <= 
//             mat_A[672] * mat_B[2] +
//             mat_A[673] * mat_B[34] +
//             mat_A[674] * mat_B[66] +
//             mat_A[675] * mat_B[98] +
//             mat_A[676] * mat_B[130] +
//             mat_A[677] * mat_B[162] +
//             mat_A[678] * mat_B[194] +
//             mat_A[679] * mat_B[226] +
//             mat_A[680] * mat_B[258] +
//             mat_A[681] * mat_B[290] +
//             mat_A[682] * mat_B[322] +
//             mat_A[683] * mat_B[354] +
//             mat_A[684] * mat_B[386] +
//             mat_A[685] * mat_B[418] +
//             mat_A[686] * mat_B[450] +
//             mat_A[687] * mat_B[482] +
//             mat_A[688] * mat_B[514] +
//             mat_A[689] * mat_B[546] +
//             mat_A[690] * mat_B[578] +
//             mat_A[691] * mat_B[610] +
//             mat_A[692] * mat_B[642] +
//             mat_A[693] * mat_B[674] +
//             mat_A[694] * mat_B[706] +
//             mat_A[695] * mat_B[738] +
//             mat_A[696] * mat_B[770] +
//             mat_A[697] * mat_B[802] +
//             mat_A[698] * mat_B[834] +
//             mat_A[699] * mat_B[866] +
//             mat_A[700] * mat_B[898] +
//             mat_A[701] * mat_B[930] +
//             mat_A[702] * mat_B[962] +
//             mat_A[703] * mat_B[994];
//  mat_C[675] <= 
//             mat_A[672] * mat_B[3] +
//             mat_A[673] * mat_B[35] +
//             mat_A[674] * mat_B[67] +
//             mat_A[675] * mat_B[99] +
//             mat_A[676] * mat_B[131] +
//             mat_A[677] * mat_B[163] +
//             mat_A[678] * mat_B[195] +
//             mat_A[679] * mat_B[227] +
//             mat_A[680] * mat_B[259] +
//             mat_A[681] * mat_B[291] +
//             mat_A[682] * mat_B[323] +
//             mat_A[683] * mat_B[355] +
//             mat_A[684] * mat_B[387] +
//             mat_A[685] * mat_B[419] +
//             mat_A[686] * mat_B[451] +
//             mat_A[687] * mat_B[483] +
//             mat_A[688] * mat_B[515] +
//             mat_A[689] * mat_B[547] +
//             mat_A[690] * mat_B[579] +
//             mat_A[691] * mat_B[611] +
//             mat_A[692] * mat_B[643] +
//             mat_A[693] * mat_B[675] +
//             mat_A[694] * mat_B[707] +
//             mat_A[695] * mat_B[739] +
//             mat_A[696] * mat_B[771] +
//             mat_A[697] * mat_B[803] +
//             mat_A[698] * mat_B[835] +
//             mat_A[699] * mat_B[867] +
//             mat_A[700] * mat_B[899] +
//             mat_A[701] * mat_B[931] +
//             mat_A[702] * mat_B[963] +
//             mat_A[703] * mat_B[995];
//  mat_C[676] <= 
//             mat_A[672] * mat_B[4] +
//             mat_A[673] * mat_B[36] +
//             mat_A[674] * mat_B[68] +
//             mat_A[675] * mat_B[100] +
//             mat_A[676] * mat_B[132] +
//             mat_A[677] * mat_B[164] +
//             mat_A[678] * mat_B[196] +
//             mat_A[679] * mat_B[228] +
//             mat_A[680] * mat_B[260] +
//             mat_A[681] * mat_B[292] +
//             mat_A[682] * mat_B[324] +
//             mat_A[683] * mat_B[356] +
//             mat_A[684] * mat_B[388] +
//             mat_A[685] * mat_B[420] +
//             mat_A[686] * mat_B[452] +
//             mat_A[687] * mat_B[484] +
//             mat_A[688] * mat_B[516] +
//             mat_A[689] * mat_B[548] +
//             mat_A[690] * mat_B[580] +
//             mat_A[691] * mat_B[612] +
//             mat_A[692] * mat_B[644] +
//             mat_A[693] * mat_B[676] +
//             mat_A[694] * mat_B[708] +
//             mat_A[695] * mat_B[740] +
//             mat_A[696] * mat_B[772] +
//             mat_A[697] * mat_B[804] +
//             mat_A[698] * mat_B[836] +
//             mat_A[699] * mat_B[868] +
//             mat_A[700] * mat_B[900] +
//             mat_A[701] * mat_B[932] +
//             mat_A[702] * mat_B[964] +
//             mat_A[703] * mat_B[996];
//  mat_C[677] <= 
//             mat_A[672] * mat_B[5] +
//             mat_A[673] * mat_B[37] +
//             mat_A[674] * mat_B[69] +
//             mat_A[675] * mat_B[101] +
//             mat_A[676] * mat_B[133] +
//             mat_A[677] * mat_B[165] +
//             mat_A[678] * mat_B[197] +
//             mat_A[679] * mat_B[229] +
//             mat_A[680] * mat_B[261] +
//             mat_A[681] * mat_B[293] +
//             mat_A[682] * mat_B[325] +
//             mat_A[683] * mat_B[357] +
//             mat_A[684] * mat_B[389] +
//             mat_A[685] * mat_B[421] +
//             mat_A[686] * mat_B[453] +
//             mat_A[687] * mat_B[485] +
//             mat_A[688] * mat_B[517] +
//             mat_A[689] * mat_B[549] +
//             mat_A[690] * mat_B[581] +
//             mat_A[691] * mat_B[613] +
//             mat_A[692] * mat_B[645] +
//             mat_A[693] * mat_B[677] +
//             mat_A[694] * mat_B[709] +
//             mat_A[695] * mat_B[741] +
//             mat_A[696] * mat_B[773] +
//             mat_A[697] * mat_B[805] +
//             mat_A[698] * mat_B[837] +
//             mat_A[699] * mat_B[869] +
//             mat_A[700] * mat_B[901] +
//             mat_A[701] * mat_B[933] +
//             mat_A[702] * mat_B[965] +
//             mat_A[703] * mat_B[997];
//  mat_C[678] <= 
//             mat_A[672] * mat_B[6] +
//             mat_A[673] * mat_B[38] +
//             mat_A[674] * mat_B[70] +
//             mat_A[675] * mat_B[102] +
//             mat_A[676] * mat_B[134] +
//             mat_A[677] * mat_B[166] +
//             mat_A[678] * mat_B[198] +
//             mat_A[679] * mat_B[230] +
//             mat_A[680] * mat_B[262] +
//             mat_A[681] * mat_B[294] +
//             mat_A[682] * mat_B[326] +
//             mat_A[683] * mat_B[358] +
//             mat_A[684] * mat_B[390] +
//             mat_A[685] * mat_B[422] +
//             mat_A[686] * mat_B[454] +
//             mat_A[687] * mat_B[486] +
//             mat_A[688] * mat_B[518] +
//             mat_A[689] * mat_B[550] +
//             mat_A[690] * mat_B[582] +
//             mat_A[691] * mat_B[614] +
//             mat_A[692] * mat_B[646] +
//             mat_A[693] * mat_B[678] +
//             mat_A[694] * mat_B[710] +
//             mat_A[695] * mat_B[742] +
//             mat_A[696] * mat_B[774] +
//             mat_A[697] * mat_B[806] +
//             mat_A[698] * mat_B[838] +
//             mat_A[699] * mat_B[870] +
//             mat_A[700] * mat_B[902] +
//             mat_A[701] * mat_B[934] +
//             mat_A[702] * mat_B[966] +
//             mat_A[703] * mat_B[998];
//  mat_C[679] <= 
//             mat_A[672] * mat_B[7] +
//             mat_A[673] * mat_B[39] +
//             mat_A[674] * mat_B[71] +
//             mat_A[675] * mat_B[103] +
//             mat_A[676] * mat_B[135] +
//             mat_A[677] * mat_B[167] +
//             mat_A[678] * mat_B[199] +
//             mat_A[679] * mat_B[231] +
//             mat_A[680] * mat_B[263] +
//             mat_A[681] * mat_B[295] +
//             mat_A[682] * mat_B[327] +
//             mat_A[683] * mat_B[359] +
//             mat_A[684] * mat_B[391] +
//             mat_A[685] * mat_B[423] +
//             mat_A[686] * mat_B[455] +
//             mat_A[687] * mat_B[487] +
//             mat_A[688] * mat_B[519] +
//             mat_A[689] * mat_B[551] +
//             mat_A[690] * mat_B[583] +
//             mat_A[691] * mat_B[615] +
//             mat_A[692] * mat_B[647] +
//             mat_A[693] * mat_B[679] +
//             mat_A[694] * mat_B[711] +
//             mat_A[695] * mat_B[743] +
//             mat_A[696] * mat_B[775] +
//             mat_A[697] * mat_B[807] +
//             mat_A[698] * mat_B[839] +
//             mat_A[699] * mat_B[871] +
//             mat_A[700] * mat_B[903] +
//             mat_A[701] * mat_B[935] +
//             mat_A[702] * mat_B[967] +
//             mat_A[703] * mat_B[999];
//  mat_C[680] <= 
//             mat_A[672] * mat_B[8] +
//             mat_A[673] * mat_B[40] +
//             mat_A[674] * mat_B[72] +
//             mat_A[675] * mat_B[104] +
//             mat_A[676] * mat_B[136] +
//             mat_A[677] * mat_B[168] +
//             mat_A[678] * mat_B[200] +
//             mat_A[679] * mat_B[232] +
//             mat_A[680] * mat_B[264] +
//             mat_A[681] * mat_B[296] +
//             mat_A[682] * mat_B[328] +
//             mat_A[683] * mat_B[360] +
//             mat_A[684] * mat_B[392] +
//             mat_A[685] * mat_B[424] +
//             mat_A[686] * mat_B[456] +
//             mat_A[687] * mat_B[488] +
//             mat_A[688] * mat_B[520] +
//             mat_A[689] * mat_B[552] +
//             mat_A[690] * mat_B[584] +
//             mat_A[691] * mat_B[616] +
//             mat_A[692] * mat_B[648] +
//             mat_A[693] * mat_B[680] +
//             mat_A[694] * mat_B[712] +
//             mat_A[695] * mat_B[744] +
//             mat_A[696] * mat_B[776] +
//             mat_A[697] * mat_B[808] +
//             mat_A[698] * mat_B[840] +
//             mat_A[699] * mat_B[872] +
//             mat_A[700] * mat_B[904] +
//             mat_A[701] * mat_B[936] +
//             mat_A[702] * mat_B[968] +
//             mat_A[703] * mat_B[1000];
//  mat_C[681] <= 
//             mat_A[672] * mat_B[9] +
//             mat_A[673] * mat_B[41] +
//             mat_A[674] * mat_B[73] +
//             mat_A[675] * mat_B[105] +
//             mat_A[676] * mat_B[137] +
//             mat_A[677] * mat_B[169] +
//             mat_A[678] * mat_B[201] +
//             mat_A[679] * mat_B[233] +
//             mat_A[680] * mat_B[265] +
//             mat_A[681] * mat_B[297] +
//             mat_A[682] * mat_B[329] +
//             mat_A[683] * mat_B[361] +
//             mat_A[684] * mat_B[393] +
//             mat_A[685] * mat_B[425] +
//             mat_A[686] * mat_B[457] +
//             mat_A[687] * mat_B[489] +
//             mat_A[688] * mat_B[521] +
//             mat_A[689] * mat_B[553] +
//             mat_A[690] * mat_B[585] +
//             mat_A[691] * mat_B[617] +
//             mat_A[692] * mat_B[649] +
//             mat_A[693] * mat_B[681] +
//             mat_A[694] * mat_B[713] +
//             mat_A[695] * mat_B[745] +
//             mat_A[696] * mat_B[777] +
//             mat_A[697] * mat_B[809] +
//             mat_A[698] * mat_B[841] +
//             mat_A[699] * mat_B[873] +
//             mat_A[700] * mat_B[905] +
//             mat_A[701] * mat_B[937] +
//             mat_A[702] * mat_B[969] +
//             mat_A[703] * mat_B[1001];
//  mat_C[682] <= 
//             mat_A[672] * mat_B[10] +
//             mat_A[673] * mat_B[42] +
//             mat_A[674] * mat_B[74] +
//             mat_A[675] * mat_B[106] +
//             mat_A[676] * mat_B[138] +
//             mat_A[677] * mat_B[170] +
//             mat_A[678] * mat_B[202] +
//             mat_A[679] * mat_B[234] +
//             mat_A[680] * mat_B[266] +
//             mat_A[681] * mat_B[298] +
//             mat_A[682] * mat_B[330] +
//             mat_A[683] * mat_B[362] +
//             mat_A[684] * mat_B[394] +
//             mat_A[685] * mat_B[426] +
//             mat_A[686] * mat_B[458] +
//             mat_A[687] * mat_B[490] +
//             mat_A[688] * mat_B[522] +
//             mat_A[689] * mat_B[554] +
//             mat_A[690] * mat_B[586] +
//             mat_A[691] * mat_B[618] +
//             mat_A[692] * mat_B[650] +
//             mat_A[693] * mat_B[682] +
//             mat_A[694] * mat_B[714] +
//             mat_A[695] * mat_B[746] +
//             mat_A[696] * mat_B[778] +
//             mat_A[697] * mat_B[810] +
//             mat_A[698] * mat_B[842] +
//             mat_A[699] * mat_B[874] +
//             mat_A[700] * mat_B[906] +
//             mat_A[701] * mat_B[938] +
//             mat_A[702] * mat_B[970] +
//             mat_A[703] * mat_B[1002];
//  mat_C[683] <= 
//             mat_A[672] * mat_B[11] +
//             mat_A[673] * mat_B[43] +
//             mat_A[674] * mat_B[75] +
//             mat_A[675] * mat_B[107] +
//             mat_A[676] * mat_B[139] +
//             mat_A[677] * mat_B[171] +
//             mat_A[678] * mat_B[203] +
//             mat_A[679] * mat_B[235] +
//             mat_A[680] * mat_B[267] +
//             mat_A[681] * mat_B[299] +
//             mat_A[682] * mat_B[331] +
//             mat_A[683] * mat_B[363] +
//             mat_A[684] * mat_B[395] +
//             mat_A[685] * mat_B[427] +
//             mat_A[686] * mat_B[459] +
//             mat_A[687] * mat_B[491] +
//             mat_A[688] * mat_B[523] +
//             mat_A[689] * mat_B[555] +
//             mat_A[690] * mat_B[587] +
//             mat_A[691] * mat_B[619] +
//             mat_A[692] * mat_B[651] +
//             mat_A[693] * mat_B[683] +
//             mat_A[694] * mat_B[715] +
//             mat_A[695] * mat_B[747] +
//             mat_A[696] * mat_B[779] +
//             mat_A[697] * mat_B[811] +
//             mat_A[698] * mat_B[843] +
//             mat_A[699] * mat_B[875] +
//             mat_A[700] * mat_B[907] +
//             mat_A[701] * mat_B[939] +
//             mat_A[702] * mat_B[971] +
//             mat_A[703] * mat_B[1003];
//  mat_C[684] <= 
//             mat_A[672] * mat_B[12] +
//             mat_A[673] * mat_B[44] +
//             mat_A[674] * mat_B[76] +
//             mat_A[675] * mat_B[108] +
//             mat_A[676] * mat_B[140] +
//             mat_A[677] * mat_B[172] +
//             mat_A[678] * mat_B[204] +
//             mat_A[679] * mat_B[236] +
//             mat_A[680] * mat_B[268] +
//             mat_A[681] * mat_B[300] +
//             mat_A[682] * mat_B[332] +
//             mat_A[683] * mat_B[364] +
//             mat_A[684] * mat_B[396] +
//             mat_A[685] * mat_B[428] +
//             mat_A[686] * mat_B[460] +
//             mat_A[687] * mat_B[492] +
//             mat_A[688] * mat_B[524] +
//             mat_A[689] * mat_B[556] +
//             mat_A[690] * mat_B[588] +
//             mat_A[691] * mat_B[620] +
//             mat_A[692] * mat_B[652] +
//             mat_A[693] * mat_B[684] +
//             mat_A[694] * mat_B[716] +
//             mat_A[695] * mat_B[748] +
//             mat_A[696] * mat_B[780] +
//             mat_A[697] * mat_B[812] +
//             mat_A[698] * mat_B[844] +
//             mat_A[699] * mat_B[876] +
//             mat_A[700] * mat_B[908] +
//             mat_A[701] * mat_B[940] +
//             mat_A[702] * mat_B[972] +
//             mat_A[703] * mat_B[1004];
//  mat_C[685] <= 
//             mat_A[672] * mat_B[13] +
//             mat_A[673] * mat_B[45] +
//             mat_A[674] * mat_B[77] +
//             mat_A[675] * mat_B[109] +
//             mat_A[676] * mat_B[141] +
//             mat_A[677] * mat_B[173] +
//             mat_A[678] * mat_B[205] +
//             mat_A[679] * mat_B[237] +
//             mat_A[680] * mat_B[269] +
//             mat_A[681] * mat_B[301] +
//             mat_A[682] * mat_B[333] +
//             mat_A[683] * mat_B[365] +
//             mat_A[684] * mat_B[397] +
//             mat_A[685] * mat_B[429] +
//             mat_A[686] * mat_B[461] +
//             mat_A[687] * mat_B[493] +
//             mat_A[688] * mat_B[525] +
//             mat_A[689] * mat_B[557] +
//             mat_A[690] * mat_B[589] +
//             mat_A[691] * mat_B[621] +
//             mat_A[692] * mat_B[653] +
//             mat_A[693] * mat_B[685] +
//             mat_A[694] * mat_B[717] +
//             mat_A[695] * mat_B[749] +
//             mat_A[696] * mat_B[781] +
//             mat_A[697] * mat_B[813] +
//             mat_A[698] * mat_B[845] +
//             mat_A[699] * mat_B[877] +
//             mat_A[700] * mat_B[909] +
//             mat_A[701] * mat_B[941] +
//             mat_A[702] * mat_B[973] +
//             mat_A[703] * mat_B[1005];
//  mat_C[686] <= 
//             mat_A[672] * mat_B[14] +
//             mat_A[673] * mat_B[46] +
//             mat_A[674] * mat_B[78] +
//             mat_A[675] * mat_B[110] +
//             mat_A[676] * mat_B[142] +
//             mat_A[677] * mat_B[174] +
//             mat_A[678] * mat_B[206] +
//             mat_A[679] * mat_B[238] +
//             mat_A[680] * mat_B[270] +
//             mat_A[681] * mat_B[302] +
//             mat_A[682] * mat_B[334] +
//             mat_A[683] * mat_B[366] +
//             mat_A[684] * mat_B[398] +
//             mat_A[685] * mat_B[430] +
//             mat_A[686] * mat_B[462] +
//             mat_A[687] * mat_B[494] +
//             mat_A[688] * mat_B[526] +
//             mat_A[689] * mat_B[558] +
//             mat_A[690] * mat_B[590] +
//             mat_A[691] * mat_B[622] +
//             mat_A[692] * mat_B[654] +
//             mat_A[693] * mat_B[686] +
//             mat_A[694] * mat_B[718] +
//             mat_A[695] * mat_B[750] +
//             mat_A[696] * mat_B[782] +
//             mat_A[697] * mat_B[814] +
//             mat_A[698] * mat_B[846] +
//             mat_A[699] * mat_B[878] +
//             mat_A[700] * mat_B[910] +
//             mat_A[701] * mat_B[942] +
//             mat_A[702] * mat_B[974] +
//             mat_A[703] * mat_B[1006];
//  mat_C[687] <= 
//             mat_A[672] * mat_B[15] +
//             mat_A[673] * mat_B[47] +
//             mat_A[674] * mat_B[79] +
//             mat_A[675] * mat_B[111] +
//             mat_A[676] * mat_B[143] +
//             mat_A[677] * mat_B[175] +
//             mat_A[678] * mat_B[207] +
//             mat_A[679] * mat_B[239] +
//             mat_A[680] * mat_B[271] +
//             mat_A[681] * mat_B[303] +
//             mat_A[682] * mat_B[335] +
//             mat_A[683] * mat_B[367] +
//             mat_A[684] * mat_B[399] +
//             mat_A[685] * mat_B[431] +
//             mat_A[686] * mat_B[463] +
//             mat_A[687] * mat_B[495] +
//             mat_A[688] * mat_B[527] +
//             mat_A[689] * mat_B[559] +
//             mat_A[690] * mat_B[591] +
//             mat_A[691] * mat_B[623] +
//             mat_A[692] * mat_B[655] +
//             mat_A[693] * mat_B[687] +
//             mat_A[694] * mat_B[719] +
//             mat_A[695] * mat_B[751] +
//             mat_A[696] * mat_B[783] +
//             mat_A[697] * mat_B[815] +
//             mat_A[698] * mat_B[847] +
//             mat_A[699] * mat_B[879] +
//             mat_A[700] * mat_B[911] +
//             mat_A[701] * mat_B[943] +
//             mat_A[702] * mat_B[975] +
//             mat_A[703] * mat_B[1007];
//  mat_C[688] <= 
//             mat_A[672] * mat_B[16] +
//             mat_A[673] * mat_B[48] +
//             mat_A[674] * mat_B[80] +
//             mat_A[675] * mat_B[112] +
//             mat_A[676] * mat_B[144] +
//             mat_A[677] * mat_B[176] +
//             mat_A[678] * mat_B[208] +
//             mat_A[679] * mat_B[240] +
//             mat_A[680] * mat_B[272] +
//             mat_A[681] * mat_B[304] +
//             mat_A[682] * mat_B[336] +
//             mat_A[683] * mat_B[368] +
//             mat_A[684] * mat_B[400] +
//             mat_A[685] * mat_B[432] +
//             mat_A[686] * mat_B[464] +
//             mat_A[687] * mat_B[496] +
//             mat_A[688] * mat_B[528] +
//             mat_A[689] * mat_B[560] +
//             mat_A[690] * mat_B[592] +
//             mat_A[691] * mat_B[624] +
//             mat_A[692] * mat_B[656] +
//             mat_A[693] * mat_B[688] +
//             mat_A[694] * mat_B[720] +
//             mat_A[695] * mat_B[752] +
//             mat_A[696] * mat_B[784] +
//             mat_A[697] * mat_B[816] +
//             mat_A[698] * mat_B[848] +
//             mat_A[699] * mat_B[880] +
//             mat_A[700] * mat_B[912] +
//             mat_A[701] * mat_B[944] +
//             mat_A[702] * mat_B[976] +
//             mat_A[703] * mat_B[1008];
//  mat_C[689] <= 
//             mat_A[672] * mat_B[17] +
//             mat_A[673] * mat_B[49] +
//             mat_A[674] * mat_B[81] +
//             mat_A[675] * mat_B[113] +
//             mat_A[676] * mat_B[145] +
//             mat_A[677] * mat_B[177] +
//             mat_A[678] * mat_B[209] +
//             mat_A[679] * mat_B[241] +
//             mat_A[680] * mat_B[273] +
//             mat_A[681] * mat_B[305] +
//             mat_A[682] * mat_B[337] +
//             mat_A[683] * mat_B[369] +
//             mat_A[684] * mat_B[401] +
//             mat_A[685] * mat_B[433] +
//             mat_A[686] * mat_B[465] +
//             mat_A[687] * mat_B[497] +
//             mat_A[688] * mat_B[529] +
//             mat_A[689] * mat_B[561] +
//             mat_A[690] * mat_B[593] +
//             mat_A[691] * mat_B[625] +
//             mat_A[692] * mat_B[657] +
//             mat_A[693] * mat_B[689] +
//             mat_A[694] * mat_B[721] +
//             mat_A[695] * mat_B[753] +
//             mat_A[696] * mat_B[785] +
//             mat_A[697] * mat_B[817] +
//             mat_A[698] * mat_B[849] +
//             mat_A[699] * mat_B[881] +
//             mat_A[700] * mat_B[913] +
//             mat_A[701] * mat_B[945] +
//             mat_A[702] * mat_B[977] +
//             mat_A[703] * mat_B[1009];
//  mat_C[690] <= 
//             mat_A[672] * mat_B[18] +
//             mat_A[673] * mat_B[50] +
//             mat_A[674] * mat_B[82] +
//             mat_A[675] * mat_B[114] +
//             mat_A[676] * mat_B[146] +
//             mat_A[677] * mat_B[178] +
//             mat_A[678] * mat_B[210] +
//             mat_A[679] * mat_B[242] +
//             mat_A[680] * mat_B[274] +
//             mat_A[681] * mat_B[306] +
//             mat_A[682] * mat_B[338] +
//             mat_A[683] * mat_B[370] +
//             mat_A[684] * mat_B[402] +
//             mat_A[685] * mat_B[434] +
//             mat_A[686] * mat_B[466] +
//             mat_A[687] * mat_B[498] +
//             mat_A[688] * mat_B[530] +
//             mat_A[689] * mat_B[562] +
//             mat_A[690] * mat_B[594] +
//             mat_A[691] * mat_B[626] +
//             mat_A[692] * mat_B[658] +
//             mat_A[693] * mat_B[690] +
//             mat_A[694] * mat_B[722] +
//             mat_A[695] * mat_B[754] +
//             mat_A[696] * mat_B[786] +
//             mat_A[697] * mat_B[818] +
//             mat_A[698] * mat_B[850] +
//             mat_A[699] * mat_B[882] +
//             mat_A[700] * mat_B[914] +
//             mat_A[701] * mat_B[946] +
//             mat_A[702] * mat_B[978] +
//             mat_A[703] * mat_B[1010];
//  mat_C[691] <= 
//             mat_A[672] * mat_B[19] +
//             mat_A[673] * mat_B[51] +
//             mat_A[674] * mat_B[83] +
//             mat_A[675] * mat_B[115] +
//             mat_A[676] * mat_B[147] +
//             mat_A[677] * mat_B[179] +
//             mat_A[678] * mat_B[211] +
//             mat_A[679] * mat_B[243] +
//             mat_A[680] * mat_B[275] +
//             mat_A[681] * mat_B[307] +
//             mat_A[682] * mat_B[339] +
//             mat_A[683] * mat_B[371] +
//             mat_A[684] * mat_B[403] +
//             mat_A[685] * mat_B[435] +
//             mat_A[686] * mat_B[467] +
//             mat_A[687] * mat_B[499] +
//             mat_A[688] * mat_B[531] +
//             mat_A[689] * mat_B[563] +
//             mat_A[690] * mat_B[595] +
//             mat_A[691] * mat_B[627] +
//             mat_A[692] * mat_B[659] +
//             mat_A[693] * mat_B[691] +
//             mat_A[694] * mat_B[723] +
//             mat_A[695] * mat_B[755] +
//             mat_A[696] * mat_B[787] +
//             mat_A[697] * mat_B[819] +
//             mat_A[698] * mat_B[851] +
//             mat_A[699] * mat_B[883] +
//             mat_A[700] * mat_B[915] +
//             mat_A[701] * mat_B[947] +
//             mat_A[702] * mat_B[979] +
//             mat_A[703] * mat_B[1011];
//  mat_C[692] <= 
//             mat_A[672] * mat_B[20] +
//             mat_A[673] * mat_B[52] +
//             mat_A[674] * mat_B[84] +
//             mat_A[675] * mat_B[116] +
//             mat_A[676] * mat_B[148] +
//             mat_A[677] * mat_B[180] +
//             mat_A[678] * mat_B[212] +
//             mat_A[679] * mat_B[244] +
//             mat_A[680] * mat_B[276] +
//             mat_A[681] * mat_B[308] +
//             mat_A[682] * mat_B[340] +
//             mat_A[683] * mat_B[372] +
//             mat_A[684] * mat_B[404] +
//             mat_A[685] * mat_B[436] +
//             mat_A[686] * mat_B[468] +
//             mat_A[687] * mat_B[500] +
//             mat_A[688] * mat_B[532] +
//             mat_A[689] * mat_B[564] +
//             mat_A[690] * mat_B[596] +
//             mat_A[691] * mat_B[628] +
//             mat_A[692] * mat_B[660] +
//             mat_A[693] * mat_B[692] +
//             mat_A[694] * mat_B[724] +
//             mat_A[695] * mat_B[756] +
//             mat_A[696] * mat_B[788] +
//             mat_A[697] * mat_B[820] +
//             mat_A[698] * mat_B[852] +
//             mat_A[699] * mat_B[884] +
//             mat_A[700] * mat_B[916] +
//             mat_A[701] * mat_B[948] +
//             mat_A[702] * mat_B[980] +
//             mat_A[703] * mat_B[1012];
//  mat_C[693] <= 
//             mat_A[672] * mat_B[21] +
//             mat_A[673] * mat_B[53] +
//             mat_A[674] * mat_B[85] +
//             mat_A[675] * mat_B[117] +
//             mat_A[676] * mat_B[149] +
//             mat_A[677] * mat_B[181] +
//             mat_A[678] * mat_B[213] +
//             mat_A[679] * mat_B[245] +
//             mat_A[680] * mat_B[277] +
//             mat_A[681] * mat_B[309] +
//             mat_A[682] * mat_B[341] +
//             mat_A[683] * mat_B[373] +
//             mat_A[684] * mat_B[405] +
//             mat_A[685] * mat_B[437] +
//             mat_A[686] * mat_B[469] +
//             mat_A[687] * mat_B[501] +
//             mat_A[688] * mat_B[533] +
//             mat_A[689] * mat_B[565] +
//             mat_A[690] * mat_B[597] +
//             mat_A[691] * mat_B[629] +
//             mat_A[692] * mat_B[661] +
//             mat_A[693] * mat_B[693] +
//             mat_A[694] * mat_B[725] +
//             mat_A[695] * mat_B[757] +
//             mat_A[696] * mat_B[789] +
//             mat_A[697] * mat_B[821] +
//             mat_A[698] * mat_B[853] +
//             mat_A[699] * mat_B[885] +
//             mat_A[700] * mat_B[917] +
//             mat_A[701] * mat_B[949] +
//             mat_A[702] * mat_B[981] +
//             mat_A[703] * mat_B[1013];
//  mat_C[694] <= 
//             mat_A[672] * mat_B[22] +
//             mat_A[673] * mat_B[54] +
//             mat_A[674] * mat_B[86] +
//             mat_A[675] * mat_B[118] +
//             mat_A[676] * mat_B[150] +
//             mat_A[677] * mat_B[182] +
//             mat_A[678] * mat_B[214] +
//             mat_A[679] * mat_B[246] +
//             mat_A[680] * mat_B[278] +
//             mat_A[681] * mat_B[310] +
//             mat_A[682] * mat_B[342] +
//             mat_A[683] * mat_B[374] +
//             mat_A[684] * mat_B[406] +
//             mat_A[685] * mat_B[438] +
//             mat_A[686] * mat_B[470] +
//             mat_A[687] * mat_B[502] +
//             mat_A[688] * mat_B[534] +
//             mat_A[689] * mat_B[566] +
//             mat_A[690] * mat_B[598] +
//             mat_A[691] * mat_B[630] +
//             mat_A[692] * mat_B[662] +
//             mat_A[693] * mat_B[694] +
//             mat_A[694] * mat_B[726] +
//             mat_A[695] * mat_B[758] +
//             mat_A[696] * mat_B[790] +
//             mat_A[697] * mat_B[822] +
//             mat_A[698] * mat_B[854] +
//             mat_A[699] * mat_B[886] +
//             mat_A[700] * mat_B[918] +
//             mat_A[701] * mat_B[950] +
//             mat_A[702] * mat_B[982] +
//             mat_A[703] * mat_B[1014];
//  mat_C[695] <= 
//             mat_A[672] * mat_B[23] +
//             mat_A[673] * mat_B[55] +
//             mat_A[674] * mat_B[87] +
//             mat_A[675] * mat_B[119] +
//             mat_A[676] * mat_B[151] +
//             mat_A[677] * mat_B[183] +
//             mat_A[678] * mat_B[215] +
//             mat_A[679] * mat_B[247] +
//             mat_A[680] * mat_B[279] +
//             mat_A[681] * mat_B[311] +
//             mat_A[682] * mat_B[343] +
//             mat_A[683] * mat_B[375] +
//             mat_A[684] * mat_B[407] +
//             mat_A[685] * mat_B[439] +
//             mat_A[686] * mat_B[471] +
//             mat_A[687] * mat_B[503] +
//             mat_A[688] * mat_B[535] +
//             mat_A[689] * mat_B[567] +
//             mat_A[690] * mat_B[599] +
//             mat_A[691] * mat_B[631] +
//             mat_A[692] * mat_B[663] +
//             mat_A[693] * mat_B[695] +
//             mat_A[694] * mat_B[727] +
//             mat_A[695] * mat_B[759] +
//             mat_A[696] * mat_B[791] +
//             mat_A[697] * mat_B[823] +
//             mat_A[698] * mat_B[855] +
//             mat_A[699] * mat_B[887] +
//             mat_A[700] * mat_B[919] +
//             mat_A[701] * mat_B[951] +
//             mat_A[702] * mat_B[983] +
//             mat_A[703] * mat_B[1015];
//  mat_C[696] <= 
//             mat_A[672] * mat_B[24] +
//             mat_A[673] * mat_B[56] +
//             mat_A[674] * mat_B[88] +
//             mat_A[675] * mat_B[120] +
//             mat_A[676] * mat_B[152] +
//             mat_A[677] * mat_B[184] +
//             mat_A[678] * mat_B[216] +
//             mat_A[679] * mat_B[248] +
//             mat_A[680] * mat_B[280] +
//             mat_A[681] * mat_B[312] +
//             mat_A[682] * mat_B[344] +
//             mat_A[683] * mat_B[376] +
//             mat_A[684] * mat_B[408] +
//             mat_A[685] * mat_B[440] +
//             mat_A[686] * mat_B[472] +
//             mat_A[687] * mat_B[504] +
//             mat_A[688] * mat_B[536] +
//             mat_A[689] * mat_B[568] +
//             mat_A[690] * mat_B[600] +
//             mat_A[691] * mat_B[632] +
//             mat_A[692] * mat_B[664] +
//             mat_A[693] * mat_B[696] +
//             mat_A[694] * mat_B[728] +
//             mat_A[695] * mat_B[760] +
//             mat_A[696] * mat_B[792] +
//             mat_A[697] * mat_B[824] +
//             mat_A[698] * mat_B[856] +
//             mat_A[699] * mat_B[888] +
//             mat_A[700] * mat_B[920] +
//             mat_A[701] * mat_B[952] +
//             mat_A[702] * mat_B[984] +
//             mat_A[703] * mat_B[1016];
//  mat_C[697] <= 
//             mat_A[672] * mat_B[25] +
//             mat_A[673] * mat_B[57] +
//             mat_A[674] * mat_B[89] +
//             mat_A[675] * mat_B[121] +
//             mat_A[676] * mat_B[153] +
//             mat_A[677] * mat_B[185] +
//             mat_A[678] * mat_B[217] +
//             mat_A[679] * mat_B[249] +
//             mat_A[680] * mat_B[281] +
//             mat_A[681] * mat_B[313] +
//             mat_A[682] * mat_B[345] +
//             mat_A[683] * mat_B[377] +
//             mat_A[684] * mat_B[409] +
//             mat_A[685] * mat_B[441] +
//             mat_A[686] * mat_B[473] +
//             mat_A[687] * mat_B[505] +
//             mat_A[688] * mat_B[537] +
//             mat_A[689] * mat_B[569] +
//             mat_A[690] * mat_B[601] +
//             mat_A[691] * mat_B[633] +
//             mat_A[692] * mat_B[665] +
//             mat_A[693] * mat_B[697] +
//             mat_A[694] * mat_B[729] +
//             mat_A[695] * mat_B[761] +
//             mat_A[696] * mat_B[793] +
//             mat_A[697] * mat_B[825] +
//             mat_A[698] * mat_B[857] +
//             mat_A[699] * mat_B[889] +
//             mat_A[700] * mat_B[921] +
//             mat_A[701] * mat_B[953] +
//             mat_A[702] * mat_B[985] +
//             mat_A[703] * mat_B[1017];
//  mat_C[698] <= 
//             mat_A[672] * mat_B[26] +
//             mat_A[673] * mat_B[58] +
//             mat_A[674] * mat_B[90] +
//             mat_A[675] * mat_B[122] +
//             mat_A[676] * mat_B[154] +
//             mat_A[677] * mat_B[186] +
//             mat_A[678] * mat_B[218] +
//             mat_A[679] * mat_B[250] +
//             mat_A[680] * mat_B[282] +
//             mat_A[681] * mat_B[314] +
//             mat_A[682] * mat_B[346] +
//             mat_A[683] * mat_B[378] +
//             mat_A[684] * mat_B[410] +
//             mat_A[685] * mat_B[442] +
//             mat_A[686] * mat_B[474] +
//             mat_A[687] * mat_B[506] +
//             mat_A[688] * mat_B[538] +
//             mat_A[689] * mat_B[570] +
//             mat_A[690] * mat_B[602] +
//             mat_A[691] * mat_B[634] +
//             mat_A[692] * mat_B[666] +
//             mat_A[693] * mat_B[698] +
//             mat_A[694] * mat_B[730] +
//             mat_A[695] * mat_B[762] +
//             mat_A[696] * mat_B[794] +
//             mat_A[697] * mat_B[826] +
//             mat_A[698] * mat_B[858] +
//             mat_A[699] * mat_B[890] +
//             mat_A[700] * mat_B[922] +
//             mat_A[701] * mat_B[954] +
//             mat_A[702] * mat_B[986] +
//             mat_A[703] * mat_B[1018];
//  mat_C[699] <= 
//             mat_A[672] * mat_B[27] +
//             mat_A[673] * mat_B[59] +
//             mat_A[674] * mat_B[91] +
//             mat_A[675] * mat_B[123] +
//             mat_A[676] * mat_B[155] +
//             mat_A[677] * mat_B[187] +
//             mat_A[678] * mat_B[219] +
//             mat_A[679] * mat_B[251] +
//             mat_A[680] * mat_B[283] +
//             mat_A[681] * mat_B[315] +
//             mat_A[682] * mat_B[347] +
//             mat_A[683] * mat_B[379] +
//             mat_A[684] * mat_B[411] +
//             mat_A[685] * mat_B[443] +
//             mat_A[686] * mat_B[475] +
//             mat_A[687] * mat_B[507] +
//             mat_A[688] * mat_B[539] +
//             mat_A[689] * mat_B[571] +
//             mat_A[690] * mat_B[603] +
//             mat_A[691] * mat_B[635] +
//             mat_A[692] * mat_B[667] +
//             mat_A[693] * mat_B[699] +
//             mat_A[694] * mat_B[731] +
//             mat_A[695] * mat_B[763] +
//             mat_A[696] * mat_B[795] +
//             mat_A[697] * mat_B[827] +
//             mat_A[698] * mat_B[859] +
//             mat_A[699] * mat_B[891] +
//             mat_A[700] * mat_B[923] +
//             mat_A[701] * mat_B[955] +
//             mat_A[702] * mat_B[987] +
//             mat_A[703] * mat_B[1019];
//  mat_C[700] <= 
//             mat_A[672] * mat_B[28] +
//             mat_A[673] * mat_B[60] +
//             mat_A[674] * mat_B[92] +
//             mat_A[675] * mat_B[124] +
//             mat_A[676] * mat_B[156] +
//             mat_A[677] * mat_B[188] +
//             mat_A[678] * mat_B[220] +
//             mat_A[679] * mat_B[252] +
//             mat_A[680] * mat_B[284] +
//             mat_A[681] * mat_B[316] +
//             mat_A[682] * mat_B[348] +
//             mat_A[683] * mat_B[380] +
//             mat_A[684] * mat_B[412] +
//             mat_A[685] * mat_B[444] +
//             mat_A[686] * mat_B[476] +
//             mat_A[687] * mat_B[508] +
//             mat_A[688] * mat_B[540] +
//             mat_A[689] * mat_B[572] +
//             mat_A[690] * mat_B[604] +
//             mat_A[691] * mat_B[636] +
//             mat_A[692] * mat_B[668] +
//             mat_A[693] * mat_B[700] +
//             mat_A[694] * mat_B[732] +
//             mat_A[695] * mat_B[764] +
//             mat_A[696] * mat_B[796] +
//             mat_A[697] * mat_B[828] +
//             mat_A[698] * mat_B[860] +
//             mat_A[699] * mat_B[892] +
//             mat_A[700] * mat_B[924] +
//             mat_A[701] * mat_B[956] +
//             mat_A[702] * mat_B[988] +
//             mat_A[703] * mat_B[1020];
//  mat_C[701] <= 
//             mat_A[672] * mat_B[29] +
//             mat_A[673] * mat_B[61] +
//             mat_A[674] * mat_B[93] +
//             mat_A[675] * mat_B[125] +
//             mat_A[676] * mat_B[157] +
//             mat_A[677] * mat_B[189] +
//             mat_A[678] * mat_B[221] +
//             mat_A[679] * mat_B[253] +
//             mat_A[680] * mat_B[285] +
//             mat_A[681] * mat_B[317] +
//             mat_A[682] * mat_B[349] +
//             mat_A[683] * mat_B[381] +
//             mat_A[684] * mat_B[413] +
//             mat_A[685] * mat_B[445] +
//             mat_A[686] * mat_B[477] +
//             mat_A[687] * mat_B[509] +
//             mat_A[688] * mat_B[541] +
//             mat_A[689] * mat_B[573] +
//             mat_A[690] * mat_B[605] +
//             mat_A[691] * mat_B[637] +
//             mat_A[692] * mat_B[669] +
//             mat_A[693] * mat_B[701] +
//             mat_A[694] * mat_B[733] +
//             mat_A[695] * mat_B[765] +
//             mat_A[696] * mat_B[797] +
//             mat_A[697] * mat_B[829] +
//             mat_A[698] * mat_B[861] +
//             mat_A[699] * mat_B[893] +
//             mat_A[700] * mat_B[925] +
//             mat_A[701] * mat_B[957] +
//             mat_A[702] * mat_B[989] +
//             mat_A[703] * mat_B[1021];
//  mat_C[702] <= 
//             mat_A[672] * mat_B[30] +
//             mat_A[673] * mat_B[62] +
//             mat_A[674] * mat_B[94] +
//             mat_A[675] * mat_B[126] +
//             mat_A[676] * mat_B[158] +
//             mat_A[677] * mat_B[190] +
//             mat_A[678] * mat_B[222] +
//             mat_A[679] * mat_B[254] +
//             mat_A[680] * mat_B[286] +
//             mat_A[681] * mat_B[318] +
//             mat_A[682] * mat_B[350] +
//             mat_A[683] * mat_B[382] +
//             mat_A[684] * mat_B[414] +
//             mat_A[685] * mat_B[446] +
//             mat_A[686] * mat_B[478] +
//             mat_A[687] * mat_B[510] +
//             mat_A[688] * mat_B[542] +
//             mat_A[689] * mat_B[574] +
//             mat_A[690] * mat_B[606] +
//             mat_A[691] * mat_B[638] +
//             mat_A[692] * mat_B[670] +
//             mat_A[693] * mat_B[702] +
//             mat_A[694] * mat_B[734] +
//             mat_A[695] * mat_B[766] +
//             mat_A[696] * mat_B[798] +
//             mat_A[697] * mat_B[830] +
//             mat_A[698] * mat_B[862] +
//             mat_A[699] * mat_B[894] +
//             mat_A[700] * mat_B[926] +
//             mat_A[701] * mat_B[958] +
//             mat_A[702] * mat_B[990] +
//             mat_A[703] * mat_B[1022];
//  mat_C[703] <= 
//             mat_A[672] * mat_B[31] +
//             mat_A[673] * mat_B[63] +
//             mat_A[674] * mat_B[95] +
//             mat_A[675] * mat_B[127] +
//             mat_A[676] * mat_B[159] +
//             mat_A[677] * mat_B[191] +
//             mat_A[678] * mat_B[223] +
//             mat_A[679] * mat_B[255] +
//             mat_A[680] * mat_B[287] +
//             mat_A[681] * mat_B[319] +
//             mat_A[682] * mat_B[351] +
//             mat_A[683] * mat_B[383] +
//             mat_A[684] * mat_B[415] +
//             mat_A[685] * mat_B[447] +
//             mat_A[686] * mat_B[479] +
//             mat_A[687] * mat_B[511] +
//             mat_A[688] * mat_B[543] +
//             mat_A[689] * mat_B[575] +
//             mat_A[690] * mat_B[607] +
//             mat_A[691] * mat_B[639] +
//             mat_A[692] * mat_B[671] +
//             mat_A[693] * mat_B[703] +
//             mat_A[694] * mat_B[735] +
//             mat_A[695] * mat_B[767] +
//             mat_A[696] * mat_B[799] +
//             mat_A[697] * mat_B[831] +
//             mat_A[698] * mat_B[863] +
//             mat_A[699] * mat_B[895] +
//             mat_A[700] * mat_B[927] +
//             mat_A[701] * mat_B[959] +
//             mat_A[702] * mat_B[991] +
//             mat_A[703] * mat_B[1023];
//  mat_C[704] <= 
//             mat_A[704] * mat_B[0] +
//             mat_A[705] * mat_B[32] +
//             mat_A[706] * mat_B[64] +
//             mat_A[707] * mat_B[96] +
//             mat_A[708] * mat_B[128] +
//             mat_A[709] * mat_B[160] +
//             mat_A[710] * mat_B[192] +
//             mat_A[711] * mat_B[224] +
//             mat_A[712] * mat_B[256] +
//             mat_A[713] * mat_B[288] +
//             mat_A[714] * mat_B[320] +
//             mat_A[715] * mat_B[352] +
//             mat_A[716] * mat_B[384] +
//             mat_A[717] * mat_B[416] +
//             mat_A[718] * mat_B[448] +
//             mat_A[719] * mat_B[480] +
//             mat_A[720] * mat_B[512] +
//             mat_A[721] * mat_B[544] +
//             mat_A[722] * mat_B[576] +
//             mat_A[723] * mat_B[608] +
//             mat_A[724] * mat_B[640] +
//             mat_A[725] * mat_B[672] +
//             mat_A[726] * mat_B[704] +
//             mat_A[727] * mat_B[736] +
//             mat_A[728] * mat_B[768] +
//             mat_A[729] * mat_B[800] +
//             mat_A[730] * mat_B[832] +
//             mat_A[731] * mat_B[864] +
//             mat_A[732] * mat_B[896] +
//             mat_A[733] * mat_B[928] +
//             mat_A[734] * mat_B[960] +
//             mat_A[735] * mat_B[992];
//  mat_C[705] <= 
//             mat_A[704] * mat_B[1] +
//             mat_A[705] * mat_B[33] +
//             mat_A[706] * mat_B[65] +
//             mat_A[707] * mat_B[97] +
//             mat_A[708] * mat_B[129] +
//             mat_A[709] * mat_B[161] +
//             mat_A[710] * mat_B[193] +
//             mat_A[711] * mat_B[225] +
//             mat_A[712] * mat_B[257] +
//             mat_A[713] * mat_B[289] +
//             mat_A[714] * mat_B[321] +
//             mat_A[715] * mat_B[353] +
//             mat_A[716] * mat_B[385] +
//             mat_A[717] * mat_B[417] +
//             mat_A[718] * mat_B[449] +
//             mat_A[719] * mat_B[481] +
//             mat_A[720] * mat_B[513] +
//             mat_A[721] * mat_B[545] +
//             mat_A[722] * mat_B[577] +
//             mat_A[723] * mat_B[609] +
//             mat_A[724] * mat_B[641] +
//             mat_A[725] * mat_B[673] +
//             mat_A[726] * mat_B[705] +
//             mat_A[727] * mat_B[737] +
//             mat_A[728] * mat_B[769] +
//             mat_A[729] * mat_B[801] +
//             mat_A[730] * mat_B[833] +
//             mat_A[731] * mat_B[865] +
//             mat_A[732] * mat_B[897] +
//             mat_A[733] * mat_B[929] +
//             mat_A[734] * mat_B[961] +
//             mat_A[735] * mat_B[993];
//  mat_C[706] <= 
//             mat_A[704] * mat_B[2] +
//             mat_A[705] * mat_B[34] +
//             mat_A[706] * mat_B[66] +
//             mat_A[707] * mat_B[98] +
//             mat_A[708] * mat_B[130] +
//             mat_A[709] * mat_B[162] +
//             mat_A[710] * mat_B[194] +
//             mat_A[711] * mat_B[226] +
//             mat_A[712] * mat_B[258] +
//             mat_A[713] * mat_B[290] +
//             mat_A[714] * mat_B[322] +
//             mat_A[715] * mat_B[354] +
//             mat_A[716] * mat_B[386] +
//             mat_A[717] * mat_B[418] +
//             mat_A[718] * mat_B[450] +
//             mat_A[719] * mat_B[482] +
//             mat_A[720] * mat_B[514] +
//             mat_A[721] * mat_B[546] +
//             mat_A[722] * mat_B[578] +
//             mat_A[723] * mat_B[610] +
//             mat_A[724] * mat_B[642] +
//             mat_A[725] * mat_B[674] +
//             mat_A[726] * mat_B[706] +
//             mat_A[727] * mat_B[738] +
//             mat_A[728] * mat_B[770] +
//             mat_A[729] * mat_B[802] +
//             mat_A[730] * mat_B[834] +
//             mat_A[731] * mat_B[866] +
//             mat_A[732] * mat_B[898] +
//             mat_A[733] * mat_B[930] +
//             mat_A[734] * mat_B[962] +
//             mat_A[735] * mat_B[994];
//  mat_C[707] <= 
//             mat_A[704] * mat_B[3] +
//             mat_A[705] * mat_B[35] +
//             mat_A[706] * mat_B[67] +
//             mat_A[707] * mat_B[99] +
//             mat_A[708] * mat_B[131] +
//             mat_A[709] * mat_B[163] +
//             mat_A[710] * mat_B[195] +
//             mat_A[711] * mat_B[227] +
//             mat_A[712] * mat_B[259] +
//             mat_A[713] * mat_B[291] +
//             mat_A[714] * mat_B[323] +
//             mat_A[715] * mat_B[355] +
//             mat_A[716] * mat_B[387] +
//             mat_A[717] * mat_B[419] +
//             mat_A[718] * mat_B[451] +
//             mat_A[719] * mat_B[483] +
//             mat_A[720] * mat_B[515] +
//             mat_A[721] * mat_B[547] +
//             mat_A[722] * mat_B[579] +
//             mat_A[723] * mat_B[611] +
//             mat_A[724] * mat_B[643] +
//             mat_A[725] * mat_B[675] +
//             mat_A[726] * mat_B[707] +
//             mat_A[727] * mat_B[739] +
//             mat_A[728] * mat_B[771] +
//             mat_A[729] * mat_B[803] +
//             mat_A[730] * mat_B[835] +
//             mat_A[731] * mat_B[867] +
//             mat_A[732] * mat_B[899] +
//             mat_A[733] * mat_B[931] +
//             mat_A[734] * mat_B[963] +
//             mat_A[735] * mat_B[995];
//  mat_C[708] <= 
//             mat_A[704] * mat_B[4] +
//             mat_A[705] * mat_B[36] +
//             mat_A[706] * mat_B[68] +
//             mat_A[707] * mat_B[100] +
//             mat_A[708] * mat_B[132] +
//             mat_A[709] * mat_B[164] +
//             mat_A[710] * mat_B[196] +
//             mat_A[711] * mat_B[228] +
//             mat_A[712] * mat_B[260] +
//             mat_A[713] * mat_B[292] +
//             mat_A[714] * mat_B[324] +
//             mat_A[715] * mat_B[356] +
//             mat_A[716] * mat_B[388] +
//             mat_A[717] * mat_B[420] +
//             mat_A[718] * mat_B[452] +
//             mat_A[719] * mat_B[484] +
//             mat_A[720] * mat_B[516] +
//             mat_A[721] * mat_B[548] +
//             mat_A[722] * mat_B[580] +
//             mat_A[723] * mat_B[612] +
//             mat_A[724] * mat_B[644] +
//             mat_A[725] * mat_B[676] +
//             mat_A[726] * mat_B[708] +
//             mat_A[727] * mat_B[740] +
//             mat_A[728] * mat_B[772] +
//             mat_A[729] * mat_B[804] +
//             mat_A[730] * mat_B[836] +
//             mat_A[731] * mat_B[868] +
//             mat_A[732] * mat_B[900] +
//             mat_A[733] * mat_B[932] +
//             mat_A[734] * mat_B[964] +
//             mat_A[735] * mat_B[996];
//  mat_C[709] <= 
//             mat_A[704] * mat_B[5] +
//             mat_A[705] * mat_B[37] +
//             mat_A[706] * mat_B[69] +
//             mat_A[707] * mat_B[101] +
//             mat_A[708] * mat_B[133] +
//             mat_A[709] * mat_B[165] +
//             mat_A[710] * mat_B[197] +
//             mat_A[711] * mat_B[229] +
//             mat_A[712] * mat_B[261] +
//             mat_A[713] * mat_B[293] +
//             mat_A[714] * mat_B[325] +
//             mat_A[715] * mat_B[357] +
//             mat_A[716] * mat_B[389] +
//             mat_A[717] * mat_B[421] +
//             mat_A[718] * mat_B[453] +
//             mat_A[719] * mat_B[485] +
//             mat_A[720] * mat_B[517] +
//             mat_A[721] * mat_B[549] +
//             mat_A[722] * mat_B[581] +
//             mat_A[723] * mat_B[613] +
//             mat_A[724] * mat_B[645] +
//             mat_A[725] * mat_B[677] +
//             mat_A[726] * mat_B[709] +
//             mat_A[727] * mat_B[741] +
//             mat_A[728] * mat_B[773] +
//             mat_A[729] * mat_B[805] +
//             mat_A[730] * mat_B[837] +
//             mat_A[731] * mat_B[869] +
//             mat_A[732] * mat_B[901] +
//             mat_A[733] * mat_B[933] +
//             mat_A[734] * mat_B[965] +
//             mat_A[735] * mat_B[997];
//  mat_C[710] <= 
//             mat_A[704] * mat_B[6] +
//             mat_A[705] * mat_B[38] +
//             mat_A[706] * mat_B[70] +
//             mat_A[707] * mat_B[102] +
//             mat_A[708] * mat_B[134] +
//             mat_A[709] * mat_B[166] +
//             mat_A[710] * mat_B[198] +
//             mat_A[711] * mat_B[230] +
//             mat_A[712] * mat_B[262] +
//             mat_A[713] * mat_B[294] +
//             mat_A[714] * mat_B[326] +
//             mat_A[715] * mat_B[358] +
//             mat_A[716] * mat_B[390] +
//             mat_A[717] * mat_B[422] +
//             mat_A[718] * mat_B[454] +
//             mat_A[719] * mat_B[486] +
//             mat_A[720] * mat_B[518] +
//             mat_A[721] * mat_B[550] +
//             mat_A[722] * mat_B[582] +
//             mat_A[723] * mat_B[614] +
//             mat_A[724] * mat_B[646] +
//             mat_A[725] * mat_B[678] +
//             mat_A[726] * mat_B[710] +
//             mat_A[727] * mat_B[742] +
//             mat_A[728] * mat_B[774] +
//             mat_A[729] * mat_B[806] +
//             mat_A[730] * mat_B[838] +
//             mat_A[731] * mat_B[870] +
//             mat_A[732] * mat_B[902] +
//             mat_A[733] * mat_B[934] +
//             mat_A[734] * mat_B[966] +
//             mat_A[735] * mat_B[998];
//  mat_C[711] <= 
//             mat_A[704] * mat_B[7] +
//             mat_A[705] * mat_B[39] +
//             mat_A[706] * mat_B[71] +
//             mat_A[707] * mat_B[103] +
//             mat_A[708] * mat_B[135] +
//             mat_A[709] * mat_B[167] +
//             mat_A[710] * mat_B[199] +
//             mat_A[711] * mat_B[231] +
//             mat_A[712] * mat_B[263] +
//             mat_A[713] * mat_B[295] +
//             mat_A[714] * mat_B[327] +
//             mat_A[715] * mat_B[359] +
//             mat_A[716] * mat_B[391] +
//             mat_A[717] * mat_B[423] +
//             mat_A[718] * mat_B[455] +
//             mat_A[719] * mat_B[487] +
//             mat_A[720] * mat_B[519] +
//             mat_A[721] * mat_B[551] +
//             mat_A[722] * mat_B[583] +
//             mat_A[723] * mat_B[615] +
//             mat_A[724] * mat_B[647] +
//             mat_A[725] * mat_B[679] +
//             mat_A[726] * mat_B[711] +
//             mat_A[727] * mat_B[743] +
//             mat_A[728] * mat_B[775] +
//             mat_A[729] * mat_B[807] +
//             mat_A[730] * mat_B[839] +
//             mat_A[731] * mat_B[871] +
//             mat_A[732] * mat_B[903] +
//             mat_A[733] * mat_B[935] +
//             mat_A[734] * mat_B[967] +
//             mat_A[735] * mat_B[999];
//  mat_C[712] <= 
//             mat_A[704] * mat_B[8] +
//             mat_A[705] * mat_B[40] +
//             mat_A[706] * mat_B[72] +
//             mat_A[707] * mat_B[104] +
//             mat_A[708] * mat_B[136] +
//             mat_A[709] * mat_B[168] +
//             mat_A[710] * mat_B[200] +
//             mat_A[711] * mat_B[232] +
//             mat_A[712] * mat_B[264] +
//             mat_A[713] * mat_B[296] +
//             mat_A[714] * mat_B[328] +
//             mat_A[715] * mat_B[360] +
//             mat_A[716] * mat_B[392] +
//             mat_A[717] * mat_B[424] +
//             mat_A[718] * mat_B[456] +
//             mat_A[719] * mat_B[488] +
//             mat_A[720] * mat_B[520] +
//             mat_A[721] * mat_B[552] +
//             mat_A[722] * mat_B[584] +
//             mat_A[723] * mat_B[616] +
//             mat_A[724] * mat_B[648] +
//             mat_A[725] * mat_B[680] +
//             mat_A[726] * mat_B[712] +
//             mat_A[727] * mat_B[744] +
//             mat_A[728] * mat_B[776] +
//             mat_A[729] * mat_B[808] +
//             mat_A[730] * mat_B[840] +
//             mat_A[731] * mat_B[872] +
//             mat_A[732] * mat_B[904] +
//             mat_A[733] * mat_B[936] +
//             mat_A[734] * mat_B[968] +
//             mat_A[735] * mat_B[1000];
//  mat_C[713] <= 
//             mat_A[704] * mat_B[9] +
//             mat_A[705] * mat_B[41] +
//             mat_A[706] * mat_B[73] +
//             mat_A[707] * mat_B[105] +
//             mat_A[708] * mat_B[137] +
//             mat_A[709] * mat_B[169] +
//             mat_A[710] * mat_B[201] +
//             mat_A[711] * mat_B[233] +
//             mat_A[712] * mat_B[265] +
//             mat_A[713] * mat_B[297] +
//             mat_A[714] * mat_B[329] +
//             mat_A[715] * mat_B[361] +
//             mat_A[716] * mat_B[393] +
//             mat_A[717] * mat_B[425] +
//             mat_A[718] * mat_B[457] +
//             mat_A[719] * mat_B[489] +
//             mat_A[720] * mat_B[521] +
//             mat_A[721] * mat_B[553] +
//             mat_A[722] * mat_B[585] +
//             mat_A[723] * mat_B[617] +
//             mat_A[724] * mat_B[649] +
//             mat_A[725] * mat_B[681] +
//             mat_A[726] * mat_B[713] +
//             mat_A[727] * mat_B[745] +
//             mat_A[728] * mat_B[777] +
//             mat_A[729] * mat_B[809] +
//             mat_A[730] * mat_B[841] +
//             mat_A[731] * mat_B[873] +
//             mat_A[732] * mat_B[905] +
//             mat_A[733] * mat_B[937] +
//             mat_A[734] * mat_B[969] +
//             mat_A[735] * mat_B[1001];
//  mat_C[714] <= 
//             mat_A[704] * mat_B[10] +
//             mat_A[705] * mat_B[42] +
//             mat_A[706] * mat_B[74] +
//             mat_A[707] * mat_B[106] +
//             mat_A[708] * mat_B[138] +
//             mat_A[709] * mat_B[170] +
//             mat_A[710] * mat_B[202] +
//             mat_A[711] * mat_B[234] +
//             mat_A[712] * mat_B[266] +
//             mat_A[713] * mat_B[298] +
//             mat_A[714] * mat_B[330] +
//             mat_A[715] * mat_B[362] +
//             mat_A[716] * mat_B[394] +
//             mat_A[717] * mat_B[426] +
//             mat_A[718] * mat_B[458] +
//             mat_A[719] * mat_B[490] +
//             mat_A[720] * mat_B[522] +
//             mat_A[721] * mat_B[554] +
//             mat_A[722] * mat_B[586] +
//             mat_A[723] * mat_B[618] +
//             mat_A[724] * mat_B[650] +
//             mat_A[725] * mat_B[682] +
//             mat_A[726] * mat_B[714] +
//             mat_A[727] * mat_B[746] +
//             mat_A[728] * mat_B[778] +
//             mat_A[729] * mat_B[810] +
//             mat_A[730] * mat_B[842] +
//             mat_A[731] * mat_B[874] +
//             mat_A[732] * mat_B[906] +
//             mat_A[733] * mat_B[938] +
//             mat_A[734] * mat_B[970] +
//             mat_A[735] * mat_B[1002];
//  mat_C[715] <= 
//             mat_A[704] * mat_B[11] +
//             mat_A[705] * mat_B[43] +
//             mat_A[706] * mat_B[75] +
//             mat_A[707] * mat_B[107] +
//             mat_A[708] * mat_B[139] +
//             mat_A[709] * mat_B[171] +
//             mat_A[710] * mat_B[203] +
//             mat_A[711] * mat_B[235] +
//             mat_A[712] * mat_B[267] +
//             mat_A[713] * mat_B[299] +
//             mat_A[714] * mat_B[331] +
//             mat_A[715] * mat_B[363] +
//             mat_A[716] * mat_B[395] +
//             mat_A[717] * mat_B[427] +
//             mat_A[718] * mat_B[459] +
//             mat_A[719] * mat_B[491] +
//             mat_A[720] * mat_B[523] +
//             mat_A[721] * mat_B[555] +
//             mat_A[722] * mat_B[587] +
//             mat_A[723] * mat_B[619] +
//             mat_A[724] * mat_B[651] +
//             mat_A[725] * mat_B[683] +
//             mat_A[726] * mat_B[715] +
//             mat_A[727] * mat_B[747] +
//             mat_A[728] * mat_B[779] +
//             mat_A[729] * mat_B[811] +
//             mat_A[730] * mat_B[843] +
//             mat_A[731] * mat_B[875] +
//             mat_A[732] * mat_B[907] +
//             mat_A[733] * mat_B[939] +
//             mat_A[734] * mat_B[971] +
//             mat_A[735] * mat_B[1003];
//  mat_C[716] <= 
//             mat_A[704] * mat_B[12] +
//             mat_A[705] * mat_B[44] +
//             mat_A[706] * mat_B[76] +
//             mat_A[707] * mat_B[108] +
//             mat_A[708] * mat_B[140] +
//             mat_A[709] * mat_B[172] +
//             mat_A[710] * mat_B[204] +
//             mat_A[711] * mat_B[236] +
//             mat_A[712] * mat_B[268] +
//             mat_A[713] * mat_B[300] +
//             mat_A[714] * mat_B[332] +
//             mat_A[715] * mat_B[364] +
//             mat_A[716] * mat_B[396] +
//             mat_A[717] * mat_B[428] +
//             mat_A[718] * mat_B[460] +
//             mat_A[719] * mat_B[492] +
//             mat_A[720] * mat_B[524] +
//             mat_A[721] * mat_B[556] +
//             mat_A[722] * mat_B[588] +
//             mat_A[723] * mat_B[620] +
//             mat_A[724] * mat_B[652] +
//             mat_A[725] * mat_B[684] +
//             mat_A[726] * mat_B[716] +
//             mat_A[727] * mat_B[748] +
//             mat_A[728] * mat_B[780] +
//             mat_A[729] * mat_B[812] +
//             mat_A[730] * mat_B[844] +
//             mat_A[731] * mat_B[876] +
//             mat_A[732] * mat_B[908] +
//             mat_A[733] * mat_B[940] +
//             mat_A[734] * mat_B[972] +
//             mat_A[735] * mat_B[1004];
//  mat_C[717] <= 
//             mat_A[704] * mat_B[13] +
//             mat_A[705] * mat_B[45] +
//             mat_A[706] * mat_B[77] +
//             mat_A[707] * mat_B[109] +
//             mat_A[708] * mat_B[141] +
//             mat_A[709] * mat_B[173] +
//             mat_A[710] * mat_B[205] +
//             mat_A[711] * mat_B[237] +
//             mat_A[712] * mat_B[269] +
//             mat_A[713] * mat_B[301] +
//             mat_A[714] * mat_B[333] +
//             mat_A[715] * mat_B[365] +
//             mat_A[716] * mat_B[397] +
//             mat_A[717] * mat_B[429] +
//             mat_A[718] * mat_B[461] +
//             mat_A[719] * mat_B[493] +
//             mat_A[720] * mat_B[525] +
//             mat_A[721] * mat_B[557] +
//             mat_A[722] * mat_B[589] +
//             mat_A[723] * mat_B[621] +
//             mat_A[724] * mat_B[653] +
//             mat_A[725] * mat_B[685] +
//             mat_A[726] * mat_B[717] +
//             mat_A[727] * mat_B[749] +
//             mat_A[728] * mat_B[781] +
//             mat_A[729] * mat_B[813] +
//             mat_A[730] * mat_B[845] +
//             mat_A[731] * mat_B[877] +
//             mat_A[732] * mat_B[909] +
//             mat_A[733] * mat_B[941] +
//             mat_A[734] * mat_B[973] +
//             mat_A[735] * mat_B[1005];
//  mat_C[718] <= 
//             mat_A[704] * mat_B[14] +
//             mat_A[705] * mat_B[46] +
//             mat_A[706] * mat_B[78] +
//             mat_A[707] * mat_B[110] +
//             mat_A[708] * mat_B[142] +
//             mat_A[709] * mat_B[174] +
//             mat_A[710] * mat_B[206] +
//             mat_A[711] * mat_B[238] +
//             mat_A[712] * mat_B[270] +
//             mat_A[713] * mat_B[302] +
//             mat_A[714] * mat_B[334] +
//             mat_A[715] * mat_B[366] +
//             mat_A[716] * mat_B[398] +
//             mat_A[717] * mat_B[430] +
//             mat_A[718] * mat_B[462] +
//             mat_A[719] * mat_B[494] +
//             mat_A[720] * mat_B[526] +
//             mat_A[721] * mat_B[558] +
//             mat_A[722] * mat_B[590] +
//             mat_A[723] * mat_B[622] +
//             mat_A[724] * mat_B[654] +
//             mat_A[725] * mat_B[686] +
//             mat_A[726] * mat_B[718] +
//             mat_A[727] * mat_B[750] +
//             mat_A[728] * mat_B[782] +
//             mat_A[729] * mat_B[814] +
//             mat_A[730] * mat_B[846] +
//             mat_A[731] * mat_B[878] +
//             mat_A[732] * mat_B[910] +
//             mat_A[733] * mat_B[942] +
//             mat_A[734] * mat_B[974] +
//             mat_A[735] * mat_B[1006];
//  mat_C[719] <= 
//             mat_A[704] * mat_B[15] +
//             mat_A[705] * mat_B[47] +
//             mat_A[706] * mat_B[79] +
//             mat_A[707] * mat_B[111] +
//             mat_A[708] * mat_B[143] +
//             mat_A[709] * mat_B[175] +
//             mat_A[710] * mat_B[207] +
//             mat_A[711] * mat_B[239] +
//             mat_A[712] * mat_B[271] +
//             mat_A[713] * mat_B[303] +
//             mat_A[714] * mat_B[335] +
//             mat_A[715] * mat_B[367] +
//             mat_A[716] * mat_B[399] +
//             mat_A[717] * mat_B[431] +
//             mat_A[718] * mat_B[463] +
//             mat_A[719] * mat_B[495] +
//             mat_A[720] * mat_B[527] +
//             mat_A[721] * mat_B[559] +
//             mat_A[722] * mat_B[591] +
//             mat_A[723] * mat_B[623] +
//             mat_A[724] * mat_B[655] +
//             mat_A[725] * mat_B[687] +
//             mat_A[726] * mat_B[719] +
//             mat_A[727] * mat_B[751] +
//             mat_A[728] * mat_B[783] +
//             mat_A[729] * mat_B[815] +
//             mat_A[730] * mat_B[847] +
//             mat_A[731] * mat_B[879] +
//             mat_A[732] * mat_B[911] +
//             mat_A[733] * mat_B[943] +
//             mat_A[734] * mat_B[975] +
//             mat_A[735] * mat_B[1007];
//  mat_C[720] <= 
//             mat_A[704] * mat_B[16] +
//             mat_A[705] * mat_B[48] +
//             mat_A[706] * mat_B[80] +
//             mat_A[707] * mat_B[112] +
//             mat_A[708] * mat_B[144] +
//             mat_A[709] * mat_B[176] +
//             mat_A[710] * mat_B[208] +
//             mat_A[711] * mat_B[240] +
//             mat_A[712] * mat_B[272] +
//             mat_A[713] * mat_B[304] +
//             mat_A[714] * mat_B[336] +
//             mat_A[715] * mat_B[368] +
//             mat_A[716] * mat_B[400] +
//             mat_A[717] * mat_B[432] +
//             mat_A[718] * mat_B[464] +
//             mat_A[719] * mat_B[496] +
//             mat_A[720] * mat_B[528] +
//             mat_A[721] * mat_B[560] +
//             mat_A[722] * mat_B[592] +
//             mat_A[723] * mat_B[624] +
//             mat_A[724] * mat_B[656] +
//             mat_A[725] * mat_B[688] +
//             mat_A[726] * mat_B[720] +
//             mat_A[727] * mat_B[752] +
//             mat_A[728] * mat_B[784] +
//             mat_A[729] * mat_B[816] +
//             mat_A[730] * mat_B[848] +
//             mat_A[731] * mat_B[880] +
//             mat_A[732] * mat_B[912] +
//             mat_A[733] * mat_B[944] +
//             mat_A[734] * mat_B[976] +
//             mat_A[735] * mat_B[1008];
//  mat_C[721] <= 
//             mat_A[704] * mat_B[17] +
//             mat_A[705] * mat_B[49] +
//             mat_A[706] * mat_B[81] +
//             mat_A[707] * mat_B[113] +
//             mat_A[708] * mat_B[145] +
//             mat_A[709] * mat_B[177] +
//             mat_A[710] * mat_B[209] +
//             mat_A[711] * mat_B[241] +
//             mat_A[712] * mat_B[273] +
//             mat_A[713] * mat_B[305] +
//             mat_A[714] * mat_B[337] +
//             mat_A[715] * mat_B[369] +
//             mat_A[716] * mat_B[401] +
//             mat_A[717] * mat_B[433] +
//             mat_A[718] * mat_B[465] +
//             mat_A[719] * mat_B[497] +
//             mat_A[720] * mat_B[529] +
//             mat_A[721] * mat_B[561] +
//             mat_A[722] * mat_B[593] +
//             mat_A[723] * mat_B[625] +
//             mat_A[724] * mat_B[657] +
//             mat_A[725] * mat_B[689] +
//             mat_A[726] * mat_B[721] +
//             mat_A[727] * mat_B[753] +
//             mat_A[728] * mat_B[785] +
//             mat_A[729] * mat_B[817] +
//             mat_A[730] * mat_B[849] +
//             mat_A[731] * mat_B[881] +
//             mat_A[732] * mat_B[913] +
//             mat_A[733] * mat_B[945] +
//             mat_A[734] * mat_B[977] +
//             mat_A[735] * mat_B[1009];
//  mat_C[722] <= 
//             mat_A[704] * mat_B[18] +
//             mat_A[705] * mat_B[50] +
//             mat_A[706] * mat_B[82] +
//             mat_A[707] * mat_B[114] +
//             mat_A[708] * mat_B[146] +
//             mat_A[709] * mat_B[178] +
//             mat_A[710] * mat_B[210] +
//             mat_A[711] * mat_B[242] +
//             mat_A[712] * mat_B[274] +
//             mat_A[713] * mat_B[306] +
//             mat_A[714] * mat_B[338] +
//             mat_A[715] * mat_B[370] +
//             mat_A[716] * mat_B[402] +
//             mat_A[717] * mat_B[434] +
//             mat_A[718] * mat_B[466] +
//             mat_A[719] * mat_B[498] +
//             mat_A[720] * mat_B[530] +
//             mat_A[721] * mat_B[562] +
//             mat_A[722] * mat_B[594] +
//             mat_A[723] * mat_B[626] +
//             mat_A[724] * mat_B[658] +
//             mat_A[725] * mat_B[690] +
//             mat_A[726] * mat_B[722] +
//             mat_A[727] * mat_B[754] +
//             mat_A[728] * mat_B[786] +
//             mat_A[729] * mat_B[818] +
//             mat_A[730] * mat_B[850] +
//             mat_A[731] * mat_B[882] +
//             mat_A[732] * mat_B[914] +
//             mat_A[733] * mat_B[946] +
//             mat_A[734] * mat_B[978] +
//             mat_A[735] * mat_B[1010];
//  mat_C[723] <= 
//             mat_A[704] * mat_B[19] +
//             mat_A[705] * mat_B[51] +
//             mat_A[706] * mat_B[83] +
//             mat_A[707] * mat_B[115] +
//             mat_A[708] * mat_B[147] +
//             mat_A[709] * mat_B[179] +
//             mat_A[710] * mat_B[211] +
//             mat_A[711] * mat_B[243] +
//             mat_A[712] * mat_B[275] +
//             mat_A[713] * mat_B[307] +
//             mat_A[714] * mat_B[339] +
//             mat_A[715] * mat_B[371] +
//             mat_A[716] * mat_B[403] +
//             mat_A[717] * mat_B[435] +
//             mat_A[718] * mat_B[467] +
//             mat_A[719] * mat_B[499] +
//             mat_A[720] * mat_B[531] +
//             mat_A[721] * mat_B[563] +
//             mat_A[722] * mat_B[595] +
//             mat_A[723] * mat_B[627] +
//             mat_A[724] * mat_B[659] +
//             mat_A[725] * mat_B[691] +
//             mat_A[726] * mat_B[723] +
//             mat_A[727] * mat_B[755] +
//             mat_A[728] * mat_B[787] +
//             mat_A[729] * mat_B[819] +
//             mat_A[730] * mat_B[851] +
//             mat_A[731] * mat_B[883] +
//             mat_A[732] * mat_B[915] +
//             mat_A[733] * mat_B[947] +
//             mat_A[734] * mat_B[979] +
//             mat_A[735] * mat_B[1011];
//  mat_C[724] <= 
//             mat_A[704] * mat_B[20] +
//             mat_A[705] * mat_B[52] +
//             mat_A[706] * mat_B[84] +
//             mat_A[707] * mat_B[116] +
//             mat_A[708] * mat_B[148] +
//             mat_A[709] * mat_B[180] +
//             mat_A[710] * mat_B[212] +
//             mat_A[711] * mat_B[244] +
//             mat_A[712] * mat_B[276] +
//             mat_A[713] * mat_B[308] +
//             mat_A[714] * mat_B[340] +
//             mat_A[715] * mat_B[372] +
//             mat_A[716] * mat_B[404] +
//             mat_A[717] * mat_B[436] +
//             mat_A[718] * mat_B[468] +
//             mat_A[719] * mat_B[500] +
//             mat_A[720] * mat_B[532] +
//             mat_A[721] * mat_B[564] +
//             mat_A[722] * mat_B[596] +
//             mat_A[723] * mat_B[628] +
//             mat_A[724] * mat_B[660] +
//             mat_A[725] * mat_B[692] +
//             mat_A[726] * mat_B[724] +
//             mat_A[727] * mat_B[756] +
//             mat_A[728] * mat_B[788] +
//             mat_A[729] * mat_B[820] +
//             mat_A[730] * mat_B[852] +
//             mat_A[731] * mat_B[884] +
//             mat_A[732] * mat_B[916] +
//             mat_A[733] * mat_B[948] +
//             mat_A[734] * mat_B[980] +
//             mat_A[735] * mat_B[1012];
//  mat_C[725] <= 
//             mat_A[704] * mat_B[21] +
//             mat_A[705] * mat_B[53] +
//             mat_A[706] * mat_B[85] +
//             mat_A[707] * mat_B[117] +
//             mat_A[708] * mat_B[149] +
//             mat_A[709] * mat_B[181] +
//             mat_A[710] * mat_B[213] +
//             mat_A[711] * mat_B[245] +
//             mat_A[712] * mat_B[277] +
//             mat_A[713] * mat_B[309] +
//             mat_A[714] * mat_B[341] +
//             mat_A[715] * mat_B[373] +
//             mat_A[716] * mat_B[405] +
//             mat_A[717] * mat_B[437] +
//             mat_A[718] * mat_B[469] +
//             mat_A[719] * mat_B[501] +
//             mat_A[720] * mat_B[533] +
//             mat_A[721] * mat_B[565] +
//             mat_A[722] * mat_B[597] +
//             mat_A[723] * mat_B[629] +
//             mat_A[724] * mat_B[661] +
//             mat_A[725] * mat_B[693] +
//             mat_A[726] * mat_B[725] +
//             mat_A[727] * mat_B[757] +
//             mat_A[728] * mat_B[789] +
//             mat_A[729] * mat_B[821] +
//             mat_A[730] * mat_B[853] +
//             mat_A[731] * mat_B[885] +
//             mat_A[732] * mat_B[917] +
//             mat_A[733] * mat_B[949] +
//             mat_A[734] * mat_B[981] +
//             mat_A[735] * mat_B[1013];
//  mat_C[726] <= 
//             mat_A[704] * mat_B[22] +
//             mat_A[705] * mat_B[54] +
//             mat_A[706] * mat_B[86] +
//             mat_A[707] * mat_B[118] +
//             mat_A[708] * mat_B[150] +
//             mat_A[709] * mat_B[182] +
//             mat_A[710] * mat_B[214] +
//             mat_A[711] * mat_B[246] +
//             mat_A[712] * mat_B[278] +
//             mat_A[713] * mat_B[310] +
//             mat_A[714] * mat_B[342] +
//             mat_A[715] * mat_B[374] +
//             mat_A[716] * mat_B[406] +
//             mat_A[717] * mat_B[438] +
//             mat_A[718] * mat_B[470] +
//             mat_A[719] * mat_B[502] +
//             mat_A[720] * mat_B[534] +
//             mat_A[721] * mat_B[566] +
//             mat_A[722] * mat_B[598] +
//             mat_A[723] * mat_B[630] +
//             mat_A[724] * mat_B[662] +
//             mat_A[725] * mat_B[694] +
//             mat_A[726] * mat_B[726] +
//             mat_A[727] * mat_B[758] +
//             mat_A[728] * mat_B[790] +
//             mat_A[729] * mat_B[822] +
//             mat_A[730] * mat_B[854] +
//             mat_A[731] * mat_B[886] +
//             mat_A[732] * mat_B[918] +
//             mat_A[733] * mat_B[950] +
//             mat_A[734] * mat_B[982] +
//             mat_A[735] * mat_B[1014];
//  mat_C[727] <= 
//             mat_A[704] * mat_B[23] +
//             mat_A[705] * mat_B[55] +
//             mat_A[706] * mat_B[87] +
//             mat_A[707] * mat_B[119] +
//             mat_A[708] * mat_B[151] +
//             mat_A[709] * mat_B[183] +
//             mat_A[710] * mat_B[215] +
//             mat_A[711] * mat_B[247] +
//             mat_A[712] * mat_B[279] +
//             mat_A[713] * mat_B[311] +
//             mat_A[714] * mat_B[343] +
//             mat_A[715] * mat_B[375] +
//             mat_A[716] * mat_B[407] +
//             mat_A[717] * mat_B[439] +
//             mat_A[718] * mat_B[471] +
//             mat_A[719] * mat_B[503] +
//             mat_A[720] * mat_B[535] +
//             mat_A[721] * mat_B[567] +
//             mat_A[722] * mat_B[599] +
//             mat_A[723] * mat_B[631] +
//             mat_A[724] * mat_B[663] +
//             mat_A[725] * mat_B[695] +
//             mat_A[726] * mat_B[727] +
//             mat_A[727] * mat_B[759] +
//             mat_A[728] * mat_B[791] +
//             mat_A[729] * mat_B[823] +
//             mat_A[730] * mat_B[855] +
//             mat_A[731] * mat_B[887] +
//             mat_A[732] * mat_B[919] +
//             mat_A[733] * mat_B[951] +
//             mat_A[734] * mat_B[983] +
//             mat_A[735] * mat_B[1015];
//  mat_C[728] <= 
//             mat_A[704] * mat_B[24] +
//             mat_A[705] * mat_B[56] +
//             mat_A[706] * mat_B[88] +
//             mat_A[707] * mat_B[120] +
//             mat_A[708] * mat_B[152] +
//             mat_A[709] * mat_B[184] +
//             mat_A[710] * mat_B[216] +
//             mat_A[711] * mat_B[248] +
//             mat_A[712] * mat_B[280] +
//             mat_A[713] * mat_B[312] +
//             mat_A[714] * mat_B[344] +
//             mat_A[715] * mat_B[376] +
//             mat_A[716] * mat_B[408] +
//             mat_A[717] * mat_B[440] +
//             mat_A[718] * mat_B[472] +
//             mat_A[719] * mat_B[504] +
//             mat_A[720] * mat_B[536] +
//             mat_A[721] * mat_B[568] +
//             mat_A[722] * mat_B[600] +
//             mat_A[723] * mat_B[632] +
//             mat_A[724] * mat_B[664] +
//             mat_A[725] * mat_B[696] +
//             mat_A[726] * mat_B[728] +
//             mat_A[727] * mat_B[760] +
//             mat_A[728] * mat_B[792] +
//             mat_A[729] * mat_B[824] +
//             mat_A[730] * mat_B[856] +
//             mat_A[731] * mat_B[888] +
//             mat_A[732] * mat_B[920] +
//             mat_A[733] * mat_B[952] +
//             mat_A[734] * mat_B[984] +
//             mat_A[735] * mat_B[1016];
//  mat_C[729] <= 
//             mat_A[704] * mat_B[25] +
//             mat_A[705] * mat_B[57] +
//             mat_A[706] * mat_B[89] +
//             mat_A[707] * mat_B[121] +
//             mat_A[708] * mat_B[153] +
//             mat_A[709] * mat_B[185] +
//             mat_A[710] * mat_B[217] +
//             mat_A[711] * mat_B[249] +
//             mat_A[712] * mat_B[281] +
//             mat_A[713] * mat_B[313] +
//             mat_A[714] * mat_B[345] +
//             mat_A[715] * mat_B[377] +
//             mat_A[716] * mat_B[409] +
//             mat_A[717] * mat_B[441] +
//             mat_A[718] * mat_B[473] +
//             mat_A[719] * mat_B[505] +
//             mat_A[720] * mat_B[537] +
//             mat_A[721] * mat_B[569] +
//             mat_A[722] * mat_B[601] +
//             mat_A[723] * mat_B[633] +
//             mat_A[724] * mat_B[665] +
//             mat_A[725] * mat_B[697] +
//             mat_A[726] * mat_B[729] +
//             mat_A[727] * mat_B[761] +
//             mat_A[728] * mat_B[793] +
//             mat_A[729] * mat_B[825] +
//             mat_A[730] * mat_B[857] +
//             mat_A[731] * mat_B[889] +
//             mat_A[732] * mat_B[921] +
//             mat_A[733] * mat_B[953] +
//             mat_A[734] * mat_B[985] +
//             mat_A[735] * mat_B[1017];
//  mat_C[730] <= 
//             mat_A[704] * mat_B[26] +
//             mat_A[705] * mat_B[58] +
//             mat_A[706] * mat_B[90] +
//             mat_A[707] * mat_B[122] +
//             mat_A[708] * mat_B[154] +
//             mat_A[709] * mat_B[186] +
//             mat_A[710] * mat_B[218] +
//             mat_A[711] * mat_B[250] +
//             mat_A[712] * mat_B[282] +
//             mat_A[713] * mat_B[314] +
//             mat_A[714] * mat_B[346] +
//             mat_A[715] * mat_B[378] +
//             mat_A[716] * mat_B[410] +
//             mat_A[717] * mat_B[442] +
//             mat_A[718] * mat_B[474] +
//             mat_A[719] * mat_B[506] +
//             mat_A[720] * mat_B[538] +
//             mat_A[721] * mat_B[570] +
//             mat_A[722] * mat_B[602] +
//             mat_A[723] * mat_B[634] +
//             mat_A[724] * mat_B[666] +
//             mat_A[725] * mat_B[698] +
//             mat_A[726] * mat_B[730] +
//             mat_A[727] * mat_B[762] +
//             mat_A[728] * mat_B[794] +
//             mat_A[729] * mat_B[826] +
//             mat_A[730] * mat_B[858] +
//             mat_A[731] * mat_B[890] +
//             mat_A[732] * mat_B[922] +
//             mat_A[733] * mat_B[954] +
//             mat_A[734] * mat_B[986] +
//             mat_A[735] * mat_B[1018];
//  mat_C[731] <= 
//             mat_A[704] * mat_B[27] +
//             mat_A[705] * mat_B[59] +
//             mat_A[706] * mat_B[91] +
//             mat_A[707] * mat_B[123] +
//             mat_A[708] * mat_B[155] +
//             mat_A[709] * mat_B[187] +
//             mat_A[710] * mat_B[219] +
//             mat_A[711] * mat_B[251] +
//             mat_A[712] * mat_B[283] +
//             mat_A[713] * mat_B[315] +
//             mat_A[714] * mat_B[347] +
//             mat_A[715] * mat_B[379] +
//             mat_A[716] * mat_B[411] +
//             mat_A[717] * mat_B[443] +
//             mat_A[718] * mat_B[475] +
//             mat_A[719] * mat_B[507] +
//             mat_A[720] * mat_B[539] +
//             mat_A[721] * mat_B[571] +
//             mat_A[722] * mat_B[603] +
//             mat_A[723] * mat_B[635] +
//             mat_A[724] * mat_B[667] +
//             mat_A[725] * mat_B[699] +
//             mat_A[726] * mat_B[731] +
//             mat_A[727] * mat_B[763] +
//             mat_A[728] * mat_B[795] +
//             mat_A[729] * mat_B[827] +
//             mat_A[730] * mat_B[859] +
//             mat_A[731] * mat_B[891] +
//             mat_A[732] * mat_B[923] +
//             mat_A[733] * mat_B[955] +
//             mat_A[734] * mat_B[987] +
//             mat_A[735] * mat_B[1019];
//  mat_C[732] <= 
//             mat_A[704] * mat_B[28] +
//             mat_A[705] * mat_B[60] +
//             mat_A[706] * mat_B[92] +
//             mat_A[707] * mat_B[124] +
//             mat_A[708] * mat_B[156] +
//             mat_A[709] * mat_B[188] +
//             mat_A[710] * mat_B[220] +
//             mat_A[711] * mat_B[252] +
//             mat_A[712] * mat_B[284] +
//             mat_A[713] * mat_B[316] +
//             mat_A[714] * mat_B[348] +
//             mat_A[715] * mat_B[380] +
//             mat_A[716] * mat_B[412] +
//             mat_A[717] * mat_B[444] +
//             mat_A[718] * mat_B[476] +
//             mat_A[719] * mat_B[508] +
//             mat_A[720] * mat_B[540] +
//             mat_A[721] * mat_B[572] +
//             mat_A[722] * mat_B[604] +
//             mat_A[723] * mat_B[636] +
//             mat_A[724] * mat_B[668] +
//             mat_A[725] * mat_B[700] +
//             mat_A[726] * mat_B[732] +
//             mat_A[727] * mat_B[764] +
//             mat_A[728] * mat_B[796] +
//             mat_A[729] * mat_B[828] +
//             mat_A[730] * mat_B[860] +
//             mat_A[731] * mat_B[892] +
//             mat_A[732] * mat_B[924] +
//             mat_A[733] * mat_B[956] +
//             mat_A[734] * mat_B[988] +
//             mat_A[735] * mat_B[1020];
//  mat_C[733] <= 
//             mat_A[704] * mat_B[29] +
//             mat_A[705] * mat_B[61] +
//             mat_A[706] * mat_B[93] +
//             mat_A[707] * mat_B[125] +
//             mat_A[708] * mat_B[157] +
//             mat_A[709] * mat_B[189] +
//             mat_A[710] * mat_B[221] +
//             mat_A[711] * mat_B[253] +
//             mat_A[712] * mat_B[285] +
//             mat_A[713] * mat_B[317] +
//             mat_A[714] * mat_B[349] +
//             mat_A[715] * mat_B[381] +
//             mat_A[716] * mat_B[413] +
//             mat_A[717] * mat_B[445] +
//             mat_A[718] * mat_B[477] +
//             mat_A[719] * mat_B[509] +
//             mat_A[720] * mat_B[541] +
//             mat_A[721] * mat_B[573] +
//             mat_A[722] * mat_B[605] +
//             mat_A[723] * mat_B[637] +
//             mat_A[724] * mat_B[669] +
//             mat_A[725] * mat_B[701] +
//             mat_A[726] * mat_B[733] +
//             mat_A[727] * mat_B[765] +
//             mat_A[728] * mat_B[797] +
//             mat_A[729] * mat_B[829] +
//             mat_A[730] * mat_B[861] +
//             mat_A[731] * mat_B[893] +
//             mat_A[732] * mat_B[925] +
//             mat_A[733] * mat_B[957] +
//             mat_A[734] * mat_B[989] +
//             mat_A[735] * mat_B[1021];
//  mat_C[734] <= 
//             mat_A[704] * mat_B[30] +
//             mat_A[705] * mat_B[62] +
//             mat_A[706] * mat_B[94] +
//             mat_A[707] * mat_B[126] +
//             mat_A[708] * mat_B[158] +
//             mat_A[709] * mat_B[190] +
//             mat_A[710] * mat_B[222] +
//             mat_A[711] * mat_B[254] +
//             mat_A[712] * mat_B[286] +
//             mat_A[713] * mat_B[318] +
//             mat_A[714] * mat_B[350] +
//             mat_A[715] * mat_B[382] +
//             mat_A[716] * mat_B[414] +
//             mat_A[717] * mat_B[446] +
//             mat_A[718] * mat_B[478] +
//             mat_A[719] * mat_B[510] +
//             mat_A[720] * mat_B[542] +
//             mat_A[721] * mat_B[574] +
//             mat_A[722] * mat_B[606] +
//             mat_A[723] * mat_B[638] +
//             mat_A[724] * mat_B[670] +
//             mat_A[725] * mat_B[702] +
//             mat_A[726] * mat_B[734] +
//             mat_A[727] * mat_B[766] +
//             mat_A[728] * mat_B[798] +
//             mat_A[729] * mat_B[830] +
//             mat_A[730] * mat_B[862] +
//             mat_A[731] * mat_B[894] +
//             mat_A[732] * mat_B[926] +
//             mat_A[733] * mat_B[958] +
//             mat_A[734] * mat_B[990] +
//             mat_A[735] * mat_B[1022];
//  mat_C[735] <= 
//             mat_A[704] * mat_B[31] +
//             mat_A[705] * mat_B[63] +
//             mat_A[706] * mat_B[95] +
//             mat_A[707] * mat_B[127] +
//             mat_A[708] * mat_B[159] +
//             mat_A[709] * mat_B[191] +
//             mat_A[710] * mat_B[223] +
//             mat_A[711] * mat_B[255] +
//             mat_A[712] * mat_B[287] +
//             mat_A[713] * mat_B[319] +
//             mat_A[714] * mat_B[351] +
//             mat_A[715] * mat_B[383] +
//             mat_A[716] * mat_B[415] +
//             mat_A[717] * mat_B[447] +
//             mat_A[718] * mat_B[479] +
//             mat_A[719] * mat_B[511] +
//             mat_A[720] * mat_B[543] +
//             mat_A[721] * mat_B[575] +
//             mat_A[722] * mat_B[607] +
//             mat_A[723] * mat_B[639] +
//             mat_A[724] * mat_B[671] +
//             mat_A[725] * mat_B[703] +
//             mat_A[726] * mat_B[735] +
//             mat_A[727] * mat_B[767] +
//             mat_A[728] * mat_B[799] +
//             mat_A[729] * mat_B[831] +
//             mat_A[730] * mat_B[863] +
//             mat_A[731] * mat_B[895] +
//             mat_A[732] * mat_B[927] +
//             mat_A[733] * mat_B[959] +
//             mat_A[734] * mat_B[991] +
//             mat_A[735] * mat_B[1023];
//  mat_C[736] <= 
//             mat_A[736] * mat_B[0] +
//             mat_A[737] * mat_B[32] +
//             mat_A[738] * mat_B[64] +
//             mat_A[739] * mat_B[96] +
//             mat_A[740] * mat_B[128] +
//             mat_A[741] * mat_B[160] +
//             mat_A[742] * mat_B[192] +
//             mat_A[743] * mat_B[224] +
//             mat_A[744] * mat_B[256] +
//             mat_A[745] * mat_B[288] +
//             mat_A[746] * mat_B[320] +
//             mat_A[747] * mat_B[352] +
//             mat_A[748] * mat_B[384] +
//             mat_A[749] * mat_B[416] +
//             mat_A[750] * mat_B[448] +
//             mat_A[751] * mat_B[480] +
//             mat_A[752] * mat_B[512] +
//             mat_A[753] * mat_B[544] +
//             mat_A[754] * mat_B[576] +
//             mat_A[755] * mat_B[608] +
//             mat_A[756] * mat_B[640] +
//             mat_A[757] * mat_B[672] +
//             mat_A[758] * mat_B[704] +
//             mat_A[759] * mat_B[736] +
//             mat_A[760] * mat_B[768] +
//             mat_A[761] * mat_B[800] +
//             mat_A[762] * mat_B[832] +
//             mat_A[763] * mat_B[864] +
//             mat_A[764] * mat_B[896] +
//             mat_A[765] * mat_B[928] +
//             mat_A[766] * mat_B[960] +
//             mat_A[767] * mat_B[992];
//  mat_C[737] <= 
//             mat_A[736] * mat_B[1] +
//             mat_A[737] * mat_B[33] +
//             mat_A[738] * mat_B[65] +
//             mat_A[739] * mat_B[97] +
//             mat_A[740] * mat_B[129] +
//             mat_A[741] * mat_B[161] +
//             mat_A[742] * mat_B[193] +
//             mat_A[743] * mat_B[225] +
//             mat_A[744] * mat_B[257] +
//             mat_A[745] * mat_B[289] +
//             mat_A[746] * mat_B[321] +
//             mat_A[747] * mat_B[353] +
//             mat_A[748] * mat_B[385] +
//             mat_A[749] * mat_B[417] +
//             mat_A[750] * mat_B[449] +
//             mat_A[751] * mat_B[481] +
//             mat_A[752] * mat_B[513] +
//             mat_A[753] * mat_B[545] +
//             mat_A[754] * mat_B[577] +
//             mat_A[755] * mat_B[609] +
//             mat_A[756] * mat_B[641] +
//             mat_A[757] * mat_B[673] +
//             mat_A[758] * mat_B[705] +
//             mat_A[759] * mat_B[737] +
//             mat_A[760] * mat_B[769] +
//             mat_A[761] * mat_B[801] +
//             mat_A[762] * mat_B[833] +
//             mat_A[763] * mat_B[865] +
//             mat_A[764] * mat_B[897] +
//             mat_A[765] * mat_B[929] +
//             mat_A[766] * mat_B[961] +
//             mat_A[767] * mat_B[993];
//  mat_C[738] <= 
//             mat_A[736] * mat_B[2] +
//             mat_A[737] * mat_B[34] +
//             mat_A[738] * mat_B[66] +
//             mat_A[739] * mat_B[98] +
//             mat_A[740] * mat_B[130] +
//             mat_A[741] * mat_B[162] +
//             mat_A[742] * mat_B[194] +
//             mat_A[743] * mat_B[226] +
//             mat_A[744] * mat_B[258] +
//             mat_A[745] * mat_B[290] +
//             mat_A[746] * mat_B[322] +
//             mat_A[747] * mat_B[354] +
//             mat_A[748] * mat_B[386] +
//             mat_A[749] * mat_B[418] +
//             mat_A[750] * mat_B[450] +
//             mat_A[751] * mat_B[482] +
//             mat_A[752] * mat_B[514] +
//             mat_A[753] * mat_B[546] +
//             mat_A[754] * mat_B[578] +
//             mat_A[755] * mat_B[610] +
//             mat_A[756] * mat_B[642] +
//             mat_A[757] * mat_B[674] +
//             mat_A[758] * mat_B[706] +
//             mat_A[759] * mat_B[738] +
//             mat_A[760] * mat_B[770] +
//             mat_A[761] * mat_B[802] +
//             mat_A[762] * mat_B[834] +
//             mat_A[763] * mat_B[866] +
//             mat_A[764] * mat_B[898] +
//             mat_A[765] * mat_B[930] +
//             mat_A[766] * mat_B[962] +
//             mat_A[767] * mat_B[994];
//  mat_C[739] <= 
//             mat_A[736] * mat_B[3] +
//             mat_A[737] * mat_B[35] +
//             mat_A[738] * mat_B[67] +
//             mat_A[739] * mat_B[99] +
//             mat_A[740] * mat_B[131] +
//             mat_A[741] * mat_B[163] +
//             mat_A[742] * mat_B[195] +
//             mat_A[743] * mat_B[227] +
//             mat_A[744] * mat_B[259] +
//             mat_A[745] * mat_B[291] +
//             mat_A[746] * mat_B[323] +
//             mat_A[747] * mat_B[355] +
//             mat_A[748] * mat_B[387] +
//             mat_A[749] * mat_B[419] +
//             mat_A[750] * mat_B[451] +
//             mat_A[751] * mat_B[483] +
//             mat_A[752] * mat_B[515] +
//             mat_A[753] * mat_B[547] +
//             mat_A[754] * mat_B[579] +
//             mat_A[755] * mat_B[611] +
//             mat_A[756] * mat_B[643] +
//             mat_A[757] * mat_B[675] +
//             mat_A[758] * mat_B[707] +
//             mat_A[759] * mat_B[739] +
//             mat_A[760] * mat_B[771] +
//             mat_A[761] * mat_B[803] +
//             mat_A[762] * mat_B[835] +
//             mat_A[763] * mat_B[867] +
//             mat_A[764] * mat_B[899] +
//             mat_A[765] * mat_B[931] +
//             mat_A[766] * mat_B[963] +
//             mat_A[767] * mat_B[995];
//  mat_C[740] <= 
//             mat_A[736] * mat_B[4] +
//             mat_A[737] * mat_B[36] +
//             mat_A[738] * mat_B[68] +
//             mat_A[739] * mat_B[100] +
//             mat_A[740] * mat_B[132] +
//             mat_A[741] * mat_B[164] +
//             mat_A[742] * mat_B[196] +
//             mat_A[743] * mat_B[228] +
//             mat_A[744] * mat_B[260] +
//             mat_A[745] * mat_B[292] +
//             mat_A[746] * mat_B[324] +
//             mat_A[747] * mat_B[356] +
//             mat_A[748] * mat_B[388] +
//             mat_A[749] * mat_B[420] +
//             mat_A[750] * mat_B[452] +
//             mat_A[751] * mat_B[484] +
//             mat_A[752] * mat_B[516] +
//             mat_A[753] * mat_B[548] +
//             mat_A[754] * mat_B[580] +
//             mat_A[755] * mat_B[612] +
//             mat_A[756] * mat_B[644] +
//             mat_A[757] * mat_B[676] +
//             mat_A[758] * mat_B[708] +
//             mat_A[759] * mat_B[740] +
//             mat_A[760] * mat_B[772] +
//             mat_A[761] * mat_B[804] +
//             mat_A[762] * mat_B[836] +
//             mat_A[763] * mat_B[868] +
//             mat_A[764] * mat_B[900] +
//             mat_A[765] * mat_B[932] +
//             mat_A[766] * mat_B[964] +
//             mat_A[767] * mat_B[996];
//  mat_C[741] <= 
//             mat_A[736] * mat_B[5] +
//             mat_A[737] * mat_B[37] +
//             mat_A[738] * mat_B[69] +
//             mat_A[739] * mat_B[101] +
//             mat_A[740] * mat_B[133] +
//             mat_A[741] * mat_B[165] +
//             mat_A[742] * mat_B[197] +
//             mat_A[743] * mat_B[229] +
//             mat_A[744] * mat_B[261] +
//             mat_A[745] * mat_B[293] +
//             mat_A[746] * mat_B[325] +
//             mat_A[747] * mat_B[357] +
//             mat_A[748] * mat_B[389] +
//             mat_A[749] * mat_B[421] +
//             mat_A[750] * mat_B[453] +
//             mat_A[751] * mat_B[485] +
//             mat_A[752] * mat_B[517] +
//             mat_A[753] * mat_B[549] +
//             mat_A[754] * mat_B[581] +
//             mat_A[755] * mat_B[613] +
//             mat_A[756] * mat_B[645] +
//             mat_A[757] * mat_B[677] +
//             mat_A[758] * mat_B[709] +
//             mat_A[759] * mat_B[741] +
//             mat_A[760] * mat_B[773] +
//             mat_A[761] * mat_B[805] +
//             mat_A[762] * mat_B[837] +
//             mat_A[763] * mat_B[869] +
//             mat_A[764] * mat_B[901] +
//             mat_A[765] * mat_B[933] +
//             mat_A[766] * mat_B[965] +
//             mat_A[767] * mat_B[997];
//  mat_C[742] <= 
//             mat_A[736] * mat_B[6] +
//             mat_A[737] * mat_B[38] +
//             mat_A[738] * mat_B[70] +
//             mat_A[739] * mat_B[102] +
//             mat_A[740] * mat_B[134] +
//             mat_A[741] * mat_B[166] +
//             mat_A[742] * mat_B[198] +
//             mat_A[743] * mat_B[230] +
//             mat_A[744] * mat_B[262] +
//             mat_A[745] * mat_B[294] +
//             mat_A[746] * mat_B[326] +
//             mat_A[747] * mat_B[358] +
//             mat_A[748] * mat_B[390] +
//             mat_A[749] * mat_B[422] +
//             mat_A[750] * mat_B[454] +
//             mat_A[751] * mat_B[486] +
//             mat_A[752] * mat_B[518] +
//             mat_A[753] * mat_B[550] +
//             mat_A[754] * mat_B[582] +
//             mat_A[755] * mat_B[614] +
//             mat_A[756] * mat_B[646] +
//             mat_A[757] * mat_B[678] +
//             mat_A[758] * mat_B[710] +
//             mat_A[759] * mat_B[742] +
//             mat_A[760] * mat_B[774] +
//             mat_A[761] * mat_B[806] +
//             mat_A[762] * mat_B[838] +
//             mat_A[763] * mat_B[870] +
//             mat_A[764] * mat_B[902] +
//             mat_A[765] * mat_B[934] +
//             mat_A[766] * mat_B[966] +
//             mat_A[767] * mat_B[998];
//  mat_C[743] <= 
//             mat_A[736] * mat_B[7] +
//             mat_A[737] * mat_B[39] +
//             mat_A[738] * mat_B[71] +
//             mat_A[739] * mat_B[103] +
//             mat_A[740] * mat_B[135] +
//             mat_A[741] * mat_B[167] +
//             mat_A[742] * mat_B[199] +
//             mat_A[743] * mat_B[231] +
//             mat_A[744] * mat_B[263] +
//             mat_A[745] * mat_B[295] +
//             mat_A[746] * mat_B[327] +
//             mat_A[747] * mat_B[359] +
//             mat_A[748] * mat_B[391] +
//             mat_A[749] * mat_B[423] +
//             mat_A[750] * mat_B[455] +
//             mat_A[751] * mat_B[487] +
//             mat_A[752] * mat_B[519] +
//             mat_A[753] * mat_B[551] +
//             mat_A[754] * mat_B[583] +
//             mat_A[755] * mat_B[615] +
//             mat_A[756] * mat_B[647] +
//             mat_A[757] * mat_B[679] +
//             mat_A[758] * mat_B[711] +
//             mat_A[759] * mat_B[743] +
//             mat_A[760] * mat_B[775] +
//             mat_A[761] * mat_B[807] +
//             mat_A[762] * mat_B[839] +
//             mat_A[763] * mat_B[871] +
//             mat_A[764] * mat_B[903] +
//             mat_A[765] * mat_B[935] +
//             mat_A[766] * mat_B[967] +
//             mat_A[767] * mat_B[999];
//  mat_C[744] <= 
//             mat_A[736] * mat_B[8] +
//             mat_A[737] * mat_B[40] +
//             mat_A[738] * mat_B[72] +
//             mat_A[739] * mat_B[104] +
//             mat_A[740] * mat_B[136] +
//             mat_A[741] * mat_B[168] +
//             mat_A[742] * mat_B[200] +
//             mat_A[743] * mat_B[232] +
//             mat_A[744] * mat_B[264] +
//             mat_A[745] * mat_B[296] +
//             mat_A[746] * mat_B[328] +
//             mat_A[747] * mat_B[360] +
//             mat_A[748] * mat_B[392] +
//             mat_A[749] * mat_B[424] +
//             mat_A[750] * mat_B[456] +
//             mat_A[751] * mat_B[488] +
//             mat_A[752] * mat_B[520] +
//             mat_A[753] * mat_B[552] +
//             mat_A[754] * mat_B[584] +
//             mat_A[755] * mat_B[616] +
//             mat_A[756] * mat_B[648] +
//             mat_A[757] * mat_B[680] +
//             mat_A[758] * mat_B[712] +
//             mat_A[759] * mat_B[744] +
//             mat_A[760] * mat_B[776] +
//             mat_A[761] * mat_B[808] +
//             mat_A[762] * mat_B[840] +
//             mat_A[763] * mat_B[872] +
//             mat_A[764] * mat_B[904] +
//             mat_A[765] * mat_B[936] +
//             mat_A[766] * mat_B[968] +
//             mat_A[767] * mat_B[1000];
//  mat_C[745] <= 
//             mat_A[736] * mat_B[9] +
//             mat_A[737] * mat_B[41] +
//             mat_A[738] * mat_B[73] +
//             mat_A[739] * mat_B[105] +
//             mat_A[740] * mat_B[137] +
//             mat_A[741] * mat_B[169] +
//             mat_A[742] * mat_B[201] +
//             mat_A[743] * mat_B[233] +
//             mat_A[744] * mat_B[265] +
//             mat_A[745] * mat_B[297] +
//             mat_A[746] * mat_B[329] +
//             mat_A[747] * mat_B[361] +
//             mat_A[748] * mat_B[393] +
//             mat_A[749] * mat_B[425] +
//             mat_A[750] * mat_B[457] +
//             mat_A[751] * mat_B[489] +
//             mat_A[752] * mat_B[521] +
//             mat_A[753] * mat_B[553] +
//             mat_A[754] * mat_B[585] +
//             mat_A[755] * mat_B[617] +
//             mat_A[756] * mat_B[649] +
//             mat_A[757] * mat_B[681] +
//             mat_A[758] * mat_B[713] +
//             mat_A[759] * mat_B[745] +
//             mat_A[760] * mat_B[777] +
//             mat_A[761] * mat_B[809] +
//             mat_A[762] * mat_B[841] +
//             mat_A[763] * mat_B[873] +
//             mat_A[764] * mat_B[905] +
//             mat_A[765] * mat_B[937] +
//             mat_A[766] * mat_B[969] +
//             mat_A[767] * mat_B[1001];
//  mat_C[746] <= 
//             mat_A[736] * mat_B[10] +
//             mat_A[737] * mat_B[42] +
//             mat_A[738] * mat_B[74] +
//             mat_A[739] * mat_B[106] +
//             mat_A[740] * mat_B[138] +
//             mat_A[741] * mat_B[170] +
//             mat_A[742] * mat_B[202] +
//             mat_A[743] * mat_B[234] +
//             mat_A[744] * mat_B[266] +
//             mat_A[745] * mat_B[298] +
//             mat_A[746] * mat_B[330] +
//             mat_A[747] * mat_B[362] +
//             mat_A[748] * mat_B[394] +
//             mat_A[749] * mat_B[426] +
//             mat_A[750] * mat_B[458] +
//             mat_A[751] * mat_B[490] +
//             mat_A[752] * mat_B[522] +
//             mat_A[753] * mat_B[554] +
//             mat_A[754] * mat_B[586] +
//             mat_A[755] * mat_B[618] +
//             mat_A[756] * mat_B[650] +
//             mat_A[757] * mat_B[682] +
//             mat_A[758] * mat_B[714] +
//             mat_A[759] * mat_B[746] +
//             mat_A[760] * mat_B[778] +
//             mat_A[761] * mat_B[810] +
//             mat_A[762] * mat_B[842] +
//             mat_A[763] * mat_B[874] +
//             mat_A[764] * mat_B[906] +
//             mat_A[765] * mat_B[938] +
//             mat_A[766] * mat_B[970] +
//             mat_A[767] * mat_B[1002];
//  mat_C[747] <= 
//             mat_A[736] * mat_B[11] +
//             mat_A[737] * mat_B[43] +
//             mat_A[738] * mat_B[75] +
//             mat_A[739] * mat_B[107] +
//             mat_A[740] * mat_B[139] +
//             mat_A[741] * mat_B[171] +
//             mat_A[742] * mat_B[203] +
//             mat_A[743] * mat_B[235] +
//             mat_A[744] * mat_B[267] +
//             mat_A[745] * mat_B[299] +
//             mat_A[746] * mat_B[331] +
//             mat_A[747] * mat_B[363] +
//             mat_A[748] * mat_B[395] +
//             mat_A[749] * mat_B[427] +
//             mat_A[750] * mat_B[459] +
//             mat_A[751] * mat_B[491] +
//             mat_A[752] * mat_B[523] +
//             mat_A[753] * mat_B[555] +
//             mat_A[754] * mat_B[587] +
//             mat_A[755] * mat_B[619] +
//             mat_A[756] * mat_B[651] +
//             mat_A[757] * mat_B[683] +
//             mat_A[758] * mat_B[715] +
//             mat_A[759] * mat_B[747] +
//             mat_A[760] * mat_B[779] +
//             mat_A[761] * mat_B[811] +
//             mat_A[762] * mat_B[843] +
//             mat_A[763] * mat_B[875] +
//             mat_A[764] * mat_B[907] +
//             mat_A[765] * mat_B[939] +
//             mat_A[766] * mat_B[971] +
//             mat_A[767] * mat_B[1003];
//  mat_C[748] <= 
//             mat_A[736] * mat_B[12] +
//             mat_A[737] * mat_B[44] +
//             mat_A[738] * mat_B[76] +
//             mat_A[739] * mat_B[108] +
//             mat_A[740] * mat_B[140] +
//             mat_A[741] * mat_B[172] +
//             mat_A[742] * mat_B[204] +
//             mat_A[743] * mat_B[236] +
//             mat_A[744] * mat_B[268] +
//             mat_A[745] * mat_B[300] +
//             mat_A[746] * mat_B[332] +
//             mat_A[747] * mat_B[364] +
//             mat_A[748] * mat_B[396] +
//             mat_A[749] * mat_B[428] +
//             mat_A[750] * mat_B[460] +
//             mat_A[751] * mat_B[492] +
//             mat_A[752] * mat_B[524] +
//             mat_A[753] * mat_B[556] +
//             mat_A[754] * mat_B[588] +
//             mat_A[755] * mat_B[620] +
//             mat_A[756] * mat_B[652] +
//             mat_A[757] * mat_B[684] +
//             mat_A[758] * mat_B[716] +
//             mat_A[759] * mat_B[748] +
//             mat_A[760] * mat_B[780] +
//             mat_A[761] * mat_B[812] +
//             mat_A[762] * mat_B[844] +
//             mat_A[763] * mat_B[876] +
//             mat_A[764] * mat_B[908] +
//             mat_A[765] * mat_B[940] +
//             mat_A[766] * mat_B[972] +
//             mat_A[767] * mat_B[1004];
//  mat_C[749] <= 
//             mat_A[736] * mat_B[13] +
//             mat_A[737] * mat_B[45] +
//             mat_A[738] * mat_B[77] +
//             mat_A[739] * mat_B[109] +
//             mat_A[740] * mat_B[141] +
//             mat_A[741] * mat_B[173] +
//             mat_A[742] * mat_B[205] +
//             mat_A[743] * mat_B[237] +
//             mat_A[744] * mat_B[269] +
//             mat_A[745] * mat_B[301] +
//             mat_A[746] * mat_B[333] +
//             mat_A[747] * mat_B[365] +
//             mat_A[748] * mat_B[397] +
//             mat_A[749] * mat_B[429] +
//             mat_A[750] * mat_B[461] +
//             mat_A[751] * mat_B[493] +
//             mat_A[752] * mat_B[525] +
//             mat_A[753] * mat_B[557] +
//             mat_A[754] * mat_B[589] +
//             mat_A[755] * mat_B[621] +
//             mat_A[756] * mat_B[653] +
//             mat_A[757] * mat_B[685] +
//             mat_A[758] * mat_B[717] +
//             mat_A[759] * mat_B[749] +
//             mat_A[760] * mat_B[781] +
//             mat_A[761] * mat_B[813] +
//             mat_A[762] * mat_B[845] +
//             mat_A[763] * mat_B[877] +
//             mat_A[764] * mat_B[909] +
//             mat_A[765] * mat_B[941] +
//             mat_A[766] * mat_B[973] +
//             mat_A[767] * mat_B[1005];
//  mat_C[750] <= 
//             mat_A[736] * mat_B[14] +
//             mat_A[737] * mat_B[46] +
//             mat_A[738] * mat_B[78] +
//             mat_A[739] * mat_B[110] +
//             mat_A[740] * mat_B[142] +
//             mat_A[741] * mat_B[174] +
//             mat_A[742] * mat_B[206] +
//             mat_A[743] * mat_B[238] +
//             mat_A[744] * mat_B[270] +
//             mat_A[745] * mat_B[302] +
//             mat_A[746] * mat_B[334] +
//             mat_A[747] * mat_B[366] +
//             mat_A[748] * mat_B[398] +
//             mat_A[749] * mat_B[430] +
//             mat_A[750] * mat_B[462] +
//             mat_A[751] * mat_B[494] +
//             mat_A[752] * mat_B[526] +
//             mat_A[753] * mat_B[558] +
//             mat_A[754] * mat_B[590] +
//             mat_A[755] * mat_B[622] +
//             mat_A[756] * mat_B[654] +
//             mat_A[757] * mat_B[686] +
//             mat_A[758] * mat_B[718] +
//             mat_A[759] * mat_B[750] +
//             mat_A[760] * mat_B[782] +
//             mat_A[761] * mat_B[814] +
//             mat_A[762] * mat_B[846] +
//             mat_A[763] * mat_B[878] +
//             mat_A[764] * mat_B[910] +
//             mat_A[765] * mat_B[942] +
//             mat_A[766] * mat_B[974] +
//             mat_A[767] * mat_B[1006];
//  mat_C[751] <= 
//             mat_A[736] * mat_B[15] +
//             mat_A[737] * mat_B[47] +
//             mat_A[738] * mat_B[79] +
//             mat_A[739] * mat_B[111] +
//             mat_A[740] * mat_B[143] +
//             mat_A[741] * mat_B[175] +
//             mat_A[742] * mat_B[207] +
//             mat_A[743] * mat_B[239] +
//             mat_A[744] * mat_B[271] +
//             mat_A[745] * mat_B[303] +
//             mat_A[746] * mat_B[335] +
//             mat_A[747] * mat_B[367] +
//             mat_A[748] * mat_B[399] +
//             mat_A[749] * mat_B[431] +
//             mat_A[750] * mat_B[463] +
//             mat_A[751] * mat_B[495] +
//             mat_A[752] * mat_B[527] +
//             mat_A[753] * mat_B[559] +
//             mat_A[754] * mat_B[591] +
//             mat_A[755] * mat_B[623] +
//             mat_A[756] * mat_B[655] +
//             mat_A[757] * mat_B[687] +
//             mat_A[758] * mat_B[719] +
//             mat_A[759] * mat_B[751] +
//             mat_A[760] * mat_B[783] +
//             mat_A[761] * mat_B[815] +
//             mat_A[762] * mat_B[847] +
//             mat_A[763] * mat_B[879] +
//             mat_A[764] * mat_B[911] +
//             mat_A[765] * mat_B[943] +
//             mat_A[766] * mat_B[975] +
//             mat_A[767] * mat_B[1007];
//  mat_C[752] <= 
//             mat_A[736] * mat_B[16] +
//             mat_A[737] * mat_B[48] +
//             mat_A[738] * mat_B[80] +
//             mat_A[739] * mat_B[112] +
//             mat_A[740] * mat_B[144] +
//             mat_A[741] * mat_B[176] +
//             mat_A[742] * mat_B[208] +
//             mat_A[743] * mat_B[240] +
//             mat_A[744] * mat_B[272] +
//             mat_A[745] * mat_B[304] +
//             mat_A[746] * mat_B[336] +
//             mat_A[747] * mat_B[368] +
//             mat_A[748] * mat_B[400] +
//             mat_A[749] * mat_B[432] +
//             mat_A[750] * mat_B[464] +
//             mat_A[751] * mat_B[496] +
//             mat_A[752] * mat_B[528] +
//             mat_A[753] * mat_B[560] +
//             mat_A[754] * mat_B[592] +
//             mat_A[755] * mat_B[624] +
//             mat_A[756] * mat_B[656] +
//             mat_A[757] * mat_B[688] +
//             mat_A[758] * mat_B[720] +
//             mat_A[759] * mat_B[752] +
//             mat_A[760] * mat_B[784] +
//             mat_A[761] * mat_B[816] +
//             mat_A[762] * mat_B[848] +
//             mat_A[763] * mat_B[880] +
//             mat_A[764] * mat_B[912] +
//             mat_A[765] * mat_B[944] +
//             mat_A[766] * mat_B[976] +
//             mat_A[767] * mat_B[1008];
//  mat_C[753] <= 
//             mat_A[736] * mat_B[17] +
//             mat_A[737] * mat_B[49] +
//             mat_A[738] * mat_B[81] +
//             mat_A[739] * mat_B[113] +
//             mat_A[740] * mat_B[145] +
//             mat_A[741] * mat_B[177] +
//             mat_A[742] * mat_B[209] +
//             mat_A[743] * mat_B[241] +
//             mat_A[744] * mat_B[273] +
//             mat_A[745] * mat_B[305] +
//             mat_A[746] * mat_B[337] +
//             mat_A[747] * mat_B[369] +
//             mat_A[748] * mat_B[401] +
//             mat_A[749] * mat_B[433] +
//             mat_A[750] * mat_B[465] +
//             mat_A[751] * mat_B[497] +
//             mat_A[752] * mat_B[529] +
//             mat_A[753] * mat_B[561] +
//             mat_A[754] * mat_B[593] +
//             mat_A[755] * mat_B[625] +
//             mat_A[756] * mat_B[657] +
//             mat_A[757] * mat_B[689] +
//             mat_A[758] * mat_B[721] +
//             mat_A[759] * mat_B[753] +
//             mat_A[760] * mat_B[785] +
//             mat_A[761] * mat_B[817] +
//             mat_A[762] * mat_B[849] +
//             mat_A[763] * mat_B[881] +
//             mat_A[764] * mat_B[913] +
//             mat_A[765] * mat_B[945] +
//             mat_A[766] * mat_B[977] +
//             mat_A[767] * mat_B[1009];
//  mat_C[754] <= 
//             mat_A[736] * mat_B[18] +
//             mat_A[737] * mat_B[50] +
//             mat_A[738] * mat_B[82] +
//             mat_A[739] * mat_B[114] +
//             mat_A[740] * mat_B[146] +
//             mat_A[741] * mat_B[178] +
//             mat_A[742] * mat_B[210] +
//             mat_A[743] * mat_B[242] +
//             mat_A[744] * mat_B[274] +
//             mat_A[745] * mat_B[306] +
//             mat_A[746] * mat_B[338] +
//             mat_A[747] * mat_B[370] +
//             mat_A[748] * mat_B[402] +
//             mat_A[749] * mat_B[434] +
//             mat_A[750] * mat_B[466] +
//             mat_A[751] * mat_B[498] +
//             mat_A[752] * mat_B[530] +
//             mat_A[753] * mat_B[562] +
//             mat_A[754] * mat_B[594] +
//             mat_A[755] * mat_B[626] +
//             mat_A[756] * mat_B[658] +
//             mat_A[757] * mat_B[690] +
//             mat_A[758] * mat_B[722] +
//             mat_A[759] * mat_B[754] +
//             mat_A[760] * mat_B[786] +
//             mat_A[761] * mat_B[818] +
//             mat_A[762] * mat_B[850] +
//             mat_A[763] * mat_B[882] +
//             mat_A[764] * mat_B[914] +
//             mat_A[765] * mat_B[946] +
//             mat_A[766] * mat_B[978] +
//             mat_A[767] * mat_B[1010];
//  mat_C[755] <= 
//             mat_A[736] * mat_B[19] +
//             mat_A[737] * mat_B[51] +
//             mat_A[738] * mat_B[83] +
//             mat_A[739] * mat_B[115] +
//             mat_A[740] * mat_B[147] +
//             mat_A[741] * mat_B[179] +
//             mat_A[742] * mat_B[211] +
//             mat_A[743] * mat_B[243] +
//             mat_A[744] * mat_B[275] +
//             mat_A[745] * mat_B[307] +
//             mat_A[746] * mat_B[339] +
//             mat_A[747] * mat_B[371] +
//             mat_A[748] * mat_B[403] +
//             mat_A[749] * mat_B[435] +
//             mat_A[750] * mat_B[467] +
//             mat_A[751] * mat_B[499] +
//             mat_A[752] * mat_B[531] +
//             mat_A[753] * mat_B[563] +
//             mat_A[754] * mat_B[595] +
//             mat_A[755] * mat_B[627] +
//             mat_A[756] * mat_B[659] +
//             mat_A[757] * mat_B[691] +
//             mat_A[758] * mat_B[723] +
//             mat_A[759] * mat_B[755] +
//             mat_A[760] * mat_B[787] +
//             mat_A[761] * mat_B[819] +
//             mat_A[762] * mat_B[851] +
//             mat_A[763] * mat_B[883] +
//             mat_A[764] * mat_B[915] +
//             mat_A[765] * mat_B[947] +
//             mat_A[766] * mat_B[979] +
//             mat_A[767] * mat_B[1011];
//  mat_C[756] <= 
//             mat_A[736] * mat_B[20] +
//             mat_A[737] * mat_B[52] +
//             mat_A[738] * mat_B[84] +
//             mat_A[739] * mat_B[116] +
//             mat_A[740] * mat_B[148] +
//             mat_A[741] * mat_B[180] +
//             mat_A[742] * mat_B[212] +
//             mat_A[743] * mat_B[244] +
//             mat_A[744] * mat_B[276] +
//             mat_A[745] * mat_B[308] +
//             mat_A[746] * mat_B[340] +
//             mat_A[747] * mat_B[372] +
//             mat_A[748] * mat_B[404] +
//             mat_A[749] * mat_B[436] +
//             mat_A[750] * mat_B[468] +
//             mat_A[751] * mat_B[500] +
//             mat_A[752] * mat_B[532] +
//             mat_A[753] * mat_B[564] +
//             mat_A[754] * mat_B[596] +
//             mat_A[755] * mat_B[628] +
//             mat_A[756] * mat_B[660] +
//             mat_A[757] * mat_B[692] +
//             mat_A[758] * mat_B[724] +
//             mat_A[759] * mat_B[756] +
//             mat_A[760] * mat_B[788] +
//             mat_A[761] * mat_B[820] +
//             mat_A[762] * mat_B[852] +
//             mat_A[763] * mat_B[884] +
//             mat_A[764] * mat_B[916] +
//             mat_A[765] * mat_B[948] +
//             mat_A[766] * mat_B[980] +
//             mat_A[767] * mat_B[1012];
//  mat_C[757] <= 
//             mat_A[736] * mat_B[21] +
//             mat_A[737] * mat_B[53] +
//             mat_A[738] * mat_B[85] +
//             mat_A[739] * mat_B[117] +
//             mat_A[740] * mat_B[149] +
//             mat_A[741] * mat_B[181] +
//             mat_A[742] * mat_B[213] +
//             mat_A[743] * mat_B[245] +
//             mat_A[744] * mat_B[277] +
//             mat_A[745] * mat_B[309] +
//             mat_A[746] * mat_B[341] +
//             mat_A[747] * mat_B[373] +
//             mat_A[748] * mat_B[405] +
//             mat_A[749] * mat_B[437] +
//             mat_A[750] * mat_B[469] +
//             mat_A[751] * mat_B[501] +
//             mat_A[752] * mat_B[533] +
//             mat_A[753] * mat_B[565] +
//             mat_A[754] * mat_B[597] +
//             mat_A[755] * mat_B[629] +
//             mat_A[756] * mat_B[661] +
//             mat_A[757] * mat_B[693] +
//             mat_A[758] * mat_B[725] +
//             mat_A[759] * mat_B[757] +
//             mat_A[760] * mat_B[789] +
//             mat_A[761] * mat_B[821] +
//             mat_A[762] * mat_B[853] +
//             mat_A[763] * mat_B[885] +
//             mat_A[764] * mat_B[917] +
//             mat_A[765] * mat_B[949] +
//             mat_A[766] * mat_B[981] +
//             mat_A[767] * mat_B[1013];
//  mat_C[758] <= 
//             mat_A[736] * mat_B[22] +
//             mat_A[737] * mat_B[54] +
//             mat_A[738] * mat_B[86] +
//             mat_A[739] * mat_B[118] +
//             mat_A[740] * mat_B[150] +
//             mat_A[741] * mat_B[182] +
//             mat_A[742] * mat_B[214] +
//             mat_A[743] * mat_B[246] +
//             mat_A[744] * mat_B[278] +
//             mat_A[745] * mat_B[310] +
//             mat_A[746] * mat_B[342] +
//             mat_A[747] * mat_B[374] +
//             mat_A[748] * mat_B[406] +
//             mat_A[749] * mat_B[438] +
//             mat_A[750] * mat_B[470] +
//             mat_A[751] * mat_B[502] +
//             mat_A[752] * mat_B[534] +
//             mat_A[753] * mat_B[566] +
//             mat_A[754] * mat_B[598] +
//             mat_A[755] * mat_B[630] +
//             mat_A[756] * mat_B[662] +
//             mat_A[757] * mat_B[694] +
//             mat_A[758] * mat_B[726] +
//             mat_A[759] * mat_B[758] +
//             mat_A[760] * mat_B[790] +
//             mat_A[761] * mat_B[822] +
//             mat_A[762] * mat_B[854] +
//             mat_A[763] * mat_B[886] +
//             mat_A[764] * mat_B[918] +
//             mat_A[765] * mat_B[950] +
//             mat_A[766] * mat_B[982] +
//             mat_A[767] * mat_B[1014];
//  mat_C[759] <= 
//             mat_A[736] * mat_B[23] +
//             mat_A[737] * mat_B[55] +
//             mat_A[738] * mat_B[87] +
//             mat_A[739] * mat_B[119] +
//             mat_A[740] * mat_B[151] +
//             mat_A[741] * mat_B[183] +
//             mat_A[742] * mat_B[215] +
//             mat_A[743] * mat_B[247] +
//             mat_A[744] * mat_B[279] +
//             mat_A[745] * mat_B[311] +
//             mat_A[746] * mat_B[343] +
//             mat_A[747] * mat_B[375] +
//             mat_A[748] * mat_B[407] +
//             mat_A[749] * mat_B[439] +
//             mat_A[750] * mat_B[471] +
//             mat_A[751] * mat_B[503] +
//             mat_A[752] * mat_B[535] +
//             mat_A[753] * mat_B[567] +
//             mat_A[754] * mat_B[599] +
//             mat_A[755] * mat_B[631] +
//             mat_A[756] * mat_B[663] +
//             mat_A[757] * mat_B[695] +
//             mat_A[758] * mat_B[727] +
//             mat_A[759] * mat_B[759] +
//             mat_A[760] * mat_B[791] +
//             mat_A[761] * mat_B[823] +
//             mat_A[762] * mat_B[855] +
//             mat_A[763] * mat_B[887] +
//             mat_A[764] * mat_B[919] +
//             mat_A[765] * mat_B[951] +
//             mat_A[766] * mat_B[983] +
//             mat_A[767] * mat_B[1015];
//  mat_C[760] <= 
//             mat_A[736] * mat_B[24] +
//             mat_A[737] * mat_B[56] +
//             mat_A[738] * mat_B[88] +
//             mat_A[739] * mat_B[120] +
//             mat_A[740] * mat_B[152] +
//             mat_A[741] * mat_B[184] +
//             mat_A[742] * mat_B[216] +
//             mat_A[743] * mat_B[248] +
//             mat_A[744] * mat_B[280] +
//             mat_A[745] * mat_B[312] +
//             mat_A[746] * mat_B[344] +
//             mat_A[747] * mat_B[376] +
//             mat_A[748] * mat_B[408] +
//             mat_A[749] * mat_B[440] +
//             mat_A[750] * mat_B[472] +
//             mat_A[751] * mat_B[504] +
//             mat_A[752] * mat_B[536] +
//             mat_A[753] * mat_B[568] +
//             mat_A[754] * mat_B[600] +
//             mat_A[755] * mat_B[632] +
//             mat_A[756] * mat_B[664] +
//             mat_A[757] * mat_B[696] +
//             mat_A[758] * mat_B[728] +
//             mat_A[759] * mat_B[760] +
//             mat_A[760] * mat_B[792] +
//             mat_A[761] * mat_B[824] +
//             mat_A[762] * mat_B[856] +
//             mat_A[763] * mat_B[888] +
//             mat_A[764] * mat_B[920] +
//             mat_A[765] * mat_B[952] +
//             mat_A[766] * mat_B[984] +
//             mat_A[767] * mat_B[1016];
//  mat_C[761] <= 
//             mat_A[736] * mat_B[25] +
//             mat_A[737] * mat_B[57] +
//             mat_A[738] * mat_B[89] +
//             mat_A[739] * mat_B[121] +
//             mat_A[740] * mat_B[153] +
//             mat_A[741] * mat_B[185] +
//             mat_A[742] * mat_B[217] +
//             mat_A[743] * mat_B[249] +
//             mat_A[744] * mat_B[281] +
//             mat_A[745] * mat_B[313] +
//             mat_A[746] * mat_B[345] +
//             mat_A[747] * mat_B[377] +
//             mat_A[748] * mat_B[409] +
//             mat_A[749] * mat_B[441] +
//             mat_A[750] * mat_B[473] +
//             mat_A[751] * mat_B[505] +
//             mat_A[752] * mat_B[537] +
//             mat_A[753] * mat_B[569] +
//             mat_A[754] * mat_B[601] +
//             mat_A[755] * mat_B[633] +
//             mat_A[756] * mat_B[665] +
//             mat_A[757] * mat_B[697] +
//             mat_A[758] * mat_B[729] +
//             mat_A[759] * mat_B[761] +
//             mat_A[760] * mat_B[793] +
//             mat_A[761] * mat_B[825] +
//             mat_A[762] * mat_B[857] +
//             mat_A[763] * mat_B[889] +
//             mat_A[764] * mat_B[921] +
//             mat_A[765] * mat_B[953] +
//             mat_A[766] * mat_B[985] +
//             mat_A[767] * mat_B[1017];
//  mat_C[762] <= 
//             mat_A[736] * mat_B[26] +
//             mat_A[737] * mat_B[58] +
//             mat_A[738] * mat_B[90] +
//             mat_A[739] * mat_B[122] +
//             mat_A[740] * mat_B[154] +
//             mat_A[741] * mat_B[186] +
//             mat_A[742] * mat_B[218] +
//             mat_A[743] * mat_B[250] +
//             mat_A[744] * mat_B[282] +
//             mat_A[745] * mat_B[314] +
//             mat_A[746] * mat_B[346] +
//             mat_A[747] * mat_B[378] +
//             mat_A[748] * mat_B[410] +
//             mat_A[749] * mat_B[442] +
//             mat_A[750] * mat_B[474] +
//             mat_A[751] * mat_B[506] +
//             mat_A[752] * mat_B[538] +
//             mat_A[753] * mat_B[570] +
//             mat_A[754] * mat_B[602] +
//             mat_A[755] * mat_B[634] +
//             mat_A[756] * mat_B[666] +
//             mat_A[757] * mat_B[698] +
//             mat_A[758] * mat_B[730] +
//             mat_A[759] * mat_B[762] +
//             mat_A[760] * mat_B[794] +
//             mat_A[761] * mat_B[826] +
//             mat_A[762] * mat_B[858] +
//             mat_A[763] * mat_B[890] +
//             mat_A[764] * mat_B[922] +
//             mat_A[765] * mat_B[954] +
//             mat_A[766] * mat_B[986] +
//             mat_A[767] * mat_B[1018];
//  mat_C[763] <= 
//             mat_A[736] * mat_B[27] +
//             mat_A[737] * mat_B[59] +
//             mat_A[738] * mat_B[91] +
//             mat_A[739] * mat_B[123] +
//             mat_A[740] * mat_B[155] +
//             mat_A[741] * mat_B[187] +
//             mat_A[742] * mat_B[219] +
//             mat_A[743] * mat_B[251] +
//             mat_A[744] * mat_B[283] +
//             mat_A[745] * mat_B[315] +
//             mat_A[746] * mat_B[347] +
//             mat_A[747] * mat_B[379] +
//             mat_A[748] * mat_B[411] +
//             mat_A[749] * mat_B[443] +
//             mat_A[750] * mat_B[475] +
//             mat_A[751] * mat_B[507] +
//             mat_A[752] * mat_B[539] +
//             mat_A[753] * mat_B[571] +
//             mat_A[754] * mat_B[603] +
//             mat_A[755] * mat_B[635] +
//             mat_A[756] * mat_B[667] +
//             mat_A[757] * mat_B[699] +
//             mat_A[758] * mat_B[731] +
//             mat_A[759] * mat_B[763] +
//             mat_A[760] * mat_B[795] +
//             mat_A[761] * mat_B[827] +
//             mat_A[762] * mat_B[859] +
//             mat_A[763] * mat_B[891] +
//             mat_A[764] * mat_B[923] +
//             mat_A[765] * mat_B[955] +
//             mat_A[766] * mat_B[987] +
//             mat_A[767] * mat_B[1019];
//  mat_C[764] <= 
//             mat_A[736] * mat_B[28] +
//             mat_A[737] * mat_B[60] +
//             mat_A[738] * mat_B[92] +
//             mat_A[739] * mat_B[124] +
//             mat_A[740] * mat_B[156] +
//             mat_A[741] * mat_B[188] +
//             mat_A[742] * mat_B[220] +
//             mat_A[743] * mat_B[252] +
//             mat_A[744] * mat_B[284] +
//             mat_A[745] * mat_B[316] +
//             mat_A[746] * mat_B[348] +
//             mat_A[747] * mat_B[380] +
//             mat_A[748] * mat_B[412] +
//             mat_A[749] * mat_B[444] +
//             mat_A[750] * mat_B[476] +
//             mat_A[751] * mat_B[508] +
//             mat_A[752] * mat_B[540] +
//             mat_A[753] * mat_B[572] +
//             mat_A[754] * mat_B[604] +
//             mat_A[755] * mat_B[636] +
//             mat_A[756] * mat_B[668] +
//             mat_A[757] * mat_B[700] +
//             mat_A[758] * mat_B[732] +
//             mat_A[759] * mat_B[764] +
//             mat_A[760] * mat_B[796] +
//             mat_A[761] * mat_B[828] +
//             mat_A[762] * mat_B[860] +
//             mat_A[763] * mat_B[892] +
//             mat_A[764] * mat_B[924] +
//             mat_A[765] * mat_B[956] +
//             mat_A[766] * mat_B[988] +
//             mat_A[767] * mat_B[1020];
//  mat_C[765] <= 
//             mat_A[736] * mat_B[29] +
//             mat_A[737] * mat_B[61] +
//             mat_A[738] * mat_B[93] +
//             mat_A[739] * mat_B[125] +
//             mat_A[740] * mat_B[157] +
//             mat_A[741] * mat_B[189] +
//             mat_A[742] * mat_B[221] +
//             mat_A[743] * mat_B[253] +
//             mat_A[744] * mat_B[285] +
//             mat_A[745] * mat_B[317] +
//             mat_A[746] * mat_B[349] +
//             mat_A[747] * mat_B[381] +
//             mat_A[748] * mat_B[413] +
//             mat_A[749] * mat_B[445] +
//             mat_A[750] * mat_B[477] +
//             mat_A[751] * mat_B[509] +
//             mat_A[752] * mat_B[541] +
//             mat_A[753] * mat_B[573] +
//             mat_A[754] * mat_B[605] +
//             mat_A[755] * mat_B[637] +
//             mat_A[756] * mat_B[669] +
//             mat_A[757] * mat_B[701] +
//             mat_A[758] * mat_B[733] +
//             mat_A[759] * mat_B[765] +
//             mat_A[760] * mat_B[797] +
//             mat_A[761] * mat_B[829] +
//             mat_A[762] * mat_B[861] +
//             mat_A[763] * mat_B[893] +
//             mat_A[764] * mat_B[925] +
//             mat_A[765] * mat_B[957] +
//             mat_A[766] * mat_B[989] +
//             mat_A[767] * mat_B[1021];
//  mat_C[766] <= 
//             mat_A[736] * mat_B[30] +
//             mat_A[737] * mat_B[62] +
//             mat_A[738] * mat_B[94] +
//             mat_A[739] * mat_B[126] +
//             mat_A[740] * mat_B[158] +
//             mat_A[741] * mat_B[190] +
//             mat_A[742] * mat_B[222] +
//             mat_A[743] * mat_B[254] +
//             mat_A[744] * mat_B[286] +
//             mat_A[745] * mat_B[318] +
//             mat_A[746] * mat_B[350] +
//             mat_A[747] * mat_B[382] +
//             mat_A[748] * mat_B[414] +
//             mat_A[749] * mat_B[446] +
//             mat_A[750] * mat_B[478] +
//             mat_A[751] * mat_B[510] +
//             mat_A[752] * mat_B[542] +
//             mat_A[753] * mat_B[574] +
//             mat_A[754] * mat_B[606] +
//             mat_A[755] * mat_B[638] +
//             mat_A[756] * mat_B[670] +
//             mat_A[757] * mat_B[702] +
//             mat_A[758] * mat_B[734] +
//             mat_A[759] * mat_B[766] +
//             mat_A[760] * mat_B[798] +
//             mat_A[761] * mat_B[830] +
//             mat_A[762] * mat_B[862] +
//             mat_A[763] * mat_B[894] +
//             mat_A[764] * mat_B[926] +
//             mat_A[765] * mat_B[958] +
//             mat_A[766] * mat_B[990] +
//             mat_A[767] * mat_B[1022];
//  mat_C[767] <= 
//             mat_A[736] * mat_B[31] +
//             mat_A[737] * mat_B[63] +
//             mat_A[738] * mat_B[95] +
//             mat_A[739] * mat_B[127] +
//             mat_A[740] * mat_B[159] +
//             mat_A[741] * mat_B[191] +
//             mat_A[742] * mat_B[223] +
//             mat_A[743] * mat_B[255] +
//             mat_A[744] * mat_B[287] +
//             mat_A[745] * mat_B[319] +
//             mat_A[746] * mat_B[351] +
//             mat_A[747] * mat_B[383] +
//             mat_A[748] * mat_B[415] +
//             mat_A[749] * mat_B[447] +
//             mat_A[750] * mat_B[479] +
//             mat_A[751] * mat_B[511] +
//             mat_A[752] * mat_B[543] +
//             mat_A[753] * mat_B[575] +
//             mat_A[754] * mat_B[607] +
//             mat_A[755] * mat_B[639] +
//             mat_A[756] * mat_B[671] +
//             mat_A[757] * mat_B[703] +
//             mat_A[758] * mat_B[735] +
//             mat_A[759] * mat_B[767] +
//             mat_A[760] * mat_B[799] +
//             mat_A[761] * mat_B[831] +
//             mat_A[762] * mat_B[863] +
//             mat_A[763] * mat_B[895] +
//             mat_A[764] * mat_B[927] +
//             mat_A[765] * mat_B[959] +
//             mat_A[766] * mat_B[991] +
//             mat_A[767] * mat_B[1023];
//  mat_C[768] <= 
//             mat_A[768] * mat_B[0] +
//             mat_A[769] * mat_B[32] +
//             mat_A[770] * mat_B[64] +
//             mat_A[771] * mat_B[96] +
//             mat_A[772] * mat_B[128] +
//             mat_A[773] * mat_B[160] +
//             mat_A[774] * mat_B[192] +
//             mat_A[775] * mat_B[224] +
//             mat_A[776] * mat_B[256] +
//             mat_A[777] * mat_B[288] +
//             mat_A[778] * mat_B[320] +
//             mat_A[779] * mat_B[352] +
//             mat_A[780] * mat_B[384] +
//             mat_A[781] * mat_B[416] +
//             mat_A[782] * mat_B[448] +
//             mat_A[783] * mat_B[480] +
//             mat_A[784] * mat_B[512] +
//             mat_A[785] * mat_B[544] +
//             mat_A[786] * mat_B[576] +
//             mat_A[787] * mat_B[608] +
//             mat_A[788] * mat_B[640] +
//             mat_A[789] * mat_B[672] +
//             mat_A[790] * mat_B[704] +
//             mat_A[791] * mat_B[736] +
//             mat_A[792] * mat_B[768] +
//             mat_A[793] * mat_B[800] +
//             mat_A[794] * mat_B[832] +
//             mat_A[795] * mat_B[864] +
//             mat_A[796] * mat_B[896] +
//             mat_A[797] * mat_B[928] +
//             mat_A[798] * mat_B[960] +
//             mat_A[799] * mat_B[992];
//  mat_C[769] <= 
//             mat_A[768] * mat_B[1] +
//             mat_A[769] * mat_B[33] +
//             mat_A[770] * mat_B[65] +
//             mat_A[771] * mat_B[97] +
//             mat_A[772] * mat_B[129] +
//             mat_A[773] * mat_B[161] +
//             mat_A[774] * mat_B[193] +
//             mat_A[775] * mat_B[225] +
//             mat_A[776] * mat_B[257] +
//             mat_A[777] * mat_B[289] +
//             mat_A[778] * mat_B[321] +
//             mat_A[779] * mat_B[353] +
//             mat_A[780] * mat_B[385] +
//             mat_A[781] * mat_B[417] +
//             mat_A[782] * mat_B[449] +
//             mat_A[783] * mat_B[481] +
//             mat_A[784] * mat_B[513] +
//             mat_A[785] * mat_B[545] +
//             mat_A[786] * mat_B[577] +
//             mat_A[787] * mat_B[609] +
//             mat_A[788] * mat_B[641] +
//             mat_A[789] * mat_B[673] +
//             mat_A[790] * mat_B[705] +
//             mat_A[791] * mat_B[737] +
//             mat_A[792] * mat_B[769] +
//             mat_A[793] * mat_B[801] +
//             mat_A[794] * mat_B[833] +
//             mat_A[795] * mat_B[865] +
//             mat_A[796] * mat_B[897] +
//             mat_A[797] * mat_B[929] +
//             mat_A[798] * mat_B[961] +
//             mat_A[799] * mat_B[993];
//  mat_C[770] <= 
//             mat_A[768] * mat_B[2] +
//             mat_A[769] * mat_B[34] +
//             mat_A[770] * mat_B[66] +
//             mat_A[771] * mat_B[98] +
//             mat_A[772] * mat_B[130] +
//             mat_A[773] * mat_B[162] +
//             mat_A[774] * mat_B[194] +
//             mat_A[775] * mat_B[226] +
//             mat_A[776] * mat_B[258] +
//             mat_A[777] * mat_B[290] +
//             mat_A[778] * mat_B[322] +
//             mat_A[779] * mat_B[354] +
//             mat_A[780] * mat_B[386] +
//             mat_A[781] * mat_B[418] +
//             mat_A[782] * mat_B[450] +
//             mat_A[783] * mat_B[482] +
//             mat_A[784] * mat_B[514] +
//             mat_A[785] * mat_B[546] +
//             mat_A[786] * mat_B[578] +
//             mat_A[787] * mat_B[610] +
//             mat_A[788] * mat_B[642] +
//             mat_A[789] * mat_B[674] +
//             mat_A[790] * mat_B[706] +
//             mat_A[791] * mat_B[738] +
//             mat_A[792] * mat_B[770] +
//             mat_A[793] * mat_B[802] +
//             mat_A[794] * mat_B[834] +
//             mat_A[795] * mat_B[866] +
//             mat_A[796] * mat_B[898] +
//             mat_A[797] * mat_B[930] +
//             mat_A[798] * mat_B[962] +
//             mat_A[799] * mat_B[994];
//  mat_C[771] <= 
//             mat_A[768] * mat_B[3] +
//             mat_A[769] * mat_B[35] +
//             mat_A[770] * mat_B[67] +
//             mat_A[771] * mat_B[99] +
//             mat_A[772] * mat_B[131] +
//             mat_A[773] * mat_B[163] +
//             mat_A[774] * mat_B[195] +
//             mat_A[775] * mat_B[227] +
//             mat_A[776] * mat_B[259] +
//             mat_A[777] * mat_B[291] +
//             mat_A[778] * mat_B[323] +
//             mat_A[779] * mat_B[355] +
//             mat_A[780] * mat_B[387] +
//             mat_A[781] * mat_B[419] +
//             mat_A[782] * mat_B[451] +
//             mat_A[783] * mat_B[483] +
//             mat_A[784] * mat_B[515] +
//             mat_A[785] * mat_B[547] +
//             mat_A[786] * mat_B[579] +
//             mat_A[787] * mat_B[611] +
//             mat_A[788] * mat_B[643] +
//             mat_A[789] * mat_B[675] +
//             mat_A[790] * mat_B[707] +
//             mat_A[791] * mat_B[739] +
//             mat_A[792] * mat_B[771] +
//             mat_A[793] * mat_B[803] +
//             mat_A[794] * mat_B[835] +
//             mat_A[795] * mat_B[867] +
//             mat_A[796] * mat_B[899] +
//             mat_A[797] * mat_B[931] +
//             mat_A[798] * mat_B[963] +
//             mat_A[799] * mat_B[995];
//  mat_C[772] <= 
//             mat_A[768] * mat_B[4] +
//             mat_A[769] * mat_B[36] +
//             mat_A[770] * mat_B[68] +
//             mat_A[771] * mat_B[100] +
//             mat_A[772] * mat_B[132] +
//             mat_A[773] * mat_B[164] +
//             mat_A[774] * mat_B[196] +
//             mat_A[775] * mat_B[228] +
//             mat_A[776] * mat_B[260] +
//             mat_A[777] * mat_B[292] +
//             mat_A[778] * mat_B[324] +
//             mat_A[779] * mat_B[356] +
//             mat_A[780] * mat_B[388] +
//             mat_A[781] * mat_B[420] +
//             mat_A[782] * mat_B[452] +
//             mat_A[783] * mat_B[484] +
//             mat_A[784] * mat_B[516] +
//             mat_A[785] * mat_B[548] +
//             mat_A[786] * mat_B[580] +
//             mat_A[787] * mat_B[612] +
//             mat_A[788] * mat_B[644] +
//             mat_A[789] * mat_B[676] +
//             mat_A[790] * mat_B[708] +
//             mat_A[791] * mat_B[740] +
//             mat_A[792] * mat_B[772] +
//             mat_A[793] * mat_B[804] +
//             mat_A[794] * mat_B[836] +
//             mat_A[795] * mat_B[868] +
//             mat_A[796] * mat_B[900] +
//             mat_A[797] * mat_B[932] +
//             mat_A[798] * mat_B[964] +
//             mat_A[799] * mat_B[996];
//  mat_C[773] <= 
//             mat_A[768] * mat_B[5] +
//             mat_A[769] * mat_B[37] +
//             mat_A[770] * mat_B[69] +
//             mat_A[771] * mat_B[101] +
//             mat_A[772] * mat_B[133] +
//             mat_A[773] * mat_B[165] +
//             mat_A[774] * mat_B[197] +
//             mat_A[775] * mat_B[229] +
//             mat_A[776] * mat_B[261] +
//             mat_A[777] * mat_B[293] +
//             mat_A[778] * mat_B[325] +
//             mat_A[779] * mat_B[357] +
//             mat_A[780] * mat_B[389] +
//             mat_A[781] * mat_B[421] +
//             mat_A[782] * mat_B[453] +
//             mat_A[783] * mat_B[485] +
//             mat_A[784] * mat_B[517] +
//             mat_A[785] * mat_B[549] +
//             mat_A[786] * mat_B[581] +
//             mat_A[787] * mat_B[613] +
//             mat_A[788] * mat_B[645] +
//             mat_A[789] * mat_B[677] +
//             mat_A[790] * mat_B[709] +
//             mat_A[791] * mat_B[741] +
//             mat_A[792] * mat_B[773] +
//             mat_A[793] * mat_B[805] +
//             mat_A[794] * mat_B[837] +
//             mat_A[795] * mat_B[869] +
//             mat_A[796] * mat_B[901] +
//             mat_A[797] * mat_B[933] +
//             mat_A[798] * mat_B[965] +
//             mat_A[799] * mat_B[997];
//  mat_C[774] <= 
//             mat_A[768] * mat_B[6] +
//             mat_A[769] * mat_B[38] +
//             mat_A[770] * mat_B[70] +
//             mat_A[771] * mat_B[102] +
//             mat_A[772] * mat_B[134] +
//             mat_A[773] * mat_B[166] +
//             mat_A[774] * mat_B[198] +
//             mat_A[775] * mat_B[230] +
//             mat_A[776] * mat_B[262] +
//             mat_A[777] * mat_B[294] +
//             mat_A[778] * mat_B[326] +
//             mat_A[779] * mat_B[358] +
//             mat_A[780] * mat_B[390] +
//             mat_A[781] * mat_B[422] +
//             mat_A[782] * mat_B[454] +
//             mat_A[783] * mat_B[486] +
//             mat_A[784] * mat_B[518] +
//             mat_A[785] * mat_B[550] +
//             mat_A[786] * mat_B[582] +
//             mat_A[787] * mat_B[614] +
//             mat_A[788] * mat_B[646] +
//             mat_A[789] * mat_B[678] +
//             mat_A[790] * mat_B[710] +
//             mat_A[791] * mat_B[742] +
//             mat_A[792] * mat_B[774] +
//             mat_A[793] * mat_B[806] +
//             mat_A[794] * mat_B[838] +
//             mat_A[795] * mat_B[870] +
//             mat_A[796] * mat_B[902] +
//             mat_A[797] * mat_B[934] +
//             mat_A[798] * mat_B[966] +
//             mat_A[799] * mat_B[998];
//  mat_C[775] <= 
//             mat_A[768] * mat_B[7] +
//             mat_A[769] * mat_B[39] +
//             mat_A[770] * mat_B[71] +
//             mat_A[771] * mat_B[103] +
//             mat_A[772] * mat_B[135] +
//             mat_A[773] * mat_B[167] +
//             mat_A[774] * mat_B[199] +
//             mat_A[775] * mat_B[231] +
//             mat_A[776] * mat_B[263] +
//             mat_A[777] * mat_B[295] +
//             mat_A[778] * mat_B[327] +
//             mat_A[779] * mat_B[359] +
//             mat_A[780] * mat_B[391] +
//             mat_A[781] * mat_B[423] +
//             mat_A[782] * mat_B[455] +
//             mat_A[783] * mat_B[487] +
//             mat_A[784] * mat_B[519] +
//             mat_A[785] * mat_B[551] +
//             mat_A[786] * mat_B[583] +
//             mat_A[787] * mat_B[615] +
//             mat_A[788] * mat_B[647] +
//             mat_A[789] * mat_B[679] +
//             mat_A[790] * mat_B[711] +
//             mat_A[791] * mat_B[743] +
//             mat_A[792] * mat_B[775] +
//             mat_A[793] * mat_B[807] +
//             mat_A[794] * mat_B[839] +
//             mat_A[795] * mat_B[871] +
//             mat_A[796] * mat_B[903] +
//             mat_A[797] * mat_B[935] +
//             mat_A[798] * mat_B[967] +
//             mat_A[799] * mat_B[999];
//  mat_C[776] <= 
//             mat_A[768] * mat_B[8] +
//             mat_A[769] * mat_B[40] +
//             mat_A[770] * mat_B[72] +
//             mat_A[771] * mat_B[104] +
//             mat_A[772] * mat_B[136] +
//             mat_A[773] * mat_B[168] +
//             mat_A[774] * mat_B[200] +
//             mat_A[775] * mat_B[232] +
//             mat_A[776] * mat_B[264] +
//             mat_A[777] * mat_B[296] +
//             mat_A[778] * mat_B[328] +
//             mat_A[779] * mat_B[360] +
//             mat_A[780] * mat_B[392] +
//             mat_A[781] * mat_B[424] +
//             mat_A[782] * mat_B[456] +
//             mat_A[783] * mat_B[488] +
//             mat_A[784] * mat_B[520] +
//             mat_A[785] * mat_B[552] +
//             mat_A[786] * mat_B[584] +
//             mat_A[787] * mat_B[616] +
//             mat_A[788] * mat_B[648] +
//             mat_A[789] * mat_B[680] +
//             mat_A[790] * mat_B[712] +
//             mat_A[791] * mat_B[744] +
//             mat_A[792] * mat_B[776] +
//             mat_A[793] * mat_B[808] +
//             mat_A[794] * mat_B[840] +
//             mat_A[795] * mat_B[872] +
//             mat_A[796] * mat_B[904] +
//             mat_A[797] * mat_B[936] +
//             mat_A[798] * mat_B[968] +
//             mat_A[799] * mat_B[1000];
//  mat_C[777] <= 
//             mat_A[768] * mat_B[9] +
//             mat_A[769] * mat_B[41] +
//             mat_A[770] * mat_B[73] +
//             mat_A[771] * mat_B[105] +
//             mat_A[772] * mat_B[137] +
//             mat_A[773] * mat_B[169] +
//             mat_A[774] * mat_B[201] +
//             mat_A[775] * mat_B[233] +
//             mat_A[776] * mat_B[265] +
//             mat_A[777] * mat_B[297] +
//             mat_A[778] * mat_B[329] +
//             mat_A[779] * mat_B[361] +
//             mat_A[780] * mat_B[393] +
//             mat_A[781] * mat_B[425] +
//             mat_A[782] * mat_B[457] +
//             mat_A[783] * mat_B[489] +
//             mat_A[784] * mat_B[521] +
//             mat_A[785] * mat_B[553] +
//             mat_A[786] * mat_B[585] +
//             mat_A[787] * mat_B[617] +
//             mat_A[788] * mat_B[649] +
//             mat_A[789] * mat_B[681] +
//             mat_A[790] * mat_B[713] +
//             mat_A[791] * mat_B[745] +
//             mat_A[792] * mat_B[777] +
//             mat_A[793] * mat_B[809] +
//             mat_A[794] * mat_B[841] +
//             mat_A[795] * mat_B[873] +
//             mat_A[796] * mat_B[905] +
//             mat_A[797] * mat_B[937] +
//             mat_A[798] * mat_B[969] +
//             mat_A[799] * mat_B[1001];
//  mat_C[778] <= 
//             mat_A[768] * mat_B[10] +
//             mat_A[769] * mat_B[42] +
//             mat_A[770] * mat_B[74] +
//             mat_A[771] * mat_B[106] +
//             mat_A[772] * mat_B[138] +
//             mat_A[773] * mat_B[170] +
//             mat_A[774] * mat_B[202] +
//             mat_A[775] * mat_B[234] +
//             mat_A[776] * mat_B[266] +
//             mat_A[777] * mat_B[298] +
//             mat_A[778] * mat_B[330] +
//             mat_A[779] * mat_B[362] +
//             mat_A[780] * mat_B[394] +
//             mat_A[781] * mat_B[426] +
//             mat_A[782] * mat_B[458] +
//             mat_A[783] * mat_B[490] +
//             mat_A[784] * mat_B[522] +
//             mat_A[785] * mat_B[554] +
//             mat_A[786] * mat_B[586] +
//             mat_A[787] * mat_B[618] +
//             mat_A[788] * mat_B[650] +
//             mat_A[789] * mat_B[682] +
//             mat_A[790] * mat_B[714] +
//             mat_A[791] * mat_B[746] +
//             mat_A[792] * mat_B[778] +
//             mat_A[793] * mat_B[810] +
//             mat_A[794] * mat_B[842] +
//             mat_A[795] * mat_B[874] +
//             mat_A[796] * mat_B[906] +
//             mat_A[797] * mat_B[938] +
//             mat_A[798] * mat_B[970] +
//             mat_A[799] * mat_B[1002];
//  mat_C[779] <= 
//             mat_A[768] * mat_B[11] +
//             mat_A[769] * mat_B[43] +
//             mat_A[770] * mat_B[75] +
//             mat_A[771] * mat_B[107] +
//             mat_A[772] * mat_B[139] +
//             mat_A[773] * mat_B[171] +
//             mat_A[774] * mat_B[203] +
//             mat_A[775] * mat_B[235] +
//             mat_A[776] * mat_B[267] +
//             mat_A[777] * mat_B[299] +
//             mat_A[778] * mat_B[331] +
//             mat_A[779] * mat_B[363] +
//             mat_A[780] * mat_B[395] +
//             mat_A[781] * mat_B[427] +
//             mat_A[782] * mat_B[459] +
//             mat_A[783] * mat_B[491] +
//             mat_A[784] * mat_B[523] +
//             mat_A[785] * mat_B[555] +
//             mat_A[786] * mat_B[587] +
//             mat_A[787] * mat_B[619] +
//             mat_A[788] * mat_B[651] +
//             mat_A[789] * mat_B[683] +
//             mat_A[790] * mat_B[715] +
//             mat_A[791] * mat_B[747] +
//             mat_A[792] * mat_B[779] +
//             mat_A[793] * mat_B[811] +
//             mat_A[794] * mat_B[843] +
//             mat_A[795] * mat_B[875] +
//             mat_A[796] * mat_B[907] +
//             mat_A[797] * mat_B[939] +
//             mat_A[798] * mat_B[971] +
//             mat_A[799] * mat_B[1003];
//  mat_C[780] <= 
//             mat_A[768] * mat_B[12] +
//             mat_A[769] * mat_B[44] +
//             mat_A[770] * mat_B[76] +
//             mat_A[771] * mat_B[108] +
//             mat_A[772] * mat_B[140] +
//             mat_A[773] * mat_B[172] +
//             mat_A[774] * mat_B[204] +
//             mat_A[775] * mat_B[236] +
//             mat_A[776] * mat_B[268] +
//             mat_A[777] * mat_B[300] +
//             mat_A[778] * mat_B[332] +
//             mat_A[779] * mat_B[364] +
//             mat_A[780] * mat_B[396] +
//             mat_A[781] * mat_B[428] +
//             mat_A[782] * mat_B[460] +
//             mat_A[783] * mat_B[492] +
//             mat_A[784] * mat_B[524] +
//             mat_A[785] * mat_B[556] +
//             mat_A[786] * mat_B[588] +
//             mat_A[787] * mat_B[620] +
//             mat_A[788] * mat_B[652] +
//             mat_A[789] * mat_B[684] +
//             mat_A[790] * mat_B[716] +
//             mat_A[791] * mat_B[748] +
//             mat_A[792] * mat_B[780] +
//             mat_A[793] * mat_B[812] +
//             mat_A[794] * mat_B[844] +
//             mat_A[795] * mat_B[876] +
//             mat_A[796] * mat_B[908] +
//             mat_A[797] * mat_B[940] +
//             mat_A[798] * mat_B[972] +
//             mat_A[799] * mat_B[1004];
//  mat_C[781] <= 
//             mat_A[768] * mat_B[13] +
//             mat_A[769] * mat_B[45] +
//             mat_A[770] * mat_B[77] +
//             mat_A[771] * mat_B[109] +
//             mat_A[772] * mat_B[141] +
//             mat_A[773] * mat_B[173] +
//             mat_A[774] * mat_B[205] +
//             mat_A[775] * mat_B[237] +
//             mat_A[776] * mat_B[269] +
//             mat_A[777] * mat_B[301] +
//             mat_A[778] * mat_B[333] +
//             mat_A[779] * mat_B[365] +
//             mat_A[780] * mat_B[397] +
//             mat_A[781] * mat_B[429] +
//             mat_A[782] * mat_B[461] +
//             mat_A[783] * mat_B[493] +
//             mat_A[784] * mat_B[525] +
//             mat_A[785] * mat_B[557] +
//             mat_A[786] * mat_B[589] +
//             mat_A[787] * mat_B[621] +
//             mat_A[788] * mat_B[653] +
//             mat_A[789] * mat_B[685] +
//             mat_A[790] * mat_B[717] +
//             mat_A[791] * mat_B[749] +
//             mat_A[792] * mat_B[781] +
//             mat_A[793] * mat_B[813] +
//             mat_A[794] * mat_B[845] +
//             mat_A[795] * mat_B[877] +
//             mat_A[796] * mat_B[909] +
//             mat_A[797] * mat_B[941] +
//             mat_A[798] * mat_B[973] +
//             mat_A[799] * mat_B[1005];
//  mat_C[782] <= 
//             mat_A[768] * mat_B[14] +
//             mat_A[769] * mat_B[46] +
//             mat_A[770] * mat_B[78] +
//             mat_A[771] * mat_B[110] +
//             mat_A[772] * mat_B[142] +
//             mat_A[773] * mat_B[174] +
//             mat_A[774] * mat_B[206] +
//             mat_A[775] * mat_B[238] +
//             mat_A[776] * mat_B[270] +
//             mat_A[777] * mat_B[302] +
//             mat_A[778] * mat_B[334] +
//             mat_A[779] * mat_B[366] +
//             mat_A[780] * mat_B[398] +
//             mat_A[781] * mat_B[430] +
//             mat_A[782] * mat_B[462] +
//             mat_A[783] * mat_B[494] +
//             mat_A[784] * mat_B[526] +
//             mat_A[785] * mat_B[558] +
//             mat_A[786] * mat_B[590] +
//             mat_A[787] * mat_B[622] +
//             mat_A[788] * mat_B[654] +
//             mat_A[789] * mat_B[686] +
//             mat_A[790] * mat_B[718] +
//             mat_A[791] * mat_B[750] +
//             mat_A[792] * mat_B[782] +
//             mat_A[793] * mat_B[814] +
//             mat_A[794] * mat_B[846] +
//             mat_A[795] * mat_B[878] +
//             mat_A[796] * mat_B[910] +
//             mat_A[797] * mat_B[942] +
//             mat_A[798] * mat_B[974] +
//             mat_A[799] * mat_B[1006];
//  mat_C[783] <= 
//             mat_A[768] * mat_B[15] +
//             mat_A[769] * mat_B[47] +
//             mat_A[770] * mat_B[79] +
//             mat_A[771] * mat_B[111] +
//             mat_A[772] * mat_B[143] +
//             mat_A[773] * mat_B[175] +
//             mat_A[774] * mat_B[207] +
//             mat_A[775] * mat_B[239] +
//             mat_A[776] * mat_B[271] +
//             mat_A[777] * mat_B[303] +
//             mat_A[778] * mat_B[335] +
//             mat_A[779] * mat_B[367] +
//             mat_A[780] * mat_B[399] +
//             mat_A[781] * mat_B[431] +
//             mat_A[782] * mat_B[463] +
//             mat_A[783] * mat_B[495] +
//             mat_A[784] * mat_B[527] +
//             mat_A[785] * mat_B[559] +
//             mat_A[786] * mat_B[591] +
//             mat_A[787] * mat_B[623] +
//             mat_A[788] * mat_B[655] +
//             mat_A[789] * mat_B[687] +
//             mat_A[790] * mat_B[719] +
//             mat_A[791] * mat_B[751] +
//             mat_A[792] * mat_B[783] +
//             mat_A[793] * mat_B[815] +
//             mat_A[794] * mat_B[847] +
//             mat_A[795] * mat_B[879] +
//             mat_A[796] * mat_B[911] +
//             mat_A[797] * mat_B[943] +
//             mat_A[798] * mat_B[975] +
//             mat_A[799] * mat_B[1007];
//  mat_C[784] <= 
//             mat_A[768] * mat_B[16] +
//             mat_A[769] * mat_B[48] +
//             mat_A[770] * mat_B[80] +
//             mat_A[771] * mat_B[112] +
//             mat_A[772] * mat_B[144] +
//             mat_A[773] * mat_B[176] +
//             mat_A[774] * mat_B[208] +
//             mat_A[775] * mat_B[240] +
//             mat_A[776] * mat_B[272] +
//             mat_A[777] * mat_B[304] +
//             mat_A[778] * mat_B[336] +
//             mat_A[779] * mat_B[368] +
//             mat_A[780] * mat_B[400] +
//             mat_A[781] * mat_B[432] +
//             mat_A[782] * mat_B[464] +
//             mat_A[783] * mat_B[496] +
//             mat_A[784] * mat_B[528] +
//             mat_A[785] * mat_B[560] +
//             mat_A[786] * mat_B[592] +
//             mat_A[787] * mat_B[624] +
//             mat_A[788] * mat_B[656] +
//             mat_A[789] * mat_B[688] +
//             mat_A[790] * mat_B[720] +
//             mat_A[791] * mat_B[752] +
//             mat_A[792] * mat_B[784] +
//             mat_A[793] * mat_B[816] +
//             mat_A[794] * mat_B[848] +
//             mat_A[795] * mat_B[880] +
//             mat_A[796] * mat_B[912] +
//             mat_A[797] * mat_B[944] +
//             mat_A[798] * mat_B[976] +
//             mat_A[799] * mat_B[1008];
//  mat_C[785] <= 
//             mat_A[768] * mat_B[17] +
//             mat_A[769] * mat_B[49] +
//             mat_A[770] * mat_B[81] +
//             mat_A[771] * mat_B[113] +
//             mat_A[772] * mat_B[145] +
//             mat_A[773] * mat_B[177] +
//             mat_A[774] * mat_B[209] +
//             mat_A[775] * mat_B[241] +
//             mat_A[776] * mat_B[273] +
//             mat_A[777] * mat_B[305] +
//             mat_A[778] * mat_B[337] +
//             mat_A[779] * mat_B[369] +
//             mat_A[780] * mat_B[401] +
//             mat_A[781] * mat_B[433] +
//             mat_A[782] * mat_B[465] +
//             mat_A[783] * mat_B[497] +
//             mat_A[784] * mat_B[529] +
//             mat_A[785] * mat_B[561] +
//             mat_A[786] * mat_B[593] +
//             mat_A[787] * mat_B[625] +
//             mat_A[788] * mat_B[657] +
//             mat_A[789] * mat_B[689] +
//             mat_A[790] * mat_B[721] +
//             mat_A[791] * mat_B[753] +
//             mat_A[792] * mat_B[785] +
//             mat_A[793] * mat_B[817] +
//             mat_A[794] * mat_B[849] +
//             mat_A[795] * mat_B[881] +
//             mat_A[796] * mat_B[913] +
//             mat_A[797] * mat_B[945] +
//             mat_A[798] * mat_B[977] +
//             mat_A[799] * mat_B[1009];
//  mat_C[786] <= 
//             mat_A[768] * mat_B[18] +
//             mat_A[769] * mat_B[50] +
//             mat_A[770] * mat_B[82] +
//             mat_A[771] * mat_B[114] +
//             mat_A[772] * mat_B[146] +
//             mat_A[773] * mat_B[178] +
//             mat_A[774] * mat_B[210] +
//             mat_A[775] * mat_B[242] +
//             mat_A[776] * mat_B[274] +
//             mat_A[777] * mat_B[306] +
//             mat_A[778] * mat_B[338] +
//             mat_A[779] * mat_B[370] +
//             mat_A[780] * mat_B[402] +
//             mat_A[781] * mat_B[434] +
//             mat_A[782] * mat_B[466] +
//             mat_A[783] * mat_B[498] +
//             mat_A[784] * mat_B[530] +
//             mat_A[785] * mat_B[562] +
//             mat_A[786] * mat_B[594] +
//             mat_A[787] * mat_B[626] +
//             mat_A[788] * mat_B[658] +
//             mat_A[789] * mat_B[690] +
//             mat_A[790] * mat_B[722] +
//             mat_A[791] * mat_B[754] +
//             mat_A[792] * mat_B[786] +
//             mat_A[793] * mat_B[818] +
//             mat_A[794] * mat_B[850] +
//             mat_A[795] * mat_B[882] +
//             mat_A[796] * mat_B[914] +
//             mat_A[797] * mat_B[946] +
//             mat_A[798] * mat_B[978] +
//             mat_A[799] * mat_B[1010];
//  mat_C[787] <= 
//             mat_A[768] * mat_B[19] +
//             mat_A[769] * mat_B[51] +
//             mat_A[770] * mat_B[83] +
//             mat_A[771] * mat_B[115] +
//             mat_A[772] * mat_B[147] +
//             mat_A[773] * mat_B[179] +
//             mat_A[774] * mat_B[211] +
//             mat_A[775] * mat_B[243] +
//             mat_A[776] * mat_B[275] +
//             mat_A[777] * mat_B[307] +
//             mat_A[778] * mat_B[339] +
//             mat_A[779] * mat_B[371] +
//             mat_A[780] * mat_B[403] +
//             mat_A[781] * mat_B[435] +
//             mat_A[782] * mat_B[467] +
//             mat_A[783] * mat_B[499] +
//             mat_A[784] * mat_B[531] +
//             mat_A[785] * mat_B[563] +
//             mat_A[786] * mat_B[595] +
//             mat_A[787] * mat_B[627] +
//             mat_A[788] * mat_B[659] +
//             mat_A[789] * mat_B[691] +
//             mat_A[790] * mat_B[723] +
//             mat_A[791] * mat_B[755] +
//             mat_A[792] * mat_B[787] +
//             mat_A[793] * mat_B[819] +
//             mat_A[794] * mat_B[851] +
//             mat_A[795] * mat_B[883] +
//             mat_A[796] * mat_B[915] +
//             mat_A[797] * mat_B[947] +
//             mat_A[798] * mat_B[979] +
//             mat_A[799] * mat_B[1011];
//  mat_C[788] <= 
//             mat_A[768] * mat_B[20] +
//             mat_A[769] * mat_B[52] +
//             mat_A[770] * mat_B[84] +
//             mat_A[771] * mat_B[116] +
//             mat_A[772] * mat_B[148] +
//             mat_A[773] * mat_B[180] +
//             mat_A[774] * mat_B[212] +
//             mat_A[775] * mat_B[244] +
//             mat_A[776] * mat_B[276] +
//             mat_A[777] * mat_B[308] +
//             mat_A[778] * mat_B[340] +
//             mat_A[779] * mat_B[372] +
//             mat_A[780] * mat_B[404] +
//             mat_A[781] * mat_B[436] +
//             mat_A[782] * mat_B[468] +
//             mat_A[783] * mat_B[500] +
//             mat_A[784] * mat_B[532] +
//             mat_A[785] * mat_B[564] +
//             mat_A[786] * mat_B[596] +
//             mat_A[787] * mat_B[628] +
//             mat_A[788] * mat_B[660] +
//             mat_A[789] * mat_B[692] +
//             mat_A[790] * mat_B[724] +
//             mat_A[791] * mat_B[756] +
//             mat_A[792] * mat_B[788] +
//             mat_A[793] * mat_B[820] +
//             mat_A[794] * mat_B[852] +
//             mat_A[795] * mat_B[884] +
//             mat_A[796] * mat_B[916] +
//             mat_A[797] * mat_B[948] +
//             mat_A[798] * mat_B[980] +
//             mat_A[799] * mat_B[1012];
//  mat_C[789] <= 
//             mat_A[768] * mat_B[21] +
//             mat_A[769] * mat_B[53] +
//             mat_A[770] * mat_B[85] +
//             mat_A[771] * mat_B[117] +
//             mat_A[772] * mat_B[149] +
//             mat_A[773] * mat_B[181] +
//             mat_A[774] * mat_B[213] +
//             mat_A[775] * mat_B[245] +
//             mat_A[776] * mat_B[277] +
//             mat_A[777] * mat_B[309] +
//             mat_A[778] * mat_B[341] +
//             mat_A[779] * mat_B[373] +
//             mat_A[780] * mat_B[405] +
//             mat_A[781] * mat_B[437] +
//             mat_A[782] * mat_B[469] +
//             mat_A[783] * mat_B[501] +
//             mat_A[784] * mat_B[533] +
//             mat_A[785] * mat_B[565] +
//             mat_A[786] * mat_B[597] +
//             mat_A[787] * mat_B[629] +
//             mat_A[788] * mat_B[661] +
//             mat_A[789] * mat_B[693] +
//             mat_A[790] * mat_B[725] +
//             mat_A[791] * mat_B[757] +
//             mat_A[792] * mat_B[789] +
//             mat_A[793] * mat_B[821] +
//             mat_A[794] * mat_B[853] +
//             mat_A[795] * mat_B[885] +
//             mat_A[796] * mat_B[917] +
//             mat_A[797] * mat_B[949] +
//             mat_A[798] * mat_B[981] +
//             mat_A[799] * mat_B[1013];
//  mat_C[790] <= 
//             mat_A[768] * mat_B[22] +
//             mat_A[769] * mat_B[54] +
//             mat_A[770] * mat_B[86] +
//             mat_A[771] * mat_B[118] +
//             mat_A[772] * mat_B[150] +
//             mat_A[773] * mat_B[182] +
//             mat_A[774] * mat_B[214] +
//             mat_A[775] * mat_B[246] +
//             mat_A[776] * mat_B[278] +
//             mat_A[777] * mat_B[310] +
//             mat_A[778] * mat_B[342] +
//             mat_A[779] * mat_B[374] +
//             mat_A[780] * mat_B[406] +
//             mat_A[781] * mat_B[438] +
//             mat_A[782] * mat_B[470] +
//             mat_A[783] * mat_B[502] +
//             mat_A[784] * mat_B[534] +
//             mat_A[785] * mat_B[566] +
//             mat_A[786] * mat_B[598] +
//             mat_A[787] * mat_B[630] +
//             mat_A[788] * mat_B[662] +
//             mat_A[789] * mat_B[694] +
//             mat_A[790] * mat_B[726] +
//             mat_A[791] * mat_B[758] +
//             mat_A[792] * mat_B[790] +
//             mat_A[793] * mat_B[822] +
//             mat_A[794] * mat_B[854] +
//             mat_A[795] * mat_B[886] +
//             mat_A[796] * mat_B[918] +
//             mat_A[797] * mat_B[950] +
//             mat_A[798] * mat_B[982] +
//             mat_A[799] * mat_B[1014];
//  mat_C[791] <= 
//             mat_A[768] * mat_B[23] +
//             mat_A[769] * mat_B[55] +
//             mat_A[770] * mat_B[87] +
//             mat_A[771] * mat_B[119] +
//             mat_A[772] * mat_B[151] +
//             mat_A[773] * mat_B[183] +
//             mat_A[774] * mat_B[215] +
//             mat_A[775] * mat_B[247] +
//             mat_A[776] * mat_B[279] +
//             mat_A[777] * mat_B[311] +
//             mat_A[778] * mat_B[343] +
//             mat_A[779] * mat_B[375] +
//             mat_A[780] * mat_B[407] +
//             mat_A[781] * mat_B[439] +
//             mat_A[782] * mat_B[471] +
//             mat_A[783] * mat_B[503] +
//             mat_A[784] * mat_B[535] +
//             mat_A[785] * mat_B[567] +
//             mat_A[786] * mat_B[599] +
//             mat_A[787] * mat_B[631] +
//             mat_A[788] * mat_B[663] +
//             mat_A[789] * mat_B[695] +
//             mat_A[790] * mat_B[727] +
//             mat_A[791] * mat_B[759] +
//             mat_A[792] * mat_B[791] +
//             mat_A[793] * mat_B[823] +
//             mat_A[794] * mat_B[855] +
//             mat_A[795] * mat_B[887] +
//             mat_A[796] * mat_B[919] +
//             mat_A[797] * mat_B[951] +
//             mat_A[798] * mat_B[983] +
//             mat_A[799] * mat_B[1015];
//  mat_C[792] <= 
//             mat_A[768] * mat_B[24] +
//             mat_A[769] * mat_B[56] +
//             mat_A[770] * mat_B[88] +
//             mat_A[771] * mat_B[120] +
//             mat_A[772] * mat_B[152] +
//             mat_A[773] * mat_B[184] +
//             mat_A[774] * mat_B[216] +
//             mat_A[775] * mat_B[248] +
//             mat_A[776] * mat_B[280] +
//             mat_A[777] * mat_B[312] +
//             mat_A[778] * mat_B[344] +
//             mat_A[779] * mat_B[376] +
//             mat_A[780] * mat_B[408] +
//             mat_A[781] * mat_B[440] +
//             mat_A[782] * mat_B[472] +
//             mat_A[783] * mat_B[504] +
//             mat_A[784] * mat_B[536] +
//             mat_A[785] * mat_B[568] +
//             mat_A[786] * mat_B[600] +
//             mat_A[787] * mat_B[632] +
//             mat_A[788] * mat_B[664] +
//             mat_A[789] * mat_B[696] +
//             mat_A[790] * mat_B[728] +
//             mat_A[791] * mat_B[760] +
//             mat_A[792] * mat_B[792] +
//             mat_A[793] * mat_B[824] +
//             mat_A[794] * mat_B[856] +
//             mat_A[795] * mat_B[888] +
//             mat_A[796] * mat_B[920] +
//             mat_A[797] * mat_B[952] +
//             mat_A[798] * mat_B[984] +
//             mat_A[799] * mat_B[1016];
//  mat_C[793] <= 
//             mat_A[768] * mat_B[25] +
//             mat_A[769] * mat_B[57] +
//             mat_A[770] * mat_B[89] +
//             mat_A[771] * mat_B[121] +
//             mat_A[772] * mat_B[153] +
//             mat_A[773] * mat_B[185] +
//             mat_A[774] * mat_B[217] +
//             mat_A[775] * mat_B[249] +
//             mat_A[776] * mat_B[281] +
//             mat_A[777] * mat_B[313] +
//             mat_A[778] * mat_B[345] +
//             mat_A[779] * mat_B[377] +
//             mat_A[780] * mat_B[409] +
//             mat_A[781] * mat_B[441] +
//             mat_A[782] * mat_B[473] +
//             mat_A[783] * mat_B[505] +
//             mat_A[784] * mat_B[537] +
//             mat_A[785] * mat_B[569] +
//             mat_A[786] * mat_B[601] +
//             mat_A[787] * mat_B[633] +
//             mat_A[788] * mat_B[665] +
//             mat_A[789] * mat_B[697] +
//             mat_A[790] * mat_B[729] +
//             mat_A[791] * mat_B[761] +
//             mat_A[792] * mat_B[793] +
//             mat_A[793] * mat_B[825] +
//             mat_A[794] * mat_B[857] +
//             mat_A[795] * mat_B[889] +
//             mat_A[796] * mat_B[921] +
//             mat_A[797] * mat_B[953] +
//             mat_A[798] * mat_B[985] +
//             mat_A[799] * mat_B[1017];
//  mat_C[794] <= 
//             mat_A[768] * mat_B[26] +
//             mat_A[769] * mat_B[58] +
//             mat_A[770] * mat_B[90] +
//             mat_A[771] * mat_B[122] +
//             mat_A[772] * mat_B[154] +
//             mat_A[773] * mat_B[186] +
//             mat_A[774] * mat_B[218] +
//             mat_A[775] * mat_B[250] +
//             mat_A[776] * mat_B[282] +
//             mat_A[777] * mat_B[314] +
//             mat_A[778] * mat_B[346] +
//             mat_A[779] * mat_B[378] +
//             mat_A[780] * mat_B[410] +
//             mat_A[781] * mat_B[442] +
//             mat_A[782] * mat_B[474] +
//             mat_A[783] * mat_B[506] +
//             mat_A[784] * mat_B[538] +
//             mat_A[785] * mat_B[570] +
//             mat_A[786] * mat_B[602] +
//             mat_A[787] * mat_B[634] +
//             mat_A[788] * mat_B[666] +
//             mat_A[789] * mat_B[698] +
//             mat_A[790] * mat_B[730] +
//             mat_A[791] * mat_B[762] +
//             mat_A[792] * mat_B[794] +
//             mat_A[793] * mat_B[826] +
//             mat_A[794] * mat_B[858] +
//             mat_A[795] * mat_B[890] +
//             mat_A[796] * mat_B[922] +
//             mat_A[797] * mat_B[954] +
//             mat_A[798] * mat_B[986] +
//             mat_A[799] * mat_B[1018];
//  mat_C[795] <= 
//             mat_A[768] * mat_B[27] +
//             mat_A[769] * mat_B[59] +
//             mat_A[770] * mat_B[91] +
//             mat_A[771] * mat_B[123] +
//             mat_A[772] * mat_B[155] +
//             mat_A[773] * mat_B[187] +
//             mat_A[774] * mat_B[219] +
//             mat_A[775] * mat_B[251] +
//             mat_A[776] * mat_B[283] +
//             mat_A[777] * mat_B[315] +
//             mat_A[778] * mat_B[347] +
//             mat_A[779] * mat_B[379] +
//             mat_A[780] * mat_B[411] +
//             mat_A[781] * mat_B[443] +
//             mat_A[782] * mat_B[475] +
//             mat_A[783] * mat_B[507] +
//             mat_A[784] * mat_B[539] +
//             mat_A[785] * mat_B[571] +
//             mat_A[786] * mat_B[603] +
//             mat_A[787] * mat_B[635] +
//             mat_A[788] * mat_B[667] +
//             mat_A[789] * mat_B[699] +
//             mat_A[790] * mat_B[731] +
//             mat_A[791] * mat_B[763] +
//             mat_A[792] * mat_B[795] +
//             mat_A[793] * mat_B[827] +
//             mat_A[794] * mat_B[859] +
//             mat_A[795] * mat_B[891] +
//             mat_A[796] * mat_B[923] +
//             mat_A[797] * mat_B[955] +
//             mat_A[798] * mat_B[987] +
//             mat_A[799] * mat_B[1019];
//  mat_C[796] <= 
//             mat_A[768] * mat_B[28] +
//             mat_A[769] * mat_B[60] +
//             mat_A[770] * mat_B[92] +
//             mat_A[771] * mat_B[124] +
//             mat_A[772] * mat_B[156] +
//             mat_A[773] * mat_B[188] +
//             mat_A[774] * mat_B[220] +
//             mat_A[775] * mat_B[252] +
//             mat_A[776] * mat_B[284] +
//             mat_A[777] * mat_B[316] +
//             mat_A[778] * mat_B[348] +
//             mat_A[779] * mat_B[380] +
//             mat_A[780] * mat_B[412] +
//             mat_A[781] * mat_B[444] +
//             mat_A[782] * mat_B[476] +
//             mat_A[783] * mat_B[508] +
//             mat_A[784] * mat_B[540] +
//             mat_A[785] * mat_B[572] +
//             mat_A[786] * mat_B[604] +
//             mat_A[787] * mat_B[636] +
//             mat_A[788] * mat_B[668] +
//             mat_A[789] * mat_B[700] +
//             mat_A[790] * mat_B[732] +
//             mat_A[791] * mat_B[764] +
//             mat_A[792] * mat_B[796] +
//             mat_A[793] * mat_B[828] +
//             mat_A[794] * mat_B[860] +
//             mat_A[795] * mat_B[892] +
//             mat_A[796] * mat_B[924] +
//             mat_A[797] * mat_B[956] +
//             mat_A[798] * mat_B[988] +
//             mat_A[799] * mat_B[1020];
//  mat_C[797] <= 
//             mat_A[768] * mat_B[29] +
//             mat_A[769] * mat_B[61] +
//             mat_A[770] * mat_B[93] +
//             mat_A[771] * mat_B[125] +
//             mat_A[772] * mat_B[157] +
//             mat_A[773] * mat_B[189] +
//             mat_A[774] * mat_B[221] +
//             mat_A[775] * mat_B[253] +
//             mat_A[776] * mat_B[285] +
//             mat_A[777] * mat_B[317] +
//             mat_A[778] * mat_B[349] +
//             mat_A[779] * mat_B[381] +
//             mat_A[780] * mat_B[413] +
//             mat_A[781] * mat_B[445] +
//             mat_A[782] * mat_B[477] +
//             mat_A[783] * mat_B[509] +
//             mat_A[784] * mat_B[541] +
//             mat_A[785] * mat_B[573] +
//             mat_A[786] * mat_B[605] +
//             mat_A[787] * mat_B[637] +
//             mat_A[788] * mat_B[669] +
//             mat_A[789] * mat_B[701] +
//             mat_A[790] * mat_B[733] +
//             mat_A[791] * mat_B[765] +
//             mat_A[792] * mat_B[797] +
//             mat_A[793] * mat_B[829] +
//             mat_A[794] * mat_B[861] +
//             mat_A[795] * mat_B[893] +
//             mat_A[796] * mat_B[925] +
//             mat_A[797] * mat_B[957] +
//             mat_A[798] * mat_B[989] +
//             mat_A[799] * mat_B[1021];
//  mat_C[798] <= 
//             mat_A[768] * mat_B[30] +
//             mat_A[769] * mat_B[62] +
//             mat_A[770] * mat_B[94] +
//             mat_A[771] * mat_B[126] +
//             mat_A[772] * mat_B[158] +
//             mat_A[773] * mat_B[190] +
//             mat_A[774] * mat_B[222] +
//             mat_A[775] * mat_B[254] +
//             mat_A[776] * mat_B[286] +
//             mat_A[777] * mat_B[318] +
//             mat_A[778] * mat_B[350] +
//             mat_A[779] * mat_B[382] +
//             mat_A[780] * mat_B[414] +
//             mat_A[781] * mat_B[446] +
//             mat_A[782] * mat_B[478] +
//             mat_A[783] * mat_B[510] +
//             mat_A[784] * mat_B[542] +
//             mat_A[785] * mat_B[574] +
//             mat_A[786] * mat_B[606] +
//             mat_A[787] * mat_B[638] +
//             mat_A[788] * mat_B[670] +
//             mat_A[789] * mat_B[702] +
//             mat_A[790] * mat_B[734] +
//             mat_A[791] * mat_B[766] +
//             mat_A[792] * mat_B[798] +
//             mat_A[793] * mat_B[830] +
//             mat_A[794] * mat_B[862] +
//             mat_A[795] * mat_B[894] +
//             mat_A[796] * mat_B[926] +
//             mat_A[797] * mat_B[958] +
//             mat_A[798] * mat_B[990] +
//             mat_A[799] * mat_B[1022];
//  mat_C[799] <= 
//             mat_A[768] * mat_B[31] +
//             mat_A[769] * mat_B[63] +
//             mat_A[770] * mat_B[95] +
//             mat_A[771] * mat_B[127] +
//             mat_A[772] * mat_B[159] +
//             mat_A[773] * mat_B[191] +
//             mat_A[774] * mat_B[223] +
//             mat_A[775] * mat_B[255] +
//             mat_A[776] * mat_B[287] +
//             mat_A[777] * mat_B[319] +
//             mat_A[778] * mat_B[351] +
//             mat_A[779] * mat_B[383] +
//             mat_A[780] * mat_B[415] +
//             mat_A[781] * mat_B[447] +
//             mat_A[782] * mat_B[479] +
//             mat_A[783] * mat_B[511] +
//             mat_A[784] * mat_B[543] +
//             mat_A[785] * mat_B[575] +
//             mat_A[786] * mat_B[607] +
//             mat_A[787] * mat_B[639] +
//             mat_A[788] * mat_B[671] +
//             mat_A[789] * mat_B[703] +
//             mat_A[790] * mat_B[735] +
//             mat_A[791] * mat_B[767] +
//             mat_A[792] * mat_B[799] +
//             mat_A[793] * mat_B[831] +
//             mat_A[794] * mat_B[863] +
//             mat_A[795] * mat_B[895] +
//             mat_A[796] * mat_B[927] +
//             mat_A[797] * mat_B[959] +
//             mat_A[798] * mat_B[991] +
//             mat_A[799] * mat_B[1023];
//  mat_C[800] <= 
//             mat_A[800] * mat_B[0] +
//             mat_A[801] * mat_B[32] +
//             mat_A[802] * mat_B[64] +
//             mat_A[803] * mat_B[96] +
//             mat_A[804] * mat_B[128] +
//             mat_A[805] * mat_B[160] +
//             mat_A[806] * mat_B[192] +
//             mat_A[807] * mat_B[224] +
//             mat_A[808] * mat_B[256] +
//             mat_A[809] * mat_B[288] +
//             mat_A[810] * mat_B[320] +
//             mat_A[811] * mat_B[352] +
//             mat_A[812] * mat_B[384] +
//             mat_A[813] * mat_B[416] +
//             mat_A[814] * mat_B[448] +
//             mat_A[815] * mat_B[480] +
//             mat_A[816] * mat_B[512] +
//             mat_A[817] * mat_B[544] +
//             mat_A[818] * mat_B[576] +
//             mat_A[819] * mat_B[608] +
//             mat_A[820] * mat_B[640] +
//             mat_A[821] * mat_B[672] +
//             mat_A[822] * mat_B[704] +
//             mat_A[823] * mat_B[736] +
//             mat_A[824] * mat_B[768] +
//             mat_A[825] * mat_B[800] +
//             mat_A[826] * mat_B[832] +
//             mat_A[827] * mat_B[864] +
//             mat_A[828] * mat_B[896] +
//             mat_A[829] * mat_B[928] +
//             mat_A[830] * mat_B[960] +
//             mat_A[831] * mat_B[992];
//  mat_C[801] <= 
//             mat_A[800] * mat_B[1] +
//             mat_A[801] * mat_B[33] +
//             mat_A[802] * mat_B[65] +
//             mat_A[803] * mat_B[97] +
//             mat_A[804] * mat_B[129] +
//             mat_A[805] * mat_B[161] +
//             mat_A[806] * mat_B[193] +
//             mat_A[807] * mat_B[225] +
//             mat_A[808] * mat_B[257] +
//             mat_A[809] * mat_B[289] +
//             mat_A[810] * mat_B[321] +
//             mat_A[811] * mat_B[353] +
//             mat_A[812] * mat_B[385] +
//             mat_A[813] * mat_B[417] +
//             mat_A[814] * mat_B[449] +
//             mat_A[815] * mat_B[481] +
//             mat_A[816] * mat_B[513] +
//             mat_A[817] * mat_B[545] +
//             mat_A[818] * mat_B[577] +
//             mat_A[819] * mat_B[609] +
//             mat_A[820] * mat_B[641] +
//             mat_A[821] * mat_B[673] +
//             mat_A[822] * mat_B[705] +
//             mat_A[823] * mat_B[737] +
//             mat_A[824] * mat_B[769] +
//             mat_A[825] * mat_B[801] +
//             mat_A[826] * mat_B[833] +
//             mat_A[827] * mat_B[865] +
//             mat_A[828] * mat_B[897] +
//             mat_A[829] * mat_B[929] +
//             mat_A[830] * mat_B[961] +
//             mat_A[831] * mat_B[993];
//  mat_C[802] <= 
//             mat_A[800] * mat_B[2] +
//             mat_A[801] * mat_B[34] +
//             mat_A[802] * mat_B[66] +
//             mat_A[803] * mat_B[98] +
//             mat_A[804] * mat_B[130] +
//             mat_A[805] * mat_B[162] +
//             mat_A[806] * mat_B[194] +
//             mat_A[807] * mat_B[226] +
//             mat_A[808] * mat_B[258] +
//             mat_A[809] * mat_B[290] +
//             mat_A[810] * mat_B[322] +
//             mat_A[811] * mat_B[354] +
//             mat_A[812] * mat_B[386] +
//             mat_A[813] * mat_B[418] +
//             mat_A[814] * mat_B[450] +
//             mat_A[815] * mat_B[482] +
//             mat_A[816] * mat_B[514] +
//             mat_A[817] * mat_B[546] +
//             mat_A[818] * mat_B[578] +
//             mat_A[819] * mat_B[610] +
//             mat_A[820] * mat_B[642] +
//             mat_A[821] * mat_B[674] +
//             mat_A[822] * mat_B[706] +
//             mat_A[823] * mat_B[738] +
//             mat_A[824] * mat_B[770] +
//             mat_A[825] * mat_B[802] +
//             mat_A[826] * mat_B[834] +
//             mat_A[827] * mat_B[866] +
//             mat_A[828] * mat_B[898] +
//             mat_A[829] * mat_B[930] +
//             mat_A[830] * mat_B[962] +
//             mat_A[831] * mat_B[994];
//  mat_C[803] <= 
//             mat_A[800] * mat_B[3] +
//             mat_A[801] * mat_B[35] +
//             mat_A[802] * mat_B[67] +
//             mat_A[803] * mat_B[99] +
//             mat_A[804] * mat_B[131] +
//             mat_A[805] * mat_B[163] +
//             mat_A[806] * mat_B[195] +
//             mat_A[807] * mat_B[227] +
//             mat_A[808] * mat_B[259] +
//             mat_A[809] * mat_B[291] +
//             mat_A[810] * mat_B[323] +
//             mat_A[811] * mat_B[355] +
//             mat_A[812] * mat_B[387] +
//             mat_A[813] * mat_B[419] +
//             mat_A[814] * mat_B[451] +
//             mat_A[815] * mat_B[483] +
//             mat_A[816] * mat_B[515] +
//             mat_A[817] * mat_B[547] +
//             mat_A[818] * mat_B[579] +
//             mat_A[819] * mat_B[611] +
//             mat_A[820] * mat_B[643] +
//             mat_A[821] * mat_B[675] +
//             mat_A[822] * mat_B[707] +
//             mat_A[823] * mat_B[739] +
//             mat_A[824] * mat_B[771] +
//             mat_A[825] * mat_B[803] +
//             mat_A[826] * mat_B[835] +
//             mat_A[827] * mat_B[867] +
//             mat_A[828] * mat_B[899] +
//             mat_A[829] * mat_B[931] +
//             mat_A[830] * mat_B[963] +
//             mat_A[831] * mat_B[995];
//  mat_C[804] <= 
//             mat_A[800] * mat_B[4] +
//             mat_A[801] * mat_B[36] +
//             mat_A[802] * mat_B[68] +
//             mat_A[803] * mat_B[100] +
//             mat_A[804] * mat_B[132] +
//             mat_A[805] * mat_B[164] +
//             mat_A[806] * mat_B[196] +
//             mat_A[807] * mat_B[228] +
//             mat_A[808] * mat_B[260] +
//             mat_A[809] * mat_B[292] +
//             mat_A[810] * mat_B[324] +
//             mat_A[811] * mat_B[356] +
//             mat_A[812] * mat_B[388] +
//             mat_A[813] * mat_B[420] +
//             mat_A[814] * mat_B[452] +
//             mat_A[815] * mat_B[484] +
//             mat_A[816] * mat_B[516] +
//             mat_A[817] * mat_B[548] +
//             mat_A[818] * mat_B[580] +
//             mat_A[819] * mat_B[612] +
//             mat_A[820] * mat_B[644] +
//             mat_A[821] * mat_B[676] +
//             mat_A[822] * mat_B[708] +
//             mat_A[823] * mat_B[740] +
//             mat_A[824] * mat_B[772] +
//             mat_A[825] * mat_B[804] +
//             mat_A[826] * mat_B[836] +
//             mat_A[827] * mat_B[868] +
//             mat_A[828] * mat_B[900] +
//             mat_A[829] * mat_B[932] +
//             mat_A[830] * mat_B[964] +
//             mat_A[831] * mat_B[996];
//  mat_C[805] <= 
//             mat_A[800] * mat_B[5] +
//             mat_A[801] * mat_B[37] +
//             mat_A[802] * mat_B[69] +
//             mat_A[803] * mat_B[101] +
//             mat_A[804] * mat_B[133] +
//             mat_A[805] * mat_B[165] +
//             mat_A[806] * mat_B[197] +
//             mat_A[807] * mat_B[229] +
//             mat_A[808] * mat_B[261] +
//             mat_A[809] * mat_B[293] +
//             mat_A[810] * mat_B[325] +
//             mat_A[811] * mat_B[357] +
//             mat_A[812] * mat_B[389] +
//             mat_A[813] * mat_B[421] +
//             mat_A[814] * mat_B[453] +
//             mat_A[815] * mat_B[485] +
//             mat_A[816] * mat_B[517] +
//             mat_A[817] * mat_B[549] +
//             mat_A[818] * mat_B[581] +
//             mat_A[819] * mat_B[613] +
//             mat_A[820] * mat_B[645] +
//             mat_A[821] * mat_B[677] +
//             mat_A[822] * mat_B[709] +
//             mat_A[823] * mat_B[741] +
//             mat_A[824] * mat_B[773] +
//             mat_A[825] * mat_B[805] +
//             mat_A[826] * mat_B[837] +
//             mat_A[827] * mat_B[869] +
//             mat_A[828] * mat_B[901] +
//             mat_A[829] * mat_B[933] +
//             mat_A[830] * mat_B[965] +
//             mat_A[831] * mat_B[997];
//  mat_C[806] <= 
//             mat_A[800] * mat_B[6] +
//             mat_A[801] * mat_B[38] +
//             mat_A[802] * mat_B[70] +
//             mat_A[803] * mat_B[102] +
//             mat_A[804] * mat_B[134] +
//             mat_A[805] * mat_B[166] +
//             mat_A[806] * mat_B[198] +
//             mat_A[807] * mat_B[230] +
//             mat_A[808] * mat_B[262] +
//             mat_A[809] * mat_B[294] +
//             mat_A[810] * mat_B[326] +
//             mat_A[811] * mat_B[358] +
//             mat_A[812] * mat_B[390] +
//             mat_A[813] * mat_B[422] +
//             mat_A[814] * mat_B[454] +
//             mat_A[815] * mat_B[486] +
//             mat_A[816] * mat_B[518] +
//             mat_A[817] * mat_B[550] +
//             mat_A[818] * mat_B[582] +
//             mat_A[819] * mat_B[614] +
//             mat_A[820] * mat_B[646] +
//             mat_A[821] * mat_B[678] +
//             mat_A[822] * mat_B[710] +
//             mat_A[823] * mat_B[742] +
//             mat_A[824] * mat_B[774] +
//             mat_A[825] * mat_B[806] +
//             mat_A[826] * mat_B[838] +
//             mat_A[827] * mat_B[870] +
//             mat_A[828] * mat_B[902] +
//             mat_A[829] * mat_B[934] +
//             mat_A[830] * mat_B[966] +
//             mat_A[831] * mat_B[998];
//  mat_C[807] <= 
//             mat_A[800] * mat_B[7] +
//             mat_A[801] * mat_B[39] +
//             mat_A[802] * mat_B[71] +
//             mat_A[803] * mat_B[103] +
//             mat_A[804] * mat_B[135] +
//             mat_A[805] * mat_B[167] +
//             mat_A[806] * mat_B[199] +
//             mat_A[807] * mat_B[231] +
//             mat_A[808] * mat_B[263] +
//             mat_A[809] * mat_B[295] +
//             mat_A[810] * mat_B[327] +
//             mat_A[811] * mat_B[359] +
//             mat_A[812] * mat_B[391] +
//             mat_A[813] * mat_B[423] +
//             mat_A[814] * mat_B[455] +
//             mat_A[815] * mat_B[487] +
//             mat_A[816] * mat_B[519] +
//             mat_A[817] * mat_B[551] +
//             mat_A[818] * mat_B[583] +
//             mat_A[819] * mat_B[615] +
//             mat_A[820] * mat_B[647] +
//             mat_A[821] * mat_B[679] +
//             mat_A[822] * mat_B[711] +
//             mat_A[823] * mat_B[743] +
//             mat_A[824] * mat_B[775] +
//             mat_A[825] * mat_B[807] +
//             mat_A[826] * mat_B[839] +
//             mat_A[827] * mat_B[871] +
//             mat_A[828] * mat_B[903] +
//             mat_A[829] * mat_B[935] +
//             mat_A[830] * mat_B[967] +
//             mat_A[831] * mat_B[999];
//  mat_C[808] <= 
//             mat_A[800] * mat_B[8] +
//             mat_A[801] * mat_B[40] +
//             mat_A[802] * mat_B[72] +
//             mat_A[803] * mat_B[104] +
//             mat_A[804] * mat_B[136] +
//             mat_A[805] * mat_B[168] +
//             mat_A[806] * mat_B[200] +
//             mat_A[807] * mat_B[232] +
//             mat_A[808] * mat_B[264] +
//             mat_A[809] * mat_B[296] +
//             mat_A[810] * mat_B[328] +
//             mat_A[811] * mat_B[360] +
//             mat_A[812] * mat_B[392] +
//             mat_A[813] * mat_B[424] +
//             mat_A[814] * mat_B[456] +
//             mat_A[815] * mat_B[488] +
//             mat_A[816] * mat_B[520] +
//             mat_A[817] * mat_B[552] +
//             mat_A[818] * mat_B[584] +
//             mat_A[819] * mat_B[616] +
//             mat_A[820] * mat_B[648] +
//             mat_A[821] * mat_B[680] +
//             mat_A[822] * mat_B[712] +
//             mat_A[823] * mat_B[744] +
//             mat_A[824] * mat_B[776] +
//             mat_A[825] * mat_B[808] +
//             mat_A[826] * mat_B[840] +
//             mat_A[827] * mat_B[872] +
//             mat_A[828] * mat_B[904] +
//             mat_A[829] * mat_B[936] +
//             mat_A[830] * mat_B[968] +
//             mat_A[831] * mat_B[1000];
//  mat_C[809] <= 
//             mat_A[800] * mat_B[9] +
//             mat_A[801] * mat_B[41] +
//             mat_A[802] * mat_B[73] +
//             mat_A[803] * mat_B[105] +
//             mat_A[804] * mat_B[137] +
//             mat_A[805] * mat_B[169] +
//             mat_A[806] * mat_B[201] +
//             mat_A[807] * mat_B[233] +
//             mat_A[808] * mat_B[265] +
//             mat_A[809] * mat_B[297] +
//             mat_A[810] * mat_B[329] +
//             mat_A[811] * mat_B[361] +
//             mat_A[812] * mat_B[393] +
//             mat_A[813] * mat_B[425] +
//             mat_A[814] * mat_B[457] +
//             mat_A[815] * mat_B[489] +
//             mat_A[816] * mat_B[521] +
//             mat_A[817] * mat_B[553] +
//             mat_A[818] * mat_B[585] +
//             mat_A[819] * mat_B[617] +
//             mat_A[820] * mat_B[649] +
//             mat_A[821] * mat_B[681] +
//             mat_A[822] * mat_B[713] +
//             mat_A[823] * mat_B[745] +
//             mat_A[824] * mat_B[777] +
//             mat_A[825] * mat_B[809] +
//             mat_A[826] * mat_B[841] +
//             mat_A[827] * mat_B[873] +
//             mat_A[828] * mat_B[905] +
//             mat_A[829] * mat_B[937] +
//             mat_A[830] * mat_B[969] +
//             mat_A[831] * mat_B[1001];
//  mat_C[810] <= 
//             mat_A[800] * mat_B[10] +
//             mat_A[801] * mat_B[42] +
//             mat_A[802] * mat_B[74] +
//             mat_A[803] * mat_B[106] +
//             mat_A[804] * mat_B[138] +
//             mat_A[805] * mat_B[170] +
//             mat_A[806] * mat_B[202] +
//             mat_A[807] * mat_B[234] +
//             mat_A[808] * mat_B[266] +
//             mat_A[809] * mat_B[298] +
//             mat_A[810] * mat_B[330] +
//             mat_A[811] * mat_B[362] +
//             mat_A[812] * mat_B[394] +
//             mat_A[813] * mat_B[426] +
//             mat_A[814] * mat_B[458] +
//             mat_A[815] * mat_B[490] +
//             mat_A[816] * mat_B[522] +
//             mat_A[817] * mat_B[554] +
//             mat_A[818] * mat_B[586] +
//             mat_A[819] * mat_B[618] +
//             mat_A[820] * mat_B[650] +
//             mat_A[821] * mat_B[682] +
//             mat_A[822] * mat_B[714] +
//             mat_A[823] * mat_B[746] +
//             mat_A[824] * mat_B[778] +
//             mat_A[825] * mat_B[810] +
//             mat_A[826] * mat_B[842] +
//             mat_A[827] * mat_B[874] +
//             mat_A[828] * mat_B[906] +
//             mat_A[829] * mat_B[938] +
//             mat_A[830] * mat_B[970] +
//             mat_A[831] * mat_B[1002];
//  mat_C[811] <= 
//             mat_A[800] * mat_B[11] +
//             mat_A[801] * mat_B[43] +
//             mat_A[802] * mat_B[75] +
//             mat_A[803] * mat_B[107] +
//             mat_A[804] * mat_B[139] +
//             mat_A[805] * mat_B[171] +
//             mat_A[806] * mat_B[203] +
//             mat_A[807] * mat_B[235] +
//             mat_A[808] * mat_B[267] +
//             mat_A[809] * mat_B[299] +
//             mat_A[810] * mat_B[331] +
//             mat_A[811] * mat_B[363] +
//             mat_A[812] * mat_B[395] +
//             mat_A[813] * mat_B[427] +
//             mat_A[814] * mat_B[459] +
//             mat_A[815] * mat_B[491] +
//             mat_A[816] * mat_B[523] +
//             mat_A[817] * mat_B[555] +
//             mat_A[818] * mat_B[587] +
//             mat_A[819] * mat_B[619] +
//             mat_A[820] * mat_B[651] +
//             mat_A[821] * mat_B[683] +
//             mat_A[822] * mat_B[715] +
//             mat_A[823] * mat_B[747] +
//             mat_A[824] * mat_B[779] +
//             mat_A[825] * mat_B[811] +
//             mat_A[826] * mat_B[843] +
//             mat_A[827] * mat_B[875] +
//             mat_A[828] * mat_B[907] +
//             mat_A[829] * mat_B[939] +
//             mat_A[830] * mat_B[971] +
//             mat_A[831] * mat_B[1003];
//  mat_C[812] <= 
//             mat_A[800] * mat_B[12] +
//             mat_A[801] * mat_B[44] +
//             mat_A[802] * mat_B[76] +
//             mat_A[803] * mat_B[108] +
//             mat_A[804] * mat_B[140] +
//             mat_A[805] * mat_B[172] +
//             mat_A[806] * mat_B[204] +
//             mat_A[807] * mat_B[236] +
//             mat_A[808] * mat_B[268] +
//             mat_A[809] * mat_B[300] +
//             mat_A[810] * mat_B[332] +
//             mat_A[811] * mat_B[364] +
//             mat_A[812] * mat_B[396] +
//             mat_A[813] * mat_B[428] +
//             mat_A[814] * mat_B[460] +
//             mat_A[815] * mat_B[492] +
//             mat_A[816] * mat_B[524] +
//             mat_A[817] * mat_B[556] +
//             mat_A[818] * mat_B[588] +
//             mat_A[819] * mat_B[620] +
//             mat_A[820] * mat_B[652] +
//             mat_A[821] * mat_B[684] +
//             mat_A[822] * mat_B[716] +
//             mat_A[823] * mat_B[748] +
//             mat_A[824] * mat_B[780] +
//             mat_A[825] * mat_B[812] +
//             mat_A[826] * mat_B[844] +
//             mat_A[827] * mat_B[876] +
//             mat_A[828] * mat_B[908] +
//             mat_A[829] * mat_B[940] +
//             mat_A[830] * mat_B[972] +
//             mat_A[831] * mat_B[1004];
//  mat_C[813] <= 
//             mat_A[800] * mat_B[13] +
//             mat_A[801] * mat_B[45] +
//             mat_A[802] * mat_B[77] +
//             mat_A[803] * mat_B[109] +
//             mat_A[804] * mat_B[141] +
//             mat_A[805] * mat_B[173] +
//             mat_A[806] * mat_B[205] +
//             mat_A[807] * mat_B[237] +
//             mat_A[808] * mat_B[269] +
//             mat_A[809] * mat_B[301] +
//             mat_A[810] * mat_B[333] +
//             mat_A[811] * mat_B[365] +
//             mat_A[812] * mat_B[397] +
//             mat_A[813] * mat_B[429] +
//             mat_A[814] * mat_B[461] +
//             mat_A[815] * mat_B[493] +
//             mat_A[816] * mat_B[525] +
//             mat_A[817] * mat_B[557] +
//             mat_A[818] * mat_B[589] +
//             mat_A[819] * mat_B[621] +
//             mat_A[820] * mat_B[653] +
//             mat_A[821] * mat_B[685] +
//             mat_A[822] * mat_B[717] +
//             mat_A[823] * mat_B[749] +
//             mat_A[824] * mat_B[781] +
//             mat_A[825] * mat_B[813] +
//             mat_A[826] * mat_B[845] +
//             mat_A[827] * mat_B[877] +
//             mat_A[828] * mat_B[909] +
//             mat_A[829] * mat_B[941] +
//             mat_A[830] * mat_B[973] +
//             mat_A[831] * mat_B[1005];
//  mat_C[814] <= 
//             mat_A[800] * mat_B[14] +
//             mat_A[801] * mat_B[46] +
//             mat_A[802] * mat_B[78] +
//             mat_A[803] * mat_B[110] +
//             mat_A[804] * mat_B[142] +
//             mat_A[805] * mat_B[174] +
//             mat_A[806] * mat_B[206] +
//             mat_A[807] * mat_B[238] +
//             mat_A[808] * mat_B[270] +
//             mat_A[809] * mat_B[302] +
//             mat_A[810] * mat_B[334] +
//             mat_A[811] * mat_B[366] +
//             mat_A[812] * mat_B[398] +
//             mat_A[813] * mat_B[430] +
//             mat_A[814] * mat_B[462] +
//             mat_A[815] * mat_B[494] +
//             mat_A[816] * mat_B[526] +
//             mat_A[817] * mat_B[558] +
//             mat_A[818] * mat_B[590] +
//             mat_A[819] * mat_B[622] +
//             mat_A[820] * mat_B[654] +
//             mat_A[821] * mat_B[686] +
//             mat_A[822] * mat_B[718] +
//             mat_A[823] * mat_B[750] +
//             mat_A[824] * mat_B[782] +
//             mat_A[825] * mat_B[814] +
//             mat_A[826] * mat_B[846] +
//             mat_A[827] * mat_B[878] +
//             mat_A[828] * mat_B[910] +
//             mat_A[829] * mat_B[942] +
//             mat_A[830] * mat_B[974] +
//             mat_A[831] * mat_B[1006];
//  mat_C[815] <= 
//             mat_A[800] * mat_B[15] +
//             mat_A[801] * mat_B[47] +
//             mat_A[802] * mat_B[79] +
//             mat_A[803] * mat_B[111] +
//             mat_A[804] * mat_B[143] +
//             mat_A[805] * mat_B[175] +
//             mat_A[806] * mat_B[207] +
//             mat_A[807] * mat_B[239] +
//             mat_A[808] * mat_B[271] +
//             mat_A[809] * mat_B[303] +
//             mat_A[810] * mat_B[335] +
//             mat_A[811] * mat_B[367] +
//             mat_A[812] * mat_B[399] +
//             mat_A[813] * mat_B[431] +
//             mat_A[814] * mat_B[463] +
//             mat_A[815] * mat_B[495] +
//             mat_A[816] * mat_B[527] +
//             mat_A[817] * mat_B[559] +
//             mat_A[818] * mat_B[591] +
//             mat_A[819] * mat_B[623] +
//             mat_A[820] * mat_B[655] +
//             mat_A[821] * mat_B[687] +
//             mat_A[822] * mat_B[719] +
//             mat_A[823] * mat_B[751] +
//             mat_A[824] * mat_B[783] +
//             mat_A[825] * mat_B[815] +
//             mat_A[826] * mat_B[847] +
//             mat_A[827] * mat_B[879] +
//             mat_A[828] * mat_B[911] +
//             mat_A[829] * mat_B[943] +
//             mat_A[830] * mat_B[975] +
//             mat_A[831] * mat_B[1007];
//  mat_C[816] <= 
//             mat_A[800] * mat_B[16] +
//             mat_A[801] * mat_B[48] +
//             mat_A[802] * mat_B[80] +
//             mat_A[803] * mat_B[112] +
//             mat_A[804] * mat_B[144] +
//             mat_A[805] * mat_B[176] +
//             mat_A[806] * mat_B[208] +
//             mat_A[807] * mat_B[240] +
//             mat_A[808] * mat_B[272] +
//             mat_A[809] * mat_B[304] +
//             mat_A[810] * mat_B[336] +
//             mat_A[811] * mat_B[368] +
//             mat_A[812] * mat_B[400] +
//             mat_A[813] * mat_B[432] +
//             mat_A[814] * mat_B[464] +
//             mat_A[815] * mat_B[496] +
//             mat_A[816] * mat_B[528] +
//             mat_A[817] * mat_B[560] +
//             mat_A[818] * mat_B[592] +
//             mat_A[819] * mat_B[624] +
//             mat_A[820] * mat_B[656] +
//             mat_A[821] * mat_B[688] +
//             mat_A[822] * mat_B[720] +
//             mat_A[823] * mat_B[752] +
//             mat_A[824] * mat_B[784] +
//             mat_A[825] * mat_B[816] +
//             mat_A[826] * mat_B[848] +
//             mat_A[827] * mat_B[880] +
//             mat_A[828] * mat_B[912] +
//             mat_A[829] * mat_B[944] +
//             mat_A[830] * mat_B[976] +
//             mat_A[831] * mat_B[1008];
//  mat_C[817] <= 
//             mat_A[800] * mat_B[17] +
//             mat_A[801] * mat_B[49] +
//             mat_A[802] * mat_B[81] +
//             mat_A[803] * mat_B[113] +
//             mat_A[804] * mat_B[145] +
//             mat_A[805] * mat_B[177] +
//             mat_A[806] * mat_B[209] +
//             mat_A[807] * mat_B[241] +
//             mat_A[808] * mat_B[273] +
//             mat_A[809] * mat_B[305] +
//             mat_A[810] * mat_B[337] +
//             mat_A[811] * mat_B[369] +
//             mat_A[812] * mat_B[401] +
//             mat_A[813] * mat_B[433] +
//             mat_A[814] * mat_B[465] +
//             mat_A[815] * mat_B[497] +
//             mat_A[816] * mat_B[529] +
//             mat_A[817] * mat_B[561] +
//             mat_A[818] * mat_B[593] +
//             mat_A[819] * mat_B[625] +
//             mat_A[820] * mat_B[657] +
//             mat_A[821] * mat_B[689] +
//             mat_A[822] * mat_B[721] +
//             mat_A[823] * mat_B[753] +
//             mat_A[824] * mat_B[785] +
//             mat_A[825] * mat_B[817] +
//             mat_A[826] * mat_B[849] +
//             mat_A[827] * mat_B[881] +
//             mat_A[828] * mat_B[913] +
//             mat_A[829] * mat_B[945] +
//             mat_A[830] * mat_B[977] +
//             mat_A[831] * mat_B[1009];
//  mat_C[818] <= 
//             mat_A[800] * mat_B[18] +
//             mat_A[801] * mat_B[50] +
//             mat_A[802] * mat_B[82] +
//             mat_A[803] * mat_B[114] +
//             mat_A[804] * mat_B[146] +
//             mat_A[805] * mat_B[178] +
//             mat_A[806] * mat_B[210] +
//             mat_A[807] * mat_B[242] +
//             mat_A[808] * mat_B[274] +
//             mat_A[809] * mat_B[306] +
//             mat_A[810] * mat_B[338] +
//             mat_A[811] * mat_B[370] +
//             mat_A[812] * mat_B[402] +
//             mat_A[813] * mat_B[434] +
//             mat_A[814] * mat_B[466] +
//             mat_A[815] * mat_B[498] +
//             mat_A[816] * mat_B[530] +
//             mat_A[817] * mat_B[562] +
//             mat_A[818] * mat_B[594] +
//             mat_A[819] * mat_B[626] +
//             mat_A[820] * mat_B[658] +
//             mat_A[821] * mat_B[690] +
//             mat_A[822] * mat_B[722] +
//             mat_A[823] * mat_B[754] +
//             mat_A[824] * mat_B[786] +
//             mat_A[825] * mat_B[818] +
//             mat_A[826] * mat_B[850] +
//             mat_A[827] * mat_B[882] +
//             mat_A[828] * mat_B[914] +
//             mat_A[829] * mat_B[946] +
//             mat_A[830] * mat_B[978] +
//             mat_A[831] * mat_B[1010];
//  mat_C[819] <= 
//             mat_A[800] * mat_B[19] +
//             mat_A[801] * mat_B[51] +
//             mat_A[802] * mat_B[83] +
//             mat_A[803] * mat_B[115] +
//             mat_A[804] * mat_B[147] +
//             mat_A[805] * mat_B[179] +
//             mat_A[806] * mat_B[211] +
//             mat_A[807] * mat_B[243] +
//             mat_A[808] * mat_B[275] +
//             mat_A[809] * mat_B[307] +
//             mat_A[810] * mat_B[339] +
//             mat_A[811] * mat_B[371] +
//             mat_A[812] * mat_B[403] +
//             mat_A[813] * mat_B[435] +
//             mat_A[814] * mat_B[467] +
//             mat_A[815] * mat_B[499] +
//             mat_A[816] * mat_B[531] +
//             mat_A[817] * mat_B[563] +
//             mat_A[818] * mat_B[595] +
//             mat_A[819] * mat_B[627] +
//             mat_A[820] * mat_B[659] +
//             mat_A[821] * mat_B[691] +
//             mat_A[822] * mat_B[723] +
//             mat_A[823] * mat_B[755] +
//             mat_A[824] * mat_B[787] +
//             mat_A[825] * mat_B[819] +
//             mat_A[826] * mat_B[851] +
//             mat_A[827] * mat_B[883] +
//             mat_A[828] * mat_B[915] +
//             mat_A[829] * mat_B[947] +
//             mat_A[830] * mat_B[979] +
//             mat_A[831] * mat_B[1011];
//  mat_C[820] <= 
//             mat_A[800] * mat_B[20] +
//             mat_A[801] * mat_B[52] +
//             mat_A[802] * mat_B[84] +
//             mat_A[803] * mat_B[116] +
//             mat_A[804] * mat_B[148] +
//             mat_A[805] * mat_B[180] +
//             mat_A[806] * mat_B[212] +
//             mat_A[807] * mat_B[244] +
//             mat_A[808] * mat_B[276] +
//             mat_A[809] * mat_B[308] +
//             mat_A[810] * mat_B[340] +
//             mat_A[811] * mat_B[372] +
//             mat_A[812] * mat_B[404] +
//             mat_A[813] * mat_B[436] +
//             mat_A[814] * mat_B[468] +
//             mat_A[815] * mat_B[500] +
//             mat_A[816] * mat_B[532] +
//             mat_A[817] * mat_B[564] +
//             mat_A[818] * mat_B[596] +
//             mat_A[819] * mat_B[628] +
//             mat_A[820] * mat_B[660] +
//             mat_A[821] * mat_B[692] +
//             mat_A[822] * mat_B[724] +
//             mat_A[823] * mat_B[756] +
//             mat_A[824] * mat_B[788] +
//             mat_A[825] * mat_B[820] +
//             mat_A[826] * mat_B[852] +
//             mat_A[827] * mat_B[884] +
//             mat_A[828] * mat_B[916] +
//             mat_A[829] * mat_B[948] +
//             mat_A[830] * mat_B[980] +
//             mat_A[831] * mat_B[1012];
//  mat_C[821] <= 
//             mat_A[800] * mat_B[21] +
//             mat_A[801] * mat_B[53] +
//             mat_A[802] * mat_B[85] +
//             mat_A[803] * mat_B[117] +
//             mat_A[804] * mat_B[149] +
//             mat_A[805] * mat_B[181] +
//             mat_A[806] * mat_B[213] +
//             mat_A[807] * mat_B[245] +
//             mat_A[808] * mat_B[277] +
//             mat_A[809] * mat_B[309] +
//             mat_A[810] * mat_B[341] +
//             mat_A[811] * mat_B[373] +
//             mat_A[812] * mat_B[405] +
//             mat_A[813] * mat_B[437] +
//             mat_A[814] * mat_B[469] +
//             mat_A[815] * mat_B[501] +
//             mat_A[816] * mat_B[533] +
//             mat_A[817] * mat_B[565] +
//             mat_A[818] * mat_B[597] +
//             mat_A[819] * mat_B[629] +
//             mat_A[820] * mat_B[661] +
//             mat_A[821] * mat_B[693] +
//             mat_A[822] * mat_B[725] +
//             mat_A[823] * mat_B[757] +
//             mat_A[824] * mat_B[789] +
//             mat_A[825] * mat_B[821] +
//             mat_A[826] * mat_B[853] +
//             mat_A[827] * mat_B[885] +
//             mat_A[828] * mat_B[917] +
//             mat_A[829] * mat_B[949] +
//             mat_A[830] * mat_B[981] +
//             mat_A[831] * mat_B[1013];
//  mat_C[822] <= 
//             mat_A[800] * mat_B[22] +
//             mat_A[801] * mat_B[54] +
//             mat_A[802] * mat_B[86] +
//             mat_A[803] * mat_B[118] +
//             mat_A[804] * mat_B[150] +
//             mat_A[805] * mat_B[182] +
//             mat_A[806] * mat_B[214] +
//             mat_A[807] * mat_B[246] +
//             mat_A[808] * mat_B[278] +
//             mat_A[809] * mat_B[310] +
//             mat_A[810] * mat_B[342] +
//             mat_A[811] * mat_B[374] +
//             mat_A[812] * mat_B[406] +
//             mat_A[813] * mat_B[438] +
//             mat_A[814] * mat_B[470] +
//             mat_A[815] * mat_B[502] +
//             mat_A[816] * mat_B[534] +
//             mat_A[817] * mat_B[566] +
//             mat_A[818] * mat_B[598] +
//             mat_A[819] * mat_B[630] +
//             mat_A[820] * mat_B[662] +
//             mat_A[821] * mat_B[694] +
//             mat_A[822] * mat_B[726] +
//             mat_A[823] * mat_B[758] +
//             mat_A[824] * mat_B[790] +
//             mat_A[825] * mat_B[822] +
//             mat_A[826] * mat_B[854] +
//             mat_A[827] * mat_B[886] +
//             mat_A[828] * mat_B[918] +
//             mat_A[829] * mat_B[950] +
//             mat_A[830] * mat_B[982] +
//             mat_A[831] * mat_B[1014];
//  mat_C[823] <= 
//             mat_A[800] * mat_B[23] +
//             mat_A[801] * mat_B[55] +
//             mat_A[802] * mat_B[87] +
//             mat_A[803] * mat_B[119] +
//             mat_A[804] * mat_B[151] +
//             mat_A[805] * mat_B[183] +
//             mat_A[806] * mat_B[215] +
//             mat_A[807] * mat_B[247] +
//             mat_A[808] * mat_B[279] +
//             mat_A[809] * mat_B[311] +
//             mat_A[810] * mat_B[343] +
//             mat_A[811] * mat_B[375] +
//             mat_A[812] * mat_B[407] +
//             mat_A[813] * mat_B[439] +
//             mat_A[814] * mat_B[471] +
//             mat_A[815] * mat_B[503] +
//             mat_A[816] * mat_B[535] +
//             mat_A[817] * mat_B[567] +
//             mat_A[818] * mat_B[599] +
//             mat_A[819] * mat_B[631] +
//             mat_A[820] * mat_B[663] +
//             mat_A[821] * mat_B[695] +
//             mat_A[822] * mat_B[727] +
//             mat_A[823] * mat_B[759] +
//             mat_A[824] * mat_B[791] +
//             mat_A[825] * mat_B[823] +
//             mat_A[826] * mat_B[855] +
//             mat_A[827] * mat_B[887] +
//             mat_A[828] * mat_B[919] +
//             mat_A[829] * mat_B[951] +
//             mat_A[830] * mat_B[983] +
//             mat_A[831] * mat_B[1015];
//  mat_C[824] <= 
//             mat_A[800] * mat_B[24] +
//             mat_A[801] * mat_B[56] +
//             mat_A[802] * mat_B[88] +
//             mat_A[803] * mat_B[120] +
//             mat_A[804] * mat_B[152] +
//             mat_A[805] * mat_B[184] +
//             mat_A[806] * mat_B[216] +
//             mat_A[807] * mat_B[248] +
//             mat_A[808] * mat_B[280] +
//             mat_A[809] * mat_B[312] +
//             mat_A[810] * mat_B[344] +
//             mat_A[811] * mat_B[376] +
//             mat_A[812] * mat_B[408] +
//             mat_A[813] * mat_B[440] +
//             mat_A[814] * mat_B[472] +
//             mat_A[815] * mat_B[504] +
//             mat_A[816] * mat_B[536] +
//             mat_A[817] * mat_B[568] +
//             mat_A[818] * mat_B[600] +
//             mat_A[819] * mat_B[632] +
//             mat_A[820] * mat_B[664] +
//             mat_A[821] * mat_B[696] +
//             mat_A[822] * mat_B[728] +
//             mat_A[823] * mat_B[760] +
//             mat_A[824] * mat_B[792] +
//             mat_A[825] * mat_B[824] +
//             mat_A[826] * mat_B[856] +
//             mat_A[827] * mat_B[888] +
//             mat_A[828] * mat_B[920] +
//             mat_A[829] * mat_B[952] +
//             mat_A[830] * mat_B[984] +
//             mat_A[831] * mat_B[1016];
//  mat_C[825] <= 
//             mat_A[800] * mat_B[25] +
//             mat_A[801] * mat_B[57] +
//             mat_A[802] * mat_B[89] +
//             mat_A[803] * mat_B[121] +
//             mat_A[804] * mat_B[153] +
//             mat_A[805] * mat_B[185] +
//             mat_A[806] * mat_B[217] +
//             mat_A[807] * mat_B[249] +
//             mat_A[808] * mat_B[281] +
//             mat_A[809] * mat_B[313] +
//             mat_A[810] * mat_B[345] +
//             mat_A[811] * mat_B[377] +
//             mat_A[812] * mat_B[409] +
//             mat_A[813] * mat_B[441] +
//             mat_A[814] * mat_B[473] +
//             mat_A[815] * mat_B[505] +
//             mat_A[816] * mat_B[537] +
//             mat_A[817] * mat_B[569] +
//             mat_A[818] * mat_B[601] +
//             mat_A[819] * mat_B[633] +
//             mat_A[820] * mat_B[665] +
//             mat_A[821] * mat_B[697] +
//             mat_A[822] * mat_B[729] +
//             mat_A[823] * mat_B[761] +
//             mat_A[824] * mat_B[793] +
//             mat_A[825] * mat_B[825] +
//             mat_A[826] * mat_B[857] +
//             mat_A[827] * mat_B[889] +
//             mat_A[828] * mat_B[921] +
//             mat_A[829] * mat_B[953] +
//             mat_A[830] * mat_B[985] +
//             mat_A[831] * mat_B[1017];
//  mat_C[826] <= 
//             mat_A[800] * mat_B[26] +
//             mat_A[801] * mat_B[58] +
//             mat_A[802] * mat_B[90] +
//             mat_A[803] * mat_B[122] +
//             mat_A[804] * mat_B[154] +
//             mat_A[805] * mat_B[186] +
//             mat_A[806] * mat_B[218] +
//             mat_A[807] * mat_B[250] +
//             mat_A[808] * mat_B[282] +
//             mat_A[809] * mat_B[314] +
//             mat_A[810] * mat_B[346] +
//             mat_A[811] * mat_B[378] +
//             mat_A[812] * mat_B[410] +
//             mat_A[813] * mat_B[442] +
//             mat_A[814] * mat_B[474] +
//             mat_A[815] * mat_B[506] +
//             mat_A[816] * mat_B[538] +
//             mat_A[817] * mat_B[570] +
//             mat_A[818] * mat_B[602] +
//             mat_A[819] * mat_B[634] +
//             mat_A[820] * mat_B[666] +
//             mat_A[821] * mat_B[698] +
//             mat_A[822] * mat_B[730] +
//             mat_A[823] * mat_B[762] +
//             mat_A[824] * mat_B[794] +
//             mat_A[825] * mat_B[826] +
//             mat_A[826] * mat_B[858] +
//             mat_A[827] * mat_B[890] +
//             mat_A[828] * mat_B[922] +
//             mat_A[829] * mat_B[954] +
//             mat_A[830] * mat_B[986] +
//             mat_A[831] * mat_B[1018];
//  mat_C[827] <= 
//             mat_A[800] * mat_B[27] +
//             mat_A[801] * mat_B[59] +
//             mat_A[802] * mat_B[91] +
//             mat_A[803] * mat_B[123] +
//             mat_A[804] * mat_B[155] +
//             mat_A[805] * mat_B[187] +
//             mat_A[806] * mat_B[219] +
//             mat_A[807] * mat_B[251] +
//             mat_A[808] * mat_B[283] +
//             mat_A[809] * mat_B[315] +
//             mat_A[810] * mat_B[347] +
//             mat_A[811] * mat_B[379] +
//             mat_A[812] * mat_B[411] +
//             mat_A[813] * mat_B[443] +
//             mat_A[814] * mat_B[475] +
//             mat_A[815] * mat_B[507] +
//             mat_A[816] * mat_B[539] +
//             mat_A[817] * mat_B[571] +
//             mat_A[818] * mat_B[603] +
//             mat_A[819] * mat_B[635] +
//             mat_A[820] * mat_B[667] +
//             mat_A[821] * mat_B[699] +
//             mat_A[822] * mat_B[731] +
//             mat_A[823] * mat_B[763] +
//             mat_A[824] * mat_B[795] +
//             mat_A[825] * mat_B[827] +
//             mat_A[826] * mat_B[859] +
//             mat_A[827] * mat_B[891] +
//             mat_A[828] * mat_B[923] +
//             mat_A[829] * mat_B[955] +
//             mat_A[830] * mat_B[987] +
//             mat_A[831] * mat_B[1019];
//  mat_C[828] <= 
//             mat_A[800] * mat_B[28] +
//             mat_A[801] * mat_B[60] +
//             mat_A[802] * mat_B[92] +
//             mat_A[803] * mat_B[124] +
//             mat_A[804] * mat_B[156] +
//             mat_A[805] * mat_B[188] +
//             mat_A[806] * mat_B[220] +
//             mat_A[807] * mat_B[252] +
//             mat_A[808] * mat_B[284] +
//             mat_A[809] * mat_B[316] +
//             mat_A[810] * mat_B[348] +
//             mat_A[811] * mat_B[380] +
//             mat_A[812] * mat_B[412] +
//             mat_A[813] * mat_B[444] +
//             mat_A[814] * mat_B[476] +
//             mat_A[815] * mat_B[508] +
//             mat_A[816] * mat_B[540] +
//             mat_A[817] * mat_B[572] +
//             mat_A[818] * mat_B[604] +
//             mat_A[819] * mat_B[636] +
//             mat_A[820] * mat_B[668] +
//             mat_A[821] * mat_B[700] +
//             mat_A[822] * mat_B[732] +
//             mat_A[823] * mat_B[764] +
//             mat_A[824] * mat_B[796] +
//             mat_A[825] * mat_B[828] +
//             mat_A[826] * mat_B[860] +
//             mat_A[827] * mat_B[892] +
//             mat_A[828] * mat_B[924] +
//             mat_A[829] * mat_B[956] +
//             mat_A[830] * mat_B[988] +
//             mat_A[831] * mat_B[1020];
//  mat_C[829] <= 
//             mat_A[800] * mat_B[29] +
//             mat_A[801] * mat_B[61] +
//             mat_A[802] * mat_B[93] +
//             mat_A[803] * mat_B[125] +
//             mat_A[804] * mat_B[157] +
//             mat_A[805] * mat_B[189] +
//             mat_A[806] * mat_B[221] +
//             mat_A[807] * mat_B[253] +
//             mat_A[808] * mat_B[285] +
//             mat_A[809] * mat_B[317] +
//             mat_A[810] * mat_B[349] +
//             mat_A[811] * mat_B[381] +
//             mat_A[812] * mat_B[413] +
//             mat_A[813] * mat_B[445] +
//             mat_A[814] * mat_B[477] +
//             mat_A[815] * mat_B[509] +
//             mat_A[816] * mat_B[541] +
//             mat_A[817] * mat_B[573] +
//             mat_A[818] * mat_B[605] +
//             mat_A[819] * mat_B[637] +
//             mat_A[820] * mat_B[669] +
//             mat_A[821] * mat_B[701] +
//             mat_A[822] * mat_B[733] +
//             mat_A[823] * mat_B[765] +
//             mat_A[824] * mat_B[797] +
//             mat_A[825] * mat_B[829] +
//             mat_A[826] * mat_B[861] +
//             mat_A[827] * mat_B[893] +
//             mat_A[828] * mat_B[925] +
//             mat_A[829] * mat_B[957] +
//             mat_A[830] * mat_B[989] +
//             mat_A[831] * mat_B[1021];
//  mat_C[830] <= 
//             mat_A[800] * mat_B[30] +
//             mat_A[801] * mat_B[62] +
//             mat_A[802] * mat_B[94] +
//             mat_A[803] * mat_B[126] +
//             mat_A[804] * mat_B[158] +
//             mat_A[805] * mat_B[190] +
//             mat_A[806] * mat_B[222] +
//             mat_A[807] * mat_B[254] +
//             mat_A[808] * mat_B[286] +
//             mat_A[809] * mat_B[318] +
//             mat_A[810] * mat_B[350] +
//             mat_A[811] * mat_B[382] +
//             mat_A[812] * mat_B[414] +
//             mat_A[813] * mat_B[446] +
//             mat_A[814] * mat_B[478] +
//             mat_A[815] * mat_B[510] +
//             mat_A[816] * mat_B[542] +
//             mat_A[817] * mat_B[574] +
//             mat_A[818] * mat_B[606] +
//             mat_A[819] * mat_B[638] +
//             mat_A[820] * mat_B[670] +
//             mat_A[821] * mat_B[702] +
//             mat_A[822] * mat_B[734] +
//             mat_A[823] * mat_B[766] +
//             mat_A[824] * mat_B[798] +
//             mat_A[825] * mat_B[830] +
//             mat_A[826] * mat_B[862] +
//             mat_A[827] * mat_B[894] +
//             mat_A[828] * mat_B[926] +
//             mat_A[829] * mat_B[958] +
//             mat_A[830] * mat_B[990] +
//             mat_A[831] * mat_B[1022];
//  mat_C[831] <= 
//             mat_A[800] * mat_B[31] +
//             mat_A[801] * mat_B[63] +
//             mat_A[802] * mat_B[95] +
//             mat_A[803] * mat_B[127] +
//             mat_A[804] * mat_B[159] +
//             mat_A[805] * mat_B[191] +
//             mat_A[806] * mat_B[223] +
//             mat_A[807] * mat_B[255] +
//             mat_A[808] * mat_B[287] +
//             mat_A[809] * mat_B[319] +
//             mat_A[810] * mat_B[351] +
//             mat_A[811] * mat_B[383] +
//             mat_A[812] * mat_B[415] +
//             mat_A[813] * mat_B[447] +
//             mat_A[814] * mat_B[479] +
//             mat_A[815] * mat_B[511] +
//             mat_A[816] * mat_B[543] +
//             mat_A[817] * mat_B[575] +
//             mat_A[818] * mat_B[607] +
//             mat_A[819] * mat_B[639] +
//             mat_A[820] * mat_B[671] +
//             mat_A[821] * mat_B[703] +
//             mat_A[822] * mat_B[735] +
//             mat_A[823] * mat_B[767] +
//             mat_A[824] * mat_B[799] +
//             mat_A[825] * mat_B[831] +
//             mat_A[826] * mat_B[863] +
//             mat_A[827] * mat_B[895] +
//             mat_A[828] * mat_B[927] +
//             mat_A[829] * mat_B[959] +
//             mat_A[830] * mat_B[991] +
//             mat_A[831] * mat_B[1023];
//  mat_C[832] <= 
//             mat_A[832] * mat_B[0] +
//             mat_A[833] * mat_B[32] +
//             mat_A[834] * mat_B[64] +
//             mat_A[835] * mat_B[96] +
//             mat_A[836] * mat_B[128] +
//             mat_A[837] * mat_B[160] +
//             mat_A[838] * mat_B[192] +
//             mat_A[839] * mat_B[224] +
//             mat_A[840] * mat_B[256] +
//             mat_A[841] * mat_B[288] +
//             mat_A[842] * mat_B[320] +
//             mat_A[843] * mat_B[352] +
//             mat_A[844] * mat_B[384] +
//             mat_A[845] * mat_B[416] +
//             mat_A[846] * mat_B[448] +
//             mat_A[847] * mat_B[480] +
//             mat_A[848] * mat_B[512] +
//             mat_A[849] * mat_B[544] +
//             mat_A[850] * mat_B[576] +
//             mat_A[851] * mat_B[608] +
//             mat_A[852] * mat_B[640] +
//             mat_A[853] * mat_B[672] +
//             mat_A[854] * mat_B[704] +
//             mat_A[855] * mat_B[736] +
//             mat_A[856] * mat_B[768] +
//             mat_A[857] * mat_B[800] +
//             mat_A[858] * mat_B[832] +
//             mat_A[859] * mat_B[864] +
//             mat_A[860] * mat_B[896] +
//             mat_A[861] * mat_B[928] +
//             mat_A[862] * mat_B[960] +
//             mat_A[863] * mat_B[992];
//  mat_C[833] <= 
//             mat_A[832] * mat_B[1] +
//             mat_A[833] * mat_B[33] +
//             mat_A[834] * mat_B[65] +
//             mat_A[835] * mat_B[97] +
//             mat_A[836] * mat_B[129] +
//             mat_A[837] * mat_B[161] +
//             mat_A[838] * mat_B[193] +
//             mat_A[839] * mat_B[225] +
//             mat_A[840] * mat_B[257] +
//             mat_A[841] * mat_B[289] +
//             mat_A[842] * mat_B[321] +
//             mat_A[843] * mat_B[353] +
//             mat_A[844] * mat_B[385] +
//             mat_A[845] * mat_B[417] +
//             mat_A[846] * mat_B[449] +
//             mat_A[847] * mat_B[481] +
//             mat_A[848] * mat_B[513] +
//             mat_A[849] * mat_B[545] +
//             mat_A[850] * mat_B[577] +
//             mat_A[851] * mat_B[609] +
//             mat_A[852] * mat_B[641] +
//             mat_A[853] * mat_B[673] +
//             mat_A[854] * mat_B[705] +
//             mat_A[855] * mat_B[737] +
//             mat_A[856] * mat_B[769] +
//             mat_A[857] * mat_B[801] +
//             mat_A[858] * mat_B[833] +
//             mat_A[859] * mat_B[865] +
//             mat_A[860] * mat_B[897] +
//             mat_A[861] * mat_B[929] +
//             mat_A[862] * mat_B[961] +
//             mat_A[863] * mat_B[993];
//  mat_C[834] <= 
//             mat_A[832] * mat_B[2] +
//             mat_A[833] * mat_B[34] +
//             mat_A[834] * mat_B[66] +
//             mat_A[835] * mat_B[98] +
//             mat_A[836] * mat_B[130] +
//             mat_A[837] * mat_B[162] +
//             mat_A[838] * mat_B[194] +
//             mat_A[839] * mat_B[226] +
//             mat_A[840] * mat_B[258] +
//             mat_A[841] * mat_B[290] +
//             mat_A[842] * mat_B[322] +
//             mat_A[843] * mat_B[354] +
//             mat_A[844] * mat_B[386] +
//             mat_A[845] * mat_B[418] +
//             mat_A[846] * mat_B[450] +
//             mat_A[847] * mat_B[482] +
//             mat_A[848] * mat_B[514] +
//             mat_A[849] * mat_B[546] +
//             mat_A[850] * mat_B[578] +
//             mat_A[851] * mat_B[610] +
//             mat_A[852] * mat_B[642] +
//             mat_A[853] * mat_B[674] +
//             mat_A[854] * mat_B[706] +
//             mat_A[855] * mat_B[738] +
//             mat_A[856] * mat_B[770] +
//             mat_A[857] * mat_B[802] +
//             mat_A[858] * mat_B[834] +
//             mat_A[859] * mat_B[866] +
//             mat_A[860] * mat_B[898] +
//             mat_A[861] * mat_B[930] +
//             mat_A[862] * mat_B[962] +
//             mat_A[863] * mat_B[994];
//  mat_C[835] <= 
//             mat_A[832] * mat_B[3] +
//             mat_A[833] * mat_B[35] +
//             mat_A[834] * mat_B[67] +
//             mat_A[835] * mat_B[99] +
//             mat_A[836] * mat_B[131] +
//             mat_A[837] * mat_B[163] +
//             mat_A[838] * mat_B[195] +
//             mat_A[839] * mat_B[227] +
//             mat_A[840] * mat_B[259] +
//             mat_A[841] * mat_B[291] +
//             mat_A[842] * mat_B[323] +
//             mat_A[843] * mat_B[355] +
//             mat_A[844] * mat_B[387] +
//             mat_A[845] * mat_B[419] +
//             mat_A[846] * mat_B[451] +
//             mat_A[847] * mat_B[483] +
//             mat_A[848] * mat_B[515] +
//             mat_A[849] * mat_B[547] +
//             mat_A[850] * mat_B[579] +
//             mat_A[851] * mat_B[611] +
//             mat_A[852] * mat_B[643] +
//             mat_A[853] * mat_B[675] +
//             mat_A[854] * mat_B[707] +
//             mat_A[855] * mat_B[739] +
//             mat_A[856] * mat_B[771] +
//             mat_A[857] * mat_B[803] +
//             mat_A[858] * mat_B[835] +
//             mat_A[859] * mat_B[867] +
//             mat_A[860] * mat_B[899] +
//             mat_A[861] * mat_B[931] +
//             mat_A[862] * mat_B[963] +
//             mat_A[863] * mat_B[995];
//  mat_C[836] <= 
//             mat_A[832] * mat_B[4] +
//             mat_A[833] * mat_B[36] +
//             mat_A[834] * mat_B[68] +
//             mat_A[835] * mat_B[100] +
//             mat_A[836] * mat_B[132] +
//             mat_A[837] * mat_B[164] +
//             mat_A[838] * mat_B[196] +
//             mat_A[839] * mat_B[228] +
//             mat_A[840] * mat_B[260] +
//             mat_A[841] * mat_B[292] +
//             mat_A[842] * mat_B[324] +
//             mat_A[843] * mat_B[356] +
//             mat_A[844] * mat_B[388] +
//             mat_A[845] * mat_B[420] +
//             mat_A[846] * mat_B[452] +
//             mat_A[847] * mat_B[484] +
//             mat_A[848] * mat_B[516] +
//             mat_A[849] * mat_B[548] +
//             mat_A[850] * mat_B[580] +
//             mat_A[851] * mat_B[612] +
//             mat_A[852] * mat_B[644] +
//             mat_A[853] * mat_B[676] +
//             mat_A[854] * mat_B[708] +
//             mat_A[855] * mat_B[740] +
//             mat_A[856] * mat_B[772] +
//             mat_A[857] * mat_B[804] +
//             mat_A[858] * mat_B[836] +
//             mat_A[859] * mat_B[868] +
//             mat_A[860] * mat_B[900] +
//             mat_A[861] * mat_B[932] +
//             mat_A[862] * mat_B[964] +
//             mat_A[863] * mat_B[996];
//  mat_C[837] <= 
//             mat_A[832] * mat_B[5] +
//             mat_A[833] * mat_B[37] +
//             mat_A[834] * mat_B[69] +
//             mat_A[835] * mat_B[101] +
//             mat_A[836] * mat_B[133] +
//             mat_A[837] * mat_B[165] +
//             mat_A[838] * mat_B[197] +
//             mat_A[839] * mat_B[229] +
//             mat_A[840] * mat_B[261] +
//             mat_A[841] * mat_B[293] +
//             mat_A[842] * mat_B[325] +
//             mat_A[843] * mat_B[357] +
//             mat_A[844] * mat_B[389] +
//             mat_A[845] * mat_B[421] +
//             mat_A[846] * mat_B[453] +
//             mat_A[847] * mat_B[485] +
//             mat_A[848] * mat_B[517] +
//             mat_A[849] * mat_B[549] +
//             mat_A[850] * mat_B[581] +
//             mat_A[851] * mat_B[613] +
//             mat_A[852] * mat_B[645] +
//             mat_A[853] * mat_B[677] +
//             mat_A[854] * mat_B[709] +
//             mat_A[855] * mat_B[741] +
//             mat_A[856] * mat_B[773] +
//             mat_A[857] * mat_B[805] +
//             mat_A[858] * mat_B[837] +
//             mat_A[859] * mat_B[869] +
//             mat_A[860] * mat_B[901] +
//             mat_A[861] * mat_B[933] +
//             mat_A[862] * mat_B[965] +
//             mat_A[863] * mat_B[997];
//  mat_C[838] <= 
//             mat_A[832] * mat_B[6] +
//             mat_A[833] * mat_B[38] +
//             mat_A[834] * mat_B[70] +
//             mat_A[835] * mat_B[102] +
//             mat_A[836] * mat_B[134] +
//             mat_A[837] * mat_B[166] +
//             mat_A[838] * mat_B[198] +
//             mat_A[839] * mat_B[230] +
//             mat_A[840] * mat_B[262] +
//             mat_A[841] * mat_B[294] +
//             mat_A[842] * mat_B[326] +
//             mat_A[843] * mat_B[358] +
//             mat_A[844] * mat_B[390] +
//             mat_A[845] * mat_B[422] +
//             mat_A[846] * mat_B[454] +
//             mat_A[847] * mat_B[486] +
//             mat_A[848] * mat_B[518] +
//             mat_A[849] * mat_B[550] +
//             mat_A[850] * mat_B[582] +
//             mat_A[851] * mat_B[614] +
//             mat_A[852] * mat_B[646] +
//             mat_A[853] * mat_B[678] +
//             mat_A[854] * mat_B[710] +
//             mat_A[855] * mat_B[742] +
//             mat_A[856] * mat_B[774] +
//             mat_A[857] * mat_B[806] +
//             mat_A[858] * mat_B[838] +
//             mat_A[859] * mat_B[870] +
//             mat_A[860] * mat_B[902] +
//             mat_A[861] * mat_B[934] +
//             mat_A[862] * mat_B[966] +
//             mat_A[863] * mat_B[998];
//  mat_C[839] <= 
//             mat_A[832] * mat_B[7] +
//             mat_A[833] * mat_B[39] +
//             mat_A[834] * mat_B[71] +
//             mat_A[835] * mat_B[103] +
//             mat_A[836] * mat_B[135] +
//             mat_A[837] * mat_B[167] +
//             mat_A[838] * mat_B[199] +
//             mat_A[839] * mat_B[231] +
//             mat_A[840] * mat_B[263] +
//             mat_A[841] * mat_B[295] +
//             mat_A[842] * mat_B[327] +
//             mat_A[843] * mat_B[359] +
//             mat_A[844] * mat_B[391] +
//             mat_A[845] * mat_B[423] +
//             mat_A[846] * mat_B[455] +
//             mat_A[847] * mat_B[487] +
//             mat_A[848] * mat_B[519] +
//             mat_A[849] * mat_B[551] +
//             mat_A[850] * mat_B[583] +
//             mat_A[851] * mat_B[615] +
//             mat_A[852] * mat_B[647] +
//             mat_A[853] * mat_B[679] +
//             mat_A[854] * mat_B[711] +
//             mat_A[855] * mat_B[743] +
//             mat_A[856] * mat_B[775] +
//             mat_A[857] * mat_B[807] +
//             mat_A[858] * mat_B[839] +
//             mat_A[859] * mat_B[871] +
//             mat_A[860] * mat_B[903] +
//             mat_A[861] * mat_B[935] +
//             mat_A[862] * mat_B[967] +
//             mat_A[863] * mat_B[999];
//  mat_C[840] <= 
//             mat_A[832] * mat_B[8] +
//             mat_A[833] * mat_B[40] +
//             mat_A[834] * mat_B[72] +
//             mat_A[835] * mat_B[104] +
//             mat_A[836] * mat_B[136] +
//             mat_A[837] * mat_B[168] +
//             mat_A[838] * mat_B[200] +
//             mat_A[839] * mat_B[232] +
//             mat_A[840] * mat_B[264] +
//             mat_A[841] * mat_B[296] +
//             mat_A[842] * mat_B[328] +
//             mat_A[843] * mat_B[360] +
//             mat_A[844] * mat_B[392] +
//             mat_A[845] * mat_B[424] +
//             mat_A[846] * mat_B[456] +
//             mat_A[847] * mat_B[488] +
//             mat_A[848] * mat_B[520] +
//             mat_A[849] * mat_B[552] +
//             mat_A[850] * mat_B[584] +
//             mat_A[851] * mat_B[616] +
//             mat_A[852] * mat_B[648] +
//             mat_A[853] * mat_B[680] +
//             mat_A[854] * mat_B[712] +
//             mat_A[855] * mat_B[744] +
//             mat_A[856] * mat_B[776] +
//             mat_A[857] * mat_B[808] +
//             mat_A[858] * mat_B[840] +
//             mat_A[859] * mat_B[872] +
//             mat_A[860] * mat_B[904] +
//             mat_A[861] * mat_B[936] +
//             mat_A[862] * mat_B[968] +
//             mat_A[863] * mat_B[1000];
//  mat_C[841] <= 
//             mat_A[832] * mat_B[9] +
//             mat_A[833] * mat_B[41] +
//             mat_A[834] * mat_B[73] +
//             mat_A[835] * mat_B[105] +
//             mat_A[836] * mat_B[137] +
//             mat_A[837] * mat_B[169] +
//             mat_A[838] * mat_B[201] +
//             mat_A[839] * mat_B[233] +
//             mat_A[840] * mat_B[265] +
//             mat_A[841] * mat_B[297] +
//             mat_A[842] * mat_B[329] +
//             mat_A[843] * mat_B[361] +
//             mat_A[844] * mat_B[393] +
//             mat_A[845] * mat_B[425] +
//             mat_A[846] * mat_B[457] +
//             mat_A[847] * mat_B[489] +
//             mat_A[848] * mat_B[521] +
//             mat_A[849] * mat_B[553] +
//             mat_A[850] * mat_B[585] +
//             mat_A[851] * mat_B[617] +
//             mat_A[852] * mat_B[649] +
//             mat_A[853] * mat_B[681] +
//             mat_A[854] * mat_B[713] +
//             mat_A[855] * mat_B[745] +
//             mat_A[856] * mat_B[777] +
//             mat_A[857] * mat_B[809] +
//             mat_A[858] * mat_B[841] +
//             mat_A[859] * mat_B[873] +
//             mat_A[860] * mat_B[905] +
//             mat_A[861] * mat_B[937] +
//             mat_A[862] * mat_B[969] +
//             mat_A[863] * mat_B[1001];
//  mat_C[842] <= 
//             mat_A[832] * mat_B[10] +
//             mat_A[833] * mat_B[42] +
//             mat_A[834] * mat_B[74] +
//             mat_A[835] * mat_B[106] +
//             mat_A[836] * mat_B[138] +
//             mat_A[837] * mat_B[170] +
//             mat_A[838] * mat_B[202] +
//             mat_A[839] * mat_B[234] +
//             mat_A[840] * mat_B[266] +
//             mat_A[841] * mat_B[298] +
//             mat_A[842] * mat_B[330] +
//             mat_A[843] * mat_B[362] +
//             mat_A[844] * mat_B[394] +
//             mat_A[845] * mat_B[426] +
//             mat_A[846] * mat_B[458] +
//             mat_A[847] * mat_B[490] +
//             mat_A[848] * mat_B[522] +
//             mat_A[849] * mat_B[554] +
//             mat_A[850] * mat_B[586] +
//             mat_A[851] * mat_B[618] +
//             mat_A[852] * mat_B[650] +
//             mat_A[853] * mat_B[682] +
//             mat_A[854] * mat_B[714] +
//             mat_A[855] * mat_B[746] +
//             mat_A[856] * mat_B[778] +
//             mat_A[857] * mat_B[810] +
//             mat_A[858] * mat_B[842] +
//             mat_A[859] * mat_B[874] +
//             mat_A[860] * mat_B[906] +
//             mat_A[861] * mat_B[938] +
//             mat_A[862] * mat_B[970] +
//             mat_A[863] * mat_B[1002];
//  mat_C[843] <= 
//             mat_A[832] * mat_B[11] +
//             mat_A[833] * mat_B[43] +
//             mat_A[834] * mat_B[75] +
//             mat_A[835] * mat_B[107] +
//             mat_A[836] * mat_B[139] +
//             mat_A[837] * mat_B[171] +
//             mat_A[838] * mat_B[203] +
//             mat_A[839] * mat_B[235] +
//             mat_A[840] * mat_B[267] +
//             mat_A[841] * mat_B[299] +
//             mat_A[842] * mat_B[331] +
//             mat_A[843] * mat_B[363] +
//             mat_A[844] * mat_B[395] +
//             mat_A[845] * mat_B[427] +
//             mat_A[846] * mat_B[459] +
//             mat_A[847] * mat_B[491] +
//             mat_A[848] * mat_B[523] +
//             mat_A[849] * mat_B[555] +
//             mat_A[850] * mat_B[587] +
//             mat_A[851] * mat_B[619] +
//             mat_A[852] * mat_B[651] +
//             mat_A[853] * mat_B[683] +
//             mat_A[854] * mat_B[715] +
//             mat_A[855] * mat_B[747] +
//             mat_A[856] * mat_B[779] +
//             mat_A[857] * mat_B[811] +
//             mat_A[858] * mat_B[843] +
//             mat_A[859] * mat_B[875] +
//             mat_A[860] * mat_B[907] +
//             mat_A[861] * mat_B[939] +
//             mat_A[862] * mat_B[971] +
//             mat_A[863] * mat_B[1003];
//  mat_C[844] <= 
//             mat_A[832] * mat_B[12] +
//             mat_A[833] * mat_B[44] +
//             mat_A[834] * mat_B[76] +
//             mat_A[835] * mat_B[108] +
//             mat_A[836] * mat_B[140] +
//             mat_A[837] * mat_B[172] +
//             mat_A[838] * mat_B[204] +
//             mat_A[839] * mat_B[236] +
//             mat_A[840] * mat_B[268] +
//             mat_A[841] * mat_B[300] +
//             mat_A[842] * mat_B[332] +
//             mat_A[843] * mat_B[364] +
//             mat_A[844] * mat_B[396] +
//             mat_A[845] * mat_B[428] +
//             mat_A[846] * mat_B[460] +
//             mat_A[847] * mat_B[492] +
//             mat_A[848] * mat_B[524] +
//             mat_A[849] * mat_B[556] +
//             mat_A[850] * mat_B[588] +
//             mat_A[851] * mat_B[620] +
//             mat_A[852] * mat_B[652] +
//             mat_A[853] * mat_B[684] +
//             mat_A[854] * mat_B[716] +
//             mat_A[855] * mat_B[748] +
//             mat_A[856] * mat_B[780] +
//             mat_A[857] * mat_B[812] +
//             mat_A[858] * mat_B[844] +
//             mat_A[859] * mat_B[876] +
//             mat_A[860] * mat_B[908] +
//             mat_A[861] * mat_B[940] +
//             mat_A[862] * mat_B[972] +
//             mat_A[863] * mat_B[1004];
//  mat_C[845] <= 
//             mat_A[832] * mat_B[13] +
//             mat_A[833] * mat_B[45] +
//             mat_A[834] * mat_B[77] +
//             mat_A[835] * mat_B[109] +
//             mat_A[836] * mat_B[141] +
//             mat_A[837] * mat_B[173] +
//             mat_A[838] * mat_B[205] +
//             mat_A[839] * mat_B[237] +
//             mat_A[840] * mat_B[269] +
//             mat_A[841] * mat_B[301] +
//             mat_A[842] * mat_B[333] +
//             mat_A[843] * mat_B[365] +
//             mat_A[844] * mat_B[397] +
//             mat_A[845] * mat_B[429] +
//             mat_A[846] * mat_B[461] +
//             mat_A[847] * mat_B[493] +
//             mat_A[848] * mat_B[525] +
//             mat_A[849] * mat_B[557] +
//             mat_A[850] * mat_B[589] +
//             mat_A[851] * mat_B[621] +
//             mat_A[852] * mat_B[653] +
//             mat_A[853] * mat_B[685] +
//             mat_A[854] * mat_B[717] +
//             mat_A[855] * mat_B[749] +
//             mat_A[856] * mat_B[781] +
//             mat_A[857] * mat_B[813] +
//             mat_A[858] * mat_B[845] +
//             mat_A[859] * mat_B[877] +
//             mat_A[860] * mat_B[909] +
//             mat_A[861] * mat_B[941] +
//             mat_A[862] * mat_B[973] +
//             mat_A[863] * mat_B[1005];
//  mat_C[846] <= 
//             mat_A[832] * mat_B[14] +
//             mat_A[833] * mat_B[46] +
//             mat_A[834] * mat_B[78] +
//             mat_A[835] * mat_B[110] +
//             mat_A[836] * mat_B[142] +
//             mat_A[837] * mat_B[174] +
//             mat_A[838] * mat_B[206] +
//             mat_A[839] * mat_B[238] +
//             mat_A[840] * mat_B[270] +
//             mat_A[841] * mat_B[302] +
//             mat_A[842] * mat_B[334] +
//             mat_A[843] * mat_B[366] +
//             mat_A[844] * mat_B[398] +
//             mat_A[845] * mat_B[430] +
//             mat_A[846] * mat_B[462] +
//             mat_A[847] * mat_B[494] +
//             mat_A[848] * mat_B[526] +
//             mat_A[849] * mat_B[558] +
//             mat_A[850] * mat_B[590] +
//             mat_A[851] * mat_B[622] +
//             mat_A[852] * mat_B[654] +
//             mat_A[853] * mat_B[686] +
//             mat_A[854] * mat_B[718] +
//             mat_A[855] * mat_B[750] +
//             mat_A[856] * mat_B[782] +
//             mat_A[857] * mat_B[814] +
//             mat_A[858] * mat_B[846] +
//             mat_A[859] * mat_B[878] +
//             mat_A[860] * mat_B[910] +
//             mat_A[861] * mat_B[942] +
//             mat_A[862] * mat_B[974] +
//             mat_A[863] * mat_B[1006];
//  mat_C[847] <= 
//             mat_A[832] * mat_B[15] +
//             mat_A[833] * mat_B[47] +
//             mat_A[834] * mat_B[79] +
//             mat_A[835] * mat_B[111] +
//             mat_A[836] * mat_B[143] +
//             mat_A[837] * mat_B[175] +
//             mat_A[838] * mat_B[207] +
//             mat_A[839] * mat_B[239] +
//             mat_A[840] * mat_B[271] +
//             mat_A[841] * mat_B[303] +
//             mat_A[842] * mat_B[335] +
//             mat_A[843] * mat_B[367] +
//             mat_A[844] * mat_B[399] +
//             mat_A[845] * mat_B[431] +
//             mat_A[846] * mat_B[463] +
//             mat_A[847] * mat_B[495] +
//             mat_A[848] * mat_B[527] +
//             mat_A[849] * mat_B[559] +
//             mat_A[850] * mat_B[591] +
//             mat_A[851] * mat_B[623] +
//             mat_A[852] * mat_B[655] +
//             mat_A[853] * mat_B[687] +
//             mat_A[854] * mat_B[719] +
//             mat_A[855] * mat_B[751] +
//             mat_A[856] * mat_B[783] +
//             mat_A[857] * mat_B[815] +
//             mat_A[858] * mat_B[847] +
//             mat_A[859] * mat_B[879] +
//             mat_A[860] * mat_B[911] +
//             mat_A[861] * mat_B[943] +
//             mat_A[862] * mat_B[975] +
//             mat_A[863] * mat_B[1007];
//  mat_C[848] <= 
//             mat_A[832] * mat_B[16] +
//             mat_A[833] * mat_B[48] +
//             mat_A[834] * mat_B[80] +
//             mat_A[835] * mat_B[112] +
//             mat_A[836] * mat_B[144] +
//             mat_A[837] * mat_B[176] +
//             mat_A[838] * mat_B[208] +
//             mat_A[839] * mat_B[240] +
//             mat_A[840] * mat_B[272] +
//             mat_A[841] * mat_B[304] +
//             mat_A[842] * mat_B[336] +
//             mat_A[843] * mat_B[368] +
//             mat_A[844] * mat_B[400] +
//             mat_A[845] * mat_B[432] +
//             mat_A[846] * mat_B[464] +
//             mat_A[847] * mat_B[496] +
//             mat_A[848] * mat_B[528] +
//             mat_A[849] * mat_B[560] +
//             mat_A[850] * mat_B[592] +
//             mat_A[851] * mat_B[624] +
//             mat_A[852] * mat_B[656] +
//             mat_A[853] * mat_B[688] +
//             mat_A[854] * mat_B[720] +
//             mat_A[855] * mat_B[752] +
//             mat_A[856] * mat_B[784] +
//             mat_A[857] * mat_B[816] +
//             mat_A[858] * mat_B[848] +
//             mat_A[859] * mat_B[880] +
//             mat_A[860] * mat_B[912] +
//             mat_A[861] * mat_B[944] +
//             mat_A[862] * mat_B[976] +
//             mat_A[863] * mat_B[1008];
//  mat_C[849] <= 
//             mat_A[832] * mat_B[17] +
//             mat_A[833] * mat_B[49] +
//             mat_A[834] * mat_B[81] +
//             mat_A[835] * mat_B[113] +
//             mat_A[836] * mat_B[145] +
//             mat_A[837] * mat_B[177] +
//             mat_A[838] * mat_B[209] +
//             mat_A[839] * mat_B[241] +
//             mat_A[840] * mat_B[273] +
//             mat_A[841] * mat_B[305] +
//             mat_A[842] * mat_B[337] +
//             mat_A[843] * mat_B[369] +
//             mat_A[844] * mat_B[401] +
//             mat_A[845] * mat_B[433] +
//             mat_A[846] * mat_B[465] +
//             mat_A[847] * mat_B[497] +
//             mat_A[848] * mat_B[529] +
//             mat_A[849] * mat_B[561] +
//             mat_A[850] * mat_B[593] +
//             mat_A[851] * mat_B[625] +
//             mat_A[852] * mat_B[657] +
//             mat_A[853] * mat_B[689] +
//             mat_A[854] * mat_B[721] +
//             mat_A[855] * mat_B[753] +
//             mat_A[856] * mat_B[785] +
//             mat_A[857] * mat_B[817] +
//             mat_A[858] * mat_B[849] +
//             mat_A[859] * mat_B[881] +
//             mat_A[860] * mat_B[913] +
//             mat_A[861] * mat_B[945] +
//             mat_A[862] * mat_B[977] +
//             mat_A[863] * mat_B[1009];
//  mat_C[850] <= 
//             mat_A[832] * mat_B[18] +
//             mat_A[833] * mat_B[50] +
//             mat_A[834] * mat_B[82] +
//             mat_A[835] * mat_B[114] +
//             mat_A[836] * mat_B[146] +
//             mat_A[837] * mat_B[178] +
//             mat_A[838] * mat_B[210] +
//             mat_A[839] * mat_B[242] +
//             mat_A[840] * mat_B[274] +
//             mat_A[841] * mat_B[306] +
//             mat_A[842] * mat_B[338] +
//             mat_A[843] * mat_B[370] +
//             mat_A[844] * mat_B[402] +
//             mat_A[845] * mat_B[434] +
//             mat_A[846] * mat_B[466] +
//             mat_A[847] * mat_B[498] +
//             mat_A[848] * mat_B[530] +
//             mat_A[849] * mat_B[562] +
//             mat_A[850] * mat_B[594] +
//             mat_A[851] * mat_B[626] +
//             mat_A[852] * mat_B[658] +
//             mat_A[853] * mat_B[690] +
//             mat_A[854] * mat_B[722] +
//             mat_A[855] * mat_B[754] +
//             mat_A[856] * mat_B[786] +
//             mat_A[857] * mat_B[818] +
//             mat_A[858] * mat_B[850] +
//             mat_A[859] * mat_B[882] +
//             mat_A[860] * mat_B[914] +
//             mat_A[861] * mat_B[946] +
//             mat_A[862] * mat_B[978] +
//             mat_A[863] * mat_B[1010];
//  mat_C[851] <= 
//             mat_A[832] * mat_B[19] +
//             mat_A[833] * mat_B[51] +
//             mat_A[834] * mat_B[83] +
//             mat_A[835] * mat_B[115] +
//             mat_A[836] * mat_B[147] +
//             mat_A[837] * mat_B[179] +
//             mat_A[838] * mat_B[211] +
//             mat_A[839] * mat_B[243] +
//             mat_A[840] * mat_B[275] +
//             mat_A[841] * mat_B[307] +
//             mat_A[842] * mat_B[339] +
//             mat_A[843] * mat_B[371] +
//             mat_A[844] * mat_B[403] +
//             mat_A[845] * mat_B[435] +
//             mat_A[846] * mat_B[467] +
//             mat_A[847] * mat_B[499] +
//             mat_A[848] * mat_B[531] +
//             mat_A[849] * mat_B[563] +
//             mat_A[850] * mat_B[595] +
//             mat_A[851] * mat_B[627] +
//             mat_A[852] * mat_B[659] +
//             mat_A[853] * mat_B[691] +
//             mat_A[854] * mat_B[723] +
//             mat_A[855] * mat_B[755] +
//             mat_A[856] * mat_B[787] +
//             mat_A[857] * mat_B[819] +
//             mat_A[858] * mat_B[851] +
//             mat_A[859] * mat_B[883] +
//             mat_A[860] * mat_B[915] +
//             mat_A[861] * mat_B[947] +
//             mat_A[862] * mat_B[979] +
//             mat_A[863] * mat_B[1011];
//  mat_C[852] <= 
//             mat_A[832] * mat_B[20] +
//             mat_A[833] * mat_B[52] +
//             mat_A[834] * mat_B[84] +
//             mat_A[835] * mat_B[116] +
//             mat_A[836] * mat_B[148] +
//             mat_A[837] * mat_B[180] +
//             mat_A[838] * mat_B[212] +
//             mat_A[839] * mat_B[244] +
//             mat_A[840] * mat_B[276] +
//             mat_A[841] * mat_B[308] +
//             mat_A[842] * mat_B[340] +
//             mat_A[843] * mat_B[372] +
//             mat_A[844] * mat_B[404] +
//             mat_A[845] * mat_B[436] +
//             mat_A[846] * mat_B[468] +
//             mat_A[847] * mat_B[500] +
//             mat_A[848] * mat_B[532] +
//             mat_A[849] * mat_B[564] +
//             mat_A[850] * mat_B[596] +
//             mat_A[851] * mat_B[628] +
//             mat_A[852] * mat_B[660] +
//             mat_A[853] * mat_B[692] +
//             mat_A[854] * mat_B[724] +
//             mat_A[855] * mat_B[756] +
//             mat_A[856] * mat_B[788] +
//             mat_A[857] * mat_B[820] +
//             mat_A[858] * mat_B[852] +
//             mat_A[859] * mat_B[884] +
//             mat_A[860] * mat_B[916] +
//             mat_A[861] * mat_B[948] +
//             mat_A[862] * mat_B[980] +
//             mat_A[863] * mat_B[1012];
//  mat_C[853] <= 
//             mat_A[832] * mat_B[21] +
//             mat_A[833] * mat_B[53] +
//             mat_A[834] * mat_B[85] +
//             mat_A[835] * mat_B[117] +
//             mat_A[836] * mat_B[149] +
//             mat_A[837] * mat_B[181] +
//             mat_A[838] * mat_B[213] +
//             mat_A[839] * mat_B[245] +
//             mat_A[840] * mat_B[277] +
//             mat_A[841] * mat_B[309] +
//             mat_A[842] * mat_B[341] +
//             mat_A[843] * mat_B[373] +
//             mat_A[844] * mat_B[405] +
//             mat_A[845] * mat_B[437] +
//             mat_A[846] * mat_B[469] +
//             mat_A[847] * mat_B[501] +
//             mat_A[848] * mat_B[533] +
//             mat_A[849] * mat_B[565] +
//             mat_A[850] * mat_B[597] +
//             mat_A[851] * mat_B[629] +
//             mat_A[852] * mat_B[661] +
//             mat_A[853] * mat_B[693] +
//             mat_A[854] * mat_B[725] +
//             mat_A[855] * mat_B[757] +
//             mat_A[856] * mat_B[789] +
//             mat_A[857] * mat_B[821] +
//             mat_A[858] * mat_B[853] +
//             mat_A[859] * mat_B[885] +
//             mat_A[860] * mat_B[917] +
//             mat_A[861] * mat_B[949] +
//             mat_A[862] * mat_B[981] +
//             mat_A[863] * mat_B[1013];
//  mat_C[854] <= 
//             mat_A[832] * mat_B[22] +
//             mat_A[833] * mat_B[54] +
//             mat_A[834] * mat_B[86] +
//             mat_A[835] * mat_B[118] +
//             mat_A[836] * mat_B[150] +
//             mat_A[837] * mat_B[182] +
//             mat_A[838] * mat_B[214] +
//             mat_A[839] * mat_B[246] +
//             mat_A[840] * mat_B[278] +
//             mat_A[841] * mat_B[310] +
//             mat_A[842] * mat_B[342] +
//             mat_A[843] * mat_B[374] +
//             mat_A[844] * mat_B[406] +
//             mat_A[845] * mat_B[438] +
//             mat_A[846] * mat_B[470] +
//             mat_A[847] * mat_B[502] +
//             mat_A[848] * mat_B[534] +
//             mat_A[849] * mat_B[566] +
//             mat_A[850] * mat_B[598] +
//             mat_A[851] * mat_B[630] +
//             mat_A[852] * mat_B[662] +
//             mat_A[853] * mat_B[694] +
//             mat_A[854] * mat_B[726] +
//             mat_A[855] * mat_B[758] +
//             mat_A[856] * mat_B[790] +
//             mat_A[857] * mat_B[822] +
//             mat_A[858] * mat_B[854] +
//             mat_A[859] * mat_B[886] +
//             mat_A[860] * mat_B[918] +
//             mat_A[861] * mat_B[950] +
//             mat_A[862] * mat_B[982] +
//             mat_A[863] * mat_B[1014];
//  mat_C[855] <= 
//             mat_A[832] * mat_B[23] +
//             mat_A[833] * mat_B[55] +
//             mat_A[834] * mat_B[87] +
//             mat_A[835] * mat_B[119] +
//             mat_A[836] * mat_B[151] +
//             mat_A[837] * mat_B[183] +
//             mat_A[838] * mat_B[215] +
//             mat_A[839] * mat_B[247] +
//             mat_A[840] * mat_B[279] +
//             mat_A[841] * mat_B[311] +
//             mat_A[842] * mat_B[343] +
//             mat_A[843] * mat_B[375] +
//             mat_A[844] * mat_B[407] +
//             mat_A[845] * mat_B[439] +
//             mat_A[846] * mat_B[471] +
//             mat_A[847] * mat_B[503] +
//             mat_A[848] * mat_B[535] +
//             mat_A[849] * mat_B[567] +
//             mat_A[850] * mat_B[599] +
//             mat_A[851] * mat_B[631] +
//             mat_A[852] * mat_B[663] +
//             mat_A[853] * mat_B[695] +
//             mat_A[854] * mat_B[727] +
//             mat_A[855] * mat_B[759] +
//             mat_A[856] * mat_B[791] +
//             mat_A[857] * mat_B[823] +
//             mat_A[858] * mat_B[855] +
//             mat_A[859] * mat_B[887] +
//             mat_A[860] * mat_B[919] +
//             mat_A[861] * mat_B[951] +
//             mat_A[862] * mat_B[983] +
//             mat_A[863] * mat_B[1015];
//  mat_C[856] <= 
//             mat_A[832] * mat_B[24] +
//             mat_A[833] * mat_B[56] +
//             mat_A[834] * mat_B[88] +
//             mat_A[835] * mat_B[120] +
//             mat_A[836] * mat_B[152] +
//             mat_A[837] * mat_B[184] +
//             mat_A[838] * mat_B[216] +
//             mat_A[839] * mat_B[248] +
//             mat_A[840] * mat_B[280] +
//             mat_A[841] * mat_B[312] +
//             mat_A[842] * mat_B[344] +
//             mat_A[843] * mat_B[376] +
//             mat_A[844] * mat_B[408] +
//             mat_A[845] * mat_B[440] +
//             mat_A[846] * mat_B[472] +
//             mat_A[847] * mat_B[504] +
//             mat_A[848] * mat_B[536] +
//             mat_A[849] * mat_B[568] +
//             mat_A[850] * mat_B[600] +
//             mat_A[851] * mat_B[632] +
//             mat_A[852] * mat_B[664] +
//             mat_A[853] * mat_B[696] +
//             mat_A[854] * mat_B[728] +
//             mat_A[855] * mat_B[760] +
//             mat_A[856] * mat_B[792] +
//             mat_A[857] * mat_B[824] +
//             mat_A[858] * mat_B[856] +
//             mat_A[859] * mat_B[888] +
//             mat_A[860] * mat_B[920] +
//             mat_A[861] * mat_B[952] +
//             mat_A[862] * mat_B[984] +
//             mat_A[863] * mat_B[1016];
//  mat_C[857] <= 
//             mat_A[832] * mat_B[25] +
//             mat_A[833] * mat_B[57] +
//             mat_A[834] * mat_B[89] +
//             mat_A[835] * mat_B[121] +
//             mat_A[836] * mat_B[153] +
//             mat_A[837] * mat_B[185] +
//             mat_A[838] * mat_B[217] +
//             mat_A[839] * mat_B[249] +
//             mat_A[840] * mat_B[281] +
//             mat_A[841] * mat_B[313] +
//             mat_A[842] * mat_B[345] +
//             mat_A[843] * mat_B[377] +
//             mat_A[844] * mat_B[409] +
//             mat_A[845] * mat_B[441] +
//             mat_A[846] * mat_B[473] +
//             mat_A[847] * mat_B[505] +
//             mat_A[848] * mat_B[537] +
//             mat_A[849] * mat_B[569] +
//             mat_A[850] * mat_B[601] +
//             mat_A[851] * mat_B[633] +
//             mat_A[852] * mat_B[665] +
//             mat_A[853] * mat_B[697] +
//             mat_A[854] * mat_B[729] +
//             mat_A[855] * mat_B[761] +
//             mat_A[856] * mat_B[793] +
//             mat_A[857] * mat_B[825] +
//             mat_A[858] * mat_B[857] +
//             mat_A[859] * mat_B[889] +
//             mat_A[860] * mat_B[921] +
//             mat_A[861] * mat_B[953] +
//             mat_A[862] * mat_B[985] +
//             mat_A[863] * mat_B[1017];
//  mat_C[858] <= 
//             mat_A[832] * mat_B[26] +
//             mat_A[833] * mat_B[58] +
//             mat_A[834] * mat_B[90] +
//             mat_A[835] * mat_B[122] +
//             mat_A[836] * mat_B[154] +
//             mat_A[837] * mat_B[186] +
//             mat_A[838] * mat_B[218] +
//             mat_A[839] * mat_B[250] +
//             mat_A[840] * mat_B[282] +
//             mat_A[841] * mat_B[314] +
//             mat_A[842] * mat_B[346] +
//             mat_A[843] * mat_B[378] +
//             mat_A[844] * mat_B[410] +
//             mat_A[845] * mat_B[442] +
//             mat_A[846] * mat_B[474] +
//             mat_A[847] * mat_B[506] +
//             mat_A[848] * mat_B[538] +
//             mat_A[849] * mat_B[570] +
//             mat_A[850] * mat_B[602] +
//             mat_A[851] * mat_B[634] +
//             mat_A[852] * mat_B[666] +
//             mat_A[853] * mat_B[698] +
//             mat_A[854] * mat_B[730] +
//             mat_A[855] * mat_B[762] +
//             mat_A[856] * mat_B[794] +
//             mat_A[857] * mat_B[826] +
//             mat_A[858] * mat_B[858] +
//             mat_A[859] * mat_B[890] +
//             mat_A[860] * mat_B[922] +
//             mat_A[861] * mat_B[954] +
//             mat_A[862] * mat_B[986] +
//             mat_A[863] * mat_B[1018];
//  mat_C[859] <= 
//             mat_A[832] * mat_B[27] +
//             mat_A[833] * mat_B[59] +
//             mat_A[834] * mat_B[91] +
//             mat_A[835] * mat_B[123] +
//             mat_A[836] * mat_B[155] +
//             mat_A[837] * mat_B[187] +
//             mat_A[838] * mat_B[219] +
//             mat_A[839] * mat_B[251] +
//             mat_A[840] * mat_B[283] +
//             mat_A[841] * mat_B[315] +
//             mat_A[842] * mat_B[347] +
//             mat_A[843] * mat_B[379] +
//             mat_A[844] * mat_B[411] +
//             mat_A[845] * mat_B[443] +
//             mat_A[846] * mat_B[475] +
//             mat_A[847] * mat_B[507] +
//             mat_A[848] * mat_B[539] +
//             mat_A[849] * mat_B[571] +
//             mat_A[850] * mat_B[603] +
//             mat_A[851] * mat_B[635] +
//             mat_A[852] * mat_B[667] +
//             mat_A[853] * mat_B[699] +
//             mat_A[854] * mat_B[731] +
//             mat_A[855] * mat_B[763] +
//             mat_A[856] * mat_B[795] +
//             mat_A[857] * mat_B[827] +
//             mat_A[858] * mat_B[859] +
//             mat_A[859] * mat_B[891] +
//             mat_A[860] * mat_B[923] +
//             mat_A[861] * mat_B[955] +
//             mat_A[862] * mat_B[987] +
//             mat_A[863] * mat_B[1019];
//  mat_C[860] <= 
//             mat_A[832] * mat_B[28] +
//             mat_A[833] * mat_B[60] +
//             mat_A[834] * mat_B[92] +
//             mat_A[835] * mat_B[124] +
//             mat_A[836] * mat_B[156] +
//             mat_A[837] * mat_B[188] +
//             mat_A[838] * mat_B[220] +
//             mat_A[839] * mat_B[252] +
//             mat_A[840] * mat_B[284] +
//             mat_A[841] * mat_B[316] +
//             mat_A[842] * mat_B[348] +
//             mat_A[843] * mat_B[380] +
//             mat_A[844] * mat_B[412] +
//             mat_A[845] * mat_B[444] +
//             mat_A[846] * mat_B[476] +
//             mat_A[847] * mat_B[508] +
//             mat_A[848] * mat_B[540] +
//             mat_A[849] * mat_B[572] +
//             mat_A[850] * mat_B[604] +
//             mat_A[851] * mat_B[636] +
//             mat_A[852] * mat_B[668] +
//             mat_A[853] * mat_B[700] +
//             mat_A[854] * mat_B[732] +
//             mat_A[855] * mat_B[764] +
//             mat_A[856] * mat_B[796] +
//             mat_A[857] * mat_B[828] +
//             mat_A[858] * mat_B[860] +
//             mat_A[859] * mat_B[892] +
//             mat_A[860] * mat_B[924] +
//             mat_A[861] * mat_B[956] +
//             mat_A[862] * mat_B[988] +
//             mat_A[863] * mat_B[1020];
//  mat_C[861] <= 
//             mat_A[832] * mat_B[29] +
//             mat_A[833] * mat_B[61] +
//             mat_A[834] * mat_B[93] +
//             mat_A[835] * mat_B[125] +
//             mat_A[836] * mat_B[157] +
//             mat_A[837] * mat_B[189] +
//             mat_A[838] * mat_B[221] +
//             mat_A[839] * mat_B[253] +
//             mat_A[840] * mat_B[285] +
//             mat_A[841] * mat_B[317] +
//             mat_A[842] * mat_B[349] +
//             mat_A[843] * mat_B[381] +
//             mat_A[844] * mat_B[413] +
//             mat_A[845] * mat_B[445] +
//             mat_A[846] * mat_B[477] +
//             mat_A[847] * mat_B[509] +
//             mat_A[848] * mat_B[541] +
//             mat_A[849] * mat_B[573] +
//             mat_A[850] * mat_B[605] +
//             mat_A[851] * mat_B[637] +
//             mat_A[852] * mat_B[669] +
//             mat_A[853] * mat_B[701] +
//             mat_A[854] * mat_B[733] +
//             mat_A[855] * mat_B[765] +
//             mat_A[856] * mat_B[797] +
//             mat_A[857] * mat_B[829] +
//             mat_A[858] * mat_B[861] +
//             mat_A[859] * mat_B[893] +
//             mat_A[860] * mat_B[925] +
//             mat_A[861] * mat_B[957] +
//             mat_A[862] * mat_B[989] +
//             mat_A[863] * mat_B[1021];
//  mat_C[862] <= 
//             mat_A[832] * mat_B[30] +
//             mat_A[833] * mat_B[62] +
//             mat_A[834] * mat_B[94] +
//             mat_A[835] * mat_B[126] +
//             mat_A[836] * mat_B[158] +
//             mat_A[837] * mat_B[190] +
//             mat_A[838] * mat_B[222] +
//             mat_A[839] * mat_B[254] +
//             mat_A[840] * mat_B[286] +
//             mat_A[841] * mat_B[318] +
//             mat_A[842] * mat_B[350] +
//             mat_A[843] * mat_B[382] +
//             mat_A[844] * mat_B[414] +
//             mat_A[845] * mat_B[446] +
//             mat_A[846] * mat_B[478] +
//             mat_A[847] * mat_B[510] +
//             mat_A[848] * mat_B[542] +
//             mat_A[849] * mat_B[574] +
//             mat_A[850] * mat_B[606] +
//             mat_A[851] * mat_B[638] +
//             mat_A[852] * mat_B[670] +
//             mat_A[853] * mat_B[702] +
//             mat_A[854] * mat_B[734] +
//             mat_A[855] * mat_B[766] +
//             mat_A[856] * mat_B[798] +
//             mat_A[857] * mat_B[830] +
//             mat_A[858] * mat_B[862] +
//             mat_A[859] * mat_B[894] +
//             mat_A[860] * mat_B[926] +
//             mat_A[861] * mat_B[958] +
//             mat_A[862] * mat_B[990] +
//             mat_A[863] * mat_B[1022];
//  mat_C[863] <= 
//             mat_A[832] * mat_B[31] +
//             mat_A[833] * mat_B[63] +
//             mat_A[834] * mat_B[95] +
//             mat_A[835] * mat_B[127] +
//             mat_A[836] * mat_B[159] +
//             mat_A[837] * mat_B[191] +
//             mat_A[838] * mat_B[223] +
//             mat_A[839] * mat_B[255] +
//             mat_A[840] * mat_B[287] +
//             mat_A[841] * mat_B[319] +
//             mat_A[842] * mat_B[351] +
//             mat_A[843] * mat_B[383] +
//             mat_A[844] * mat_B[415] +
//             mat_A[845] * mat_B[447] +
//             mat_A[846] * mat_B[479] +
//             mat_A[847] * mat_B[511] +
//             mat_A[848] * mat_B[543] +
//             mat_A[849] * mat_B[575] +
//             mat_A[850] * mat_B[607] +
//             mat_A[851] * mat_B[639] +
//             mat_A[852] * mat_B[671] +
//             mat_A[853] * mat_B[703] +
//             mat_A[854] * mat_B[735] +
//             mat_A[855] * mat_B[767] +
//             mat_A[856] * mat_B[799] +
//             mat_A[857] * mat_B[831] +
//             mat_A[858] * mat_B[863] +
//             mat_A[859] * mat_B[895] +
//             mat_A[860] * mat_B[927] +
//             mat_A[861] * mat_B[959] +
//             mat_A[862] * mat_B[991] +
//             mat_A[863] * mat_B[1023];
//  mat_C[864] <= 
//             mat_A[864] * mat_B[0] +
//             mat_A[865] * mat_B[32] +
//             mat_A[866] * mat_B[64] +
//             mat_A[867] * mat_B[96] +
//             mat_A[868] * mat_B[128] +
//             mat_A[869] * mat_B[160] +
//             mat_A[870] * mat_B[192] +
//             mat_A[871] * mat_B[224] +
//             mat_A[872] * mat_B[256] +
//             mat_A[873] * mat_B[288] +
//             mat_A[874] * mat_B[320] +
//             mat_A[875] * mat_B[352] +
//             mat_A[876] * mat_B[384] +
//             mat_A[877] * mat_B[416] +
//             mat_A[878] * mat_B[448] +
//             mat_A[879] * mat_B[480] +
//             mat_A[880] * mat_B[512] +
//             mat_A[881] * mat_B[544] +
//             mat_A[882] * mat_B[576] +
//             mat_A[883] * mat_B[608] +
//             mat_A[884] * mat_B[640] +
//             mat_A[885] * mat_B[672] +
//             mat_A[886] * mat_B[704] +
//             mat_A[887] * mat_B[736] +
//             mat_A[888] * mat_B[768] +
//             mat_A[889] * mat_B[800] +
//             mat_A[890] * mat_B[832] +
//             mat_A[891] * mat_B[864] +
//             mat_A[892] * mat_B[896] +
//             mat_A[893] * mat_B[928] +
//             mat_A[894] * mat_B[960] +
//             mat_A[895] * mat_B[992];
//  mat_C[865] <= 
//             mat_A[864] * mat_B[1] +
//             mat_A[865] * mat_B[33] +
//             mat_A[866] * mat_B[65] +
//             mat_A[867] * mat_B[97] +
//             mat_A[868] * mat_B[129] +
//             mat_A[869] * mat_B[161] +
//             mat_A[870] * mat_B[193] +
//             mat_A[871] * mat_B[225] +
//             mat_A[872] * mat_B[257] +
//             mat_A[873] * mat_B[289] +
//             mat_A[874] * mat_B[321] +
//             mat_A[875] * mat_B[353] +
//             mat_A[876] * mat_B[385] +
//             mat_A[877] * mat_B[417] +
//             mat_A[878] * mat_B[449] +
//             mat_A[879] * mat_B[481] +
//             mat_A[880] * mat_B[513] +
//             mat_A[881] * mat_B[545] +
//             mat_A[882] * mat_B[577] +
//             mat_A[883] * mat_B[609] +
//             mat_A[884] * mat_B[641] +
//             mat_A[885] * mat_B[673] +
//             mat_A[886] * mat_B[705] +
//             mat_A[887] * mat_B[737] +
//             mat_A[888] * mat_B[769] +
//             mat_A[889] * mat_B[801] +
//             mat_A[890] * mat_B[833] +
//             mat_A[891] * mat_B[865] +
//             mat_A[892] * mat_B[897] +
//             mat_A[893] * mat_B[929] +
//             mat_A[894] * mat_B[961] +
//             mat_A[895] * mat_B[993];
//  mat_C[866] <= 
//             mat_A[864] * mat_B[2] +
//             mat_A[865] * mat_B[34] +
//             mat_A[866] * mat_B[66] +
//             mat_A[867] * mat_B[98] +
//             mat_A[868] * mat_B[130] +
//             mat_A[869] * mat_B[162] +
//             mat_A[870] * mat_B[194] +
//             mat_A[871] * mat_B[226] +
//             mat_A[872] * mat_B[258] +
//             mat_A[873] * mat_B[290] +
//             mat_A[874] * mat_B[322] +
//             mat_A[875] * mat_B[354] +
//             mat_A[876] * mat_B[386] +
//             mat_A[877] * mat_B[418] +
//             mat_A[878] * mat_B[450] +
//             mat_A[879] * mat_B[482] +
//             mat_A[880] * mat_B[514] +
//             mat_A[881] * mat_B[546] +
//             mat_A[882] * mat_B[578] +
//             mat_A[883] * mat_B[610] +
//             mat_A[884] * mat_B[642] +
//             mat_A[885] * mat_B[674] +
//             mat_A[886] * mat_B[706] +
//             mat_A[887] * mat_B[738] +
//             mat_A[888] * mat_B[770] +
//             mat_A[889] * mat_B[802] +
//             mat_A[890] * mat_B[834] +
//             mat_A[891] * mat_B[866] +
//             mat_A[892] * mat_B[898] +
//             mat_A[893] * mat_B[930] +
//             mat_A[894] * mat_B[962] +
//             mat_A[895] * mat_B[994];
//  mat_C[867] <= 
//             mat_A[864] * mat_B[3] +
//             mat_A[865] * mat_B[35] +
//             mat_A[866] * mat_B[67] +
//             mat_A[867] * mat_B[99] +
//             mat_A[868] * mat_B[131] +
//             mat_A[869] * mat_B[163] +
//             mat_A[870] * mat_B[195] +
//             mat_A[871] * mat_B[227] +
//             mat_A[872] * mat_B[259] +
//             mat_A[873] * mat_B[291] +
//             mat_A[874] * mat_B[323] +
//             mat_A[875] * mat_B[355] +
//             mat_A[876] * mat_B[387] +
//             mat_A[877] * mat_B[419] +
//             mat_A[878] * mat_B[451] +
//             mat_A[879] * mat_B[483] +
//             mat_A[880] * mat_B[515] +
//             mat_A[881] * mat_B[547] +
//             mat_A[882] * mat_B[579] +
//             mat_A[883] * mat_B[611] +
//             mat_A[884] * mat_B[643] +
//             mat_A[885] * mat_B[675] +
//             mat_A[886] * mat_B[707] +
//             mat_A[887] * mat_B[739] +
//             mat_A[888] * mat_B[771] +
//             mat_A[889] * mat_B[803] +
//             mat_A[890] * mat_B[835] +
//             mat_A[891] * mat_B[867] +
//             mat_A[892] * mat_B[899] +
//             mat_A[893] * mat_B[931] +
//             mat_A[894] * mat_B[963] +
//             mat_A[895] * mat_B[995];
//  mat_C[868] <= 
//             mat_A[864] * mat_B[4] +
//             mat_A[865] * mat_B[36] +
//             mat_A[866] * mat_B[68] +
//             mat_A[867] * mat_B[100] +
//             mat_A[868] * mat_B[132] +
//             mat_A[869] * mat_B[164] +
//             mat_A[870] * mat_B[196] +
//             mat_A[871] * mat_B[228] +
//             mat_A[872] * mat_B[260] +
//             mat_A[873] * mat_B[292] +
//             mat_A[874] * mat_B[324] +
//             mat_A[875] * mat_B[356] +
//             mat_A[876] * mat_B[388] +
//             mat_A[877] * mat_B[420] +
//             mat_A[878] * mat_B[452] +
//             mat_A[879] * mat_B[484] +
//             mat_A[880] * mat_B[516] +
//             mat_A[881] * mat_B[548] +
//             mat_A[882] * mat_B[580] +
//             mat_A[883] * mat_B[612] +
//             mat_A[884] * mat_B[644] +
//             mat_A[885] * mat_B[676] +
//             mat_A[886] * mat_B[708] +
//             mat_A[887] * mat_B[740] +
//             mat_A[888] * mat_B[772] +
//             mat_A[889] * mat_B[804] +
//             mat_A[890] * mat_B[836] +
//             mat_A[891] * mat_B[868] +
//             mat_A[892] * mat_B[900] +
//             mat_A[893] * mat_B[932] +
//             mat_A[894] * mat_B[964] +
//             mat_A[895] * mat_B[996];
//  mat_C[869] <= 
//             mat_A[864] * mat_B[5] +
//             mat_A[865] * mat_B[37] +
//             mat_A[866] * mat_B[69] +
//             mat_A[867] * mat_B[101] +
//             mat_A[868] * mat_B[133] +
//             mat_A[869] * mat_B[165] +
//             mat_A[870] * mat_B[197] +
//             mat_A[871] * mat_B[229] +
//             mat_A[872] * mat_B[261] +
//             mat_A[873] * mat_B[293] +
//             mat_A[874] * mat_B[325] +
//             mat_A[875] * mat_B[357] +
//             mat_A[876] * mat_B[389] +
//             mat_A[877] * mat_B[421] +
//             mat_A[878] * mat_B[453] +
//             mat_A[879] * mat_B[485] +
//             mat_A[880] * mat_B[517] +
//             mat_A[881] * mat_B[549] +
//             mat_A[882] * mat_B[581] +
//             mat_A[883] * mat_B[613] +
//             mat_A[884] * mat_B[645] +
//             mat_A[885] * mat_B[677] +
//             mat_A[886] * mat_B[709] +
//             mat_A[887] * mat_B[741] +
//             mat_A[888] * mat_B[773] +
//             mat_A[889] * mat_B[805] +
//             mat_A[890] * mat_B[837] +
//             mat_A[891] * mat_B[869] +
//             mat_A[892] * mat_B[901] +
//             mat_A[893] * mat_B[933] +
//             mat_A[894] * mat_B[965] +
//             mat_A[895] * mat_B[997];
//  mat_C[870] <= 
//             mat_A[864] * mat_B[6] +
//             mat_A[865] * mat_B[38] +
//             mat_A[866] * mat_B[70] +
//             mat_A[867] * mat_B[102] +
//             mat_A[868] * mat_B[134] +
//             mat_A[869] * mat_B[166] +
//             mat_A[870] * mat_B[198] +
//             mat_A[871] * mat_B[230] +
//             mat_A[872] * mat_B[262] +
//             mat_A[873] * mat_B[294] +
//             mat_A[874] * mat_B[326] +
//             mat_A[875] * mat_B[358] +
//             mat_A[876] * mat_B[390] +
//             mat_A[877] * mat_B[422] +
//             mat_A[878] * mat_B[454] +
//             mat_A[879] * mat_B[486] +
//             mat_A[880] * mat_B[518] +
//             mat_A[881] * mat_B[550] +
//             mat_A[882] * mat_B[582] +
//             mat_A[883] * mat_B[614] +
//             mat_A[884] * mat_B[646] +
//             mat_A[885] * mat_B[678] +
//             mat_A[886] * mat_B[710] +
//             mat_A[887] * mat_B[742] +
//             mat_A[888] * mat_B[774] +
//             mat_A[889] * mat_B[806] +
//             mat_A[890] * mat_B[838] +
//             mat_A[891] * mat_B[870] +
//             mat_A[892] * mat_B[902] +
//             mat_A[893] * mat_B[934] +
//             mat_A[894] * mat_B[966] +
//             mat_A[895] * mat_B[998];
//  mat_C[871] <= 
//             mat_A[864] * mat_B[7] +
//             mat_A[865] * mat_B[39] +
//             mat_A[866] * mat_B[71] +
//             mat_A[867] * mat_B[103] +
//             mat_A[868] * mat_B[135] +
//             mat_A[869] * mat_B[167] +
//             mat_A[870] * mat_B[199] +
//             mat_A[871] * mat_B[231] +
//             mat_A[872] * mat_B[263] +
//             mat_A[873] * mat_B[295] +
//             mat_A[874] * mat_B[327] +
//             mat_A[875] * mat_B[359] +
//             mat_A[876] * mat_B[391] +
//             mat_A[877] * mat_B[423] +
//             mat_A[878] * mat_B[455] +
//             mat_A[879] * mat_B[487] +
//             mat_A[880] * mat_B[519] +
//             mat_A[881] * mat_B[551] +
//             mat_A[882] * mat_B[583] +
//             mat_A[883] * mat_B[615] +
//             mat_A[884] * mat_B[647] +
//             mat_A[885] * mat_B[679] +
//             mat_A[886] * mat_B[711] +
//             mat_A[887] * mat_B[743] +
//             mat_A[888] * mat_B[775] +
//             mat_A[889] * mat_B[807] +
//             mat_A[890] * mat_B[839] +
//             mat_A[891] * mat_B[871] +
//             mat_A[892] * mat_B[903] +
//             mat_A[893] * mat_B[935] +
//             mat_A[894] * mat_B[967] +
//             mat_A[895] * mat_B[999];
//  mat_C[872] <= 
//             mat_A[864] * mat_B[8] +
//             mat_A[865] * mat_B[40] +
//             mat_A[866] * mat_B[72] +
//             mat_A[867] * mat_B[104] +
//             mat_A[868] * mat_B[136] +
//             mat_A[869] * mat_B[168] +
//             mat_A[870] * mat_B[200] +
//             mat_A[871] * mat_B[232] +
//             mat_A[872] * mat_B[264] +
//             mat_A[873] * mat_B[296] +
//             mat_A[874] * mat_B[328] +
//             mat_A[875] * mat_B[360] +
//             mat_A[876] * mat_B[392] +
//             mat_A[877] * mat_B[424] +
//             mat_A[878] * mat_B[456] +
//             mat_A[879] * mat_B[488] +
//             mat_A[880] * mat_B[520] +
//             mat_A[881] * mat_B[552] +
//             mat_A[882] * mat_B[584] +
//             mat_A[883] * mat_B[616] +
//             mat_A[884] * mat_B[648] +
//             mat_A[885] * mat_B[680] +
//             mat_A[886] * mat_B[712] +
//             mat_A[887] * mat_B[744] +
//             mat_A[888] * mat_B[776] +
//             mat_A[889] * mat_B[808] +
//             mat_A[890] * mat_B[840] +
//             mat_A[891] * mat_B[872] +
//             mat_A[892] * mat_B[904] +
//             mat_A[893] * mat_B[936] +
//             mat_A[894] * mat_B[968] +
//             mat_A[895] * mat_B[1000];
//  mat_C[873] <= 
//             mat_A[864] * mat_B[9] +
//             mat_A[865] * mat_B[41] +
//             mat_A[866] * mat_B[73] +
//             mat_A[867] * mat_B[105] +
//             mat_A[868] * mat_B[137] +
//             mat_A[869] * mat_B[169] +
//             mat_A[870] * mat_B[201] +
//             mat_A[871] * mat_B[233] +
//             mat_A[872] * mat_B[265] +
//             mat_A[873] * mat_B[297] +
//             mat_A[874] * mat_B[329] +
//             mat_A[875] * mat_B[361] +
//             mat_A[876] * mat_B[393] +
//             mat_A[877] * mat_B[425] +
//             mat_A[878] * mat_B[457] +
//             mat_A[879] * mat_B[489] +
//             mat_A[880] * mat_B[521] +
//             mat_A[881] * mat_B[553] +
//             mat_A[882] * mat_B[585] +
//             mat_A[883] * mat_B[617] +
//             mat_A[884] * mat_B[649] +
//             mat_A[885] * mat_B[681] +
//             mat_A[886] * mat_B[713] +
//             mat_A[887] * mat_B[745] +
//             mat_A[888] * mat_B[777] +
//             mat_A[889] * mat_B[809] +
//             mat_A[890] * mat_B[841] +
//             mat_A[891] * mat_B[873] +
//             mat_A[892] * mat_B[905] +
//             mat_A[893] * mat_B[937] +
//             mat_A[894] * mat_B[969] +
//             mat_A[895] * mat_B[1001];
//  mat_C[874] <= 
//             mat_A[864] * mat_B[10] +
//             mat_A[865] * mat_B[42] +
//             mat_A[866] * mat_B[74] +
//             mat_A[867] * mat_B[106] +
//             mat_A[868] * mat_B[138] +
//             mat_A[869] * mat_B[170] +
//             mat_A[870] * mat_B[202] +
//             mat_A[871] * mat_B[234] +
//             mat_A[872] * mat_B[266] +
//             mat_A[873] * mat_B[298] +
//             mat_A[874] * mat_B[330] +
//             mat_A[875] * mat_B[362] +
//             mat_A[876] * mat_B[394] +
//             mat_A[877] * mat_B[426] +
//             mat_A[878] * mat_B[458] +
//             mat_A[879] * mat_B[490] +
//             mat_A[880] * mat_B[522] +
//             mat_A[881] * mat_B[554] +
//             mat_A[882] * mat_B[586] +
//             mat_A[883] * mat_B[618] +
//             mat_A[884] * mat_B[650] +
//             mat_A[885] * mat_B[682] +
//             mat_A[886] * mat_B[714] +
//             mat_A[887] * mat_B[746] +
//             mat_A[888] * mat_B[778] +
//             mat_A[889] * mat_B[810] +
//             mat_A[890] * mat_B[842] +
//             mat_A[891] * mat_B[874] +
//             mat_A[892] * mat_B[906] +
//             mat_A[893] * mat_B[938] +
//             mat_A[894] * mat_B[970] +
//             mat_A[895] * mat_B[1002];
//  mat_C[875] <= 
//             mat_A[864] * mat_B[11] +
//             mat_A[865] * mat_B[43] +
//             mat_A[866] * mat_B[75] +
//             mat_A[867] * mat_B[107] +
//             mat_A[868] * mat_B[139] +
//             mat_A[869] * mat_B[171] +
//             mat_A[870] * mat_B[203] +
//             mat_A[871] * mat_B[235] +
//             mat_A[872] * mat_B[267] +
//             mat_A[873] * mat_B[299] +
//             mat_A[874] * mat_B[331] +
//             mat_A[875] * mat_B[363] +
//             mat_A[876] * mat_B[395] +
//             mat_A[877] * mat_B[427] +
//             mat_A[878] * mat_B[459] +
//             mat_A[879] * mat_B[491] +
//             mat_A[880] * mat_B[523] +
//             mat_A[881] * mat_B[555] +
//             mat_A[882] * mat_B[587] +
//             mat_A[883] * mat_B[619] +
//             mat_A[884] * mat_B[651] +
//             mat_A[885] * mat_B[683] +
//             mat_A[886] * mat_B[715] +
//             mat_A[887] * mat_B[747] +
//             mat_A[888] * mat_B[779] +
//             mat_A[889] * mat_B[811] +
//             mat_A[890] * mat_B[843] +
//             mat_A[891] * mat_B[875] +
//             mat_A[892] * mat_B[907] +
//             mat_A[893] * mat_B[939] +
//             mat_A[894] * mat_B[971] +
//             mat_A[895] * mat_B[1003];
//  mat_C[876] <= 
//             mat_A[864] * mat_B[12] +
//             mat_A[865] * mat_B[44] +
//             mat_A[866] * mat_B[76] +
//             mat_A[867] * mat_B[108] +
//             mat_A[868] * mat_B[140] +
//             mat_A[869] * mat_B[172] +
//             mat_A[870] * mat_B[204] +
//             mat_A[871] * mat_B[236] +
//             mat_A[872] * mat_B[268] +
//             mat_A[873] * mat_B[300] +
//             mat_A[874] * mat_B[332] +
//             mat_A[875] * mat_B[364] +
//             mat_A[876] * mat_B[396] +
//             mat_A[877] * mat_B[428] +
//             mat_A[878] * mat_B[460] +
//             mat_A[879] * mat_B[492] +
//             mat_A[880] * mat_B[524] +
//             mat_A[881] * mat_B[556] +
//             mat_A[882] * mat_B[588] +
//             mat_A[883] * mat_B[620] +
//             mat_A[884] * mat_B[652] +
//             mat_A[885] * mat_B[684] +
//             mat_A[886] * mat_B[716] +
//             mat_A[887] * mat_B[748] +
//             mat_A[888] * mat_B[780] +
//             mat_A[889] * mat_B[812] +
//             mat_A[890] * mat_B[844] +
//             mat_A[891] * mat_B[876] +
//             mat_A[892] * mat_B[908] +
//             mat_A[893] * mat_B[940] +
//             mat_A[894] * mat_B[972] +
//             mat_A[895] * mat_B[1004];
//  mat_C[877] <= 
//             mat_A[864] * mat_B[13] +
//             mat_A[865] * mat_B[45] +
//             mat_A[866] * mat_B[77] +
//             mat_A[867] * mat_B[109] +
//             mat_A[868] * mat_B[141] +
//             mat_A[869] * mat_B[173] +
//             mat_A[870] * mat_B[205] +
//             mat_A[871] * mat_B[237] +
//             mat_A[872] * mat_B[269] +
//             mat_A[873] * mat_B[301] +
//             mat_A[874] * mat_B[333] +
//             mat_A[875] * mat_B[365] +
//             mat_A[876] * mat_B[397] +
//             mat_A[877] * mat_B[429] +
//             mat_A[878] * mat_B[461] +
//             mat_A[879] * mat_B[493] +
//             mat_A[880] * mat_B[525] +
//             mat_A[881] * mat_B[557] +
//             mat_A[882] * mat_B[589] +
//             mat_A[883] * mat_B[621] +
//             mat_A[884] * mat_B[653] +
//             mat_A[885] * mat_B[685] +
//             mat_A[886] * mat_B[717] +
//             mat_A[887] * mat_B[749] +
//             mat_A[888] * mat_B[781] +
//             mat_A[889] * mat_B[813] +
//             mat_A[890] * mat_B[845] +
//             mat_A[891] * mat_B[877] +
//             mat_A[892] * mat_B[909] +
//             mat_A[893] * mat_B[941] +
//             mat_A[894] * mat_B[973] +
//             mat_A[895] * mat_B[1005];
//  mat_C[878] <= 
//             mat_A[864] * mat_B[14] +
//             mat_A[865] * mat_B[46] +
//             mat_A[866] * mat_B[78] +
//             mat_A[867] * mat_B[110] +
//             mat_A[868] * mat_B[142] +
//             mat_A[869] * mat_B[174] +
//             mat_A[870] * mat_B[206] +
//             mat_A[871] * mat_B[238] +
//             mat_A[872] * mat_B[270] +
//             mat_A[873] * mat_B[302] +
//             mat_A[874] * mat_B[334] +
//             mat_A[875] * mat_B[366] +
//             mat_A[876] * mat_B[398] +
//             mat_A[877] * mat_B[430] +
//             mat_A[878] * mat_B[462] +
//             mat_A[879] * mat_B[494] +
//             mat_A[880] * mat_B[526] +
//             mat_A[881] * mat_B[558] +
//             mat_A[882] * mat_B[590] +
//             mat_A[883] * mat_B[622] +
//             mat_A[884] * mat_B[654] +
//             mat_A[885] * mat_B[686] +
//             mat_A[886] * mat_B[718] +
//             mat_A[887] * mat_B[750] +
//             mat_A[888] * mat_B[782] +
//             mat_A[889] * mat_B[814] +
//             mat_A[890] * mat_B[846] +
//             mat_A[891] * mat_B[878] +
//             mat_A[892] * mat_B[910] +
//             mat_A[893] * mat_B[942] +
//             mat_A[894] * mat_B[974] +
//             mat_A[895] * mat_B[1006];
//  mat_C[879] <= 
//             mat_A[864] * mat_B[15] +
//             mat_A[865] * mat_B[47] +
//             mat_A[866] * mat_B[79] +
//             mat_A[867] * mat_B[111] +
//             mat_A[868] * mat_B[143] +
//             mat_A[869] * mat_B[175] +
//             mat_A[870] * mat_B[207] +
//             mat_A[871] * mat_B[239] +
//             mat_A[872] * mat_B[271] +
//             mat_A[873] * mat_B[303] +
//             mat_A[874] * mat_B[335] +
//             mat_A[875] * mat_B[367] +
//             mat_A[876] * mat_B[399] +
//             mat_A[877] * mat_B[431] +
//             mat_A[878] * mat_B[463] +
//             mat_A[879] * mat_B[495] +
//             mat_A[880] * mat_B[527] +
//             mat_A[881] * mat_B[559] +
//             mat_A[882] * mat_B[591] +
//             mat_A[883] * mat_B[623] +
//             mat_A[884] * mat_B[655] +
//             mat_A[885] * mat_B[687] +
//             mat_A[886] * mat_B[719] +
//             mat_A[887] * mat_B[751] +
//             mat_A[888] * mat_B[783] +
//             mat_A[889] * mat_B[815] +
//             mat_A[890] * mat_B[847] +
//             mat_A[891] * mat_B[879] +
//             mat_A[892] * mat_B[911] +
//             mat_A[893] * mat_B[943] +
//             mat_A[894] * mat_B[975] +
//             mat_A[895] * mat_B[1007];
//  mat_C[880] <= 
//             mat_A[864] * mat_B[16] +
//             mat_A[865] * mat_B[48] +
//             mat_A[866] * mat_B[80] +
//             mat_A[867] * mat_B[112] +
//             mat_A[868] * mat_B[144] +
//             mat_A[869] * mat_B[176] +
//             mat_A[870] * mat_B[208] +
//             mat_A[871] * mat_B[240] +
//             mat_A[872] * mat_B[272] +
//             mat_A[873] * mat_B[304] +
//             mat_A[874] * mat_B[336] +
//             mat_A[875] * mat_B[368] +
//             mat_A[876] * mat_B[400] +
//             mat_A[877] * mat_B[432] +
//             mat_A[878] * mat_B[464] +
//             mat_A[879] * mat_B[496] +
//             mat_A[880] * mat_B[528] +
//             mat_A[881] * mat_B[560] +
//             mat_A[882] * mat_B[592] +
//             mat_A[883] * mat_B[624] +
//             mat_A[884] * mat_B[656] +
//             mat_A[885] * mat_B[688] +
//             mat_A[886] * mat_B[720] +
//             mat_A[887] * mat_B[752] +
//             mat_A[888] * mat_B[784] +
//             mat_A[889] * mat_B[816] +
//             mat_A[890] * mat_B[848] +
//             mat_A[891] * mat_B[880] +
//             mat_A[892] * mat_B[912] +
//             mat_A[893] * mat_B[944] +
//             mat_A[894] * mat_B[976] +
//             mat_A[895] * mat_B[1008];
//  mat_C[881] <= 
//             mat_A[864] * mat_B[17] +
//             mat_A[865] * mat_B[49] +
//             mat_A[866] * mat_B[81] +
//             mat_A[867] * mat_B[113] +
//             mat_A[868] * mat_B[145] +
//             mat_A[869] * mat_B[177] +
//             mat_A[870] * mat_B[209] +
//             mat_A[871] * mat_B[241] +
//             mat_A[872] * mat_B[273] +
//             mat_A[873] * mat_B[305] +
//             mat_A[874] * mat_B[337] +
//             mat_A[875] * mat_B[369] +
//             mat_A[876] * mat_B[401] +
//             mat_A[877] * mat_B[433] +
//             mat_A[878] * mat_B[465] +
//             mat_A[879] * mat_B[497] +
//             mat_A[880] * mat_B[529] +
//             mat_A[881] * mat_B[561] +
//             mat_A[882] * mat_B[593] +
//             mat_A[883] * mat_B[625] +
//             mat_A[884] * mat_B[657] +
//             mat_A[885] * mat_B[689] +
//             mat_A[886] * mat_B[721] +
//             mat_A[887] * mat_B[753] +
//             mat_A[888] * mat_B[785] +
//             mat_A[889] * mat_B[817] +
//             mat_A[890] * mat_B[849] +
//             mat_A[891] * mat_B[881] +
//             mat_A[892] * mat_B[913] +
//             mat_A[893] * mat_B[945] +
//             mat_A[894] * mat_B[977] +
//             mat_A[895] * mat_B[1009];
//  mat_C[882] <= 
//             mat_A[864] * mat_B[18] +
//             mat_A[865] * mat_B[50] +
//             mat_A[866] * mat_B[82] +
//             mat_A[867] * mat_B[114] +
//             mat_A[868] * mat_B[146] +
//             mat_A[869] * mat_B[178] +
//             mat_A[870] * mat_B[210] +
//             mat_A[871] * mat_B[242] +
//             mat_A[872] * mat_B[274] +
//             mat_A[873] * mat_B[306] +
//             mat_A[874] * mat_B[338] +
//             mat_A[875] * mat_B[370] +
//             mat_A[876] * mat_B[402] +
//             mat_A[877] * mat_B[434] +
//             mat_A[878] * mat_B[466] +
//             mat_A[879] * mat_B[498] +
//             mat_A[880] * mat_B[530] +
//             mat_A[881] * mat_B[562] +
//             mat_A[882] * mat_B[594] +
//             mat_A[883] * mat_B[626] +
//             mat_A[884] * mat_B[658] +
//             mat_A[885] * mat_B[690] +
//             mat_A[886] * mat_B[722] +
//             mat_A[887] * mat_B[754] +
//             mat_A[888] * mat_B[786] +
//             mat_A[889] * mat_B[818] +
//             mat_A[890] * mat_B[850] +
//             mat_A[891] * mat_B[882] +
//             mat_A[892] * mat_B[914] +
//             mat_A[893] * mat_B[946] +
//             mat_A[894] * mat_B[978] +
//             mat_A[895] * mat_B[1010];
//  mat_C[883] <= 
//             mat_A[864] * mat_B[19] +
//             mat_A[865] * mat_B[51] +
//             mat_A[866] * mat_B[83] +
//             mat_A[867] * mat_B[115] +
//             mat_A[868] * mat_B[147] +
//             mat_A[869] * mat_B[179] +
//             mat_A[870] * mat_B[211] +
//             mat_A[871] * mat_B[243] +
//             mat_A[872] * mat_B[275] +
//             mat_A[873] * mat_B[307] +
//             mat_A[874] * mat_B[339] +
//             mat_A[875] * mat_B[371] +
//             mat_A[876] * mat_B[403] +
//             mat_A[877] * mat_B[435] +
//             mat_A[878] * mat_B[467] +
//             mat_A[879] * mat_B[499] +
//             mat_A[880] * mat_B[531] +
//             mat_A[881] * mat_B[563] +
//             mat_A[882] * mat_B[595] +
//             mat_A[883] * mat_B[627] +
//             mat_A[884] * mat_B[659] +
//             mat_A[885] * mat_B[691] +
//             mat_A[886] * mat_B[723] +
//             mat_A[887] * mat_B[755] +
//             mat_A[888] * mat_B[787] +
//             mat_A[889] * mat_B[819] +
//             mat_A[890] * mat_B[851] +
//             mat_A[891] * mat_B[883] +
//             mat_A[892] * mat_B[915] +
//             mat_A[893] * mat_B[947] +
//             mat_A[894] * mat_B[979] +
//             mat_A[895] * mat_B[1011];
//  mat_C[884] <= 
//             mat_A[864] * mat_B[20] +
//             mat_A[865] * mat_B[52] +
//             mat_A[866] * mat_B[84] +
//             mat_A[867] * mat_B[116] +
//             mat_A[868] * mat_B[148] +
//             mat_A[869] * mat_B[180] +
//             mat_A[870] * mat_B[212] +
//             mat_A[871] * mat_B[244] +
//             mat_A[872] * mat_B[276] +
//             mat_A[873] * mat_B[308] +
//             mat_A[874] * mat_B[340] +
//             mat_A[875] * mat_B[372] +
//             mat_A[876] * mat_B[404] +
//             mat_A[877] * mat_B[436] +
//             mat_A[878] * mat_B[468] +
//             mat_A[879] * mat_B[500] +
//             mat_A[880] * mat_B[532] +
//             mat_A[881] * mat_B[564] +
//             mat_A[882] * mat_B[596] +
//             mat_A[883] * mat_B[628] +
//             mat_A[884] * mat_B[660] +
//             mat_A[885] * mat_B[692] +
//             mat_A[886] * mat_B[724] +
//             mat_A[887] * mat_B[756] +
//             mat_A[888] * mat_B[788] +
//             mat_A[889] * mat_B[820] +
//             mat_A[890] * mat_B[852] +
//             mat_A[891] * mat_B[884] +
//             mat_A[892] * mat_B[916] +
//             mat_A[893] * mat_B[948] +
//             mat_A[894] * mat_B[980] +
//             mat_A[895] * mat_B[1012];
//  mat_C[885] <= 
//             mat_A[864] * mat_B[21] +
//             mat_A[865] * mat_B[53] +
//             mat_A[866] * mat_B[85] +
//             mat_A[867] * mat_B[117] +
//             mat_A[868] * mat_B[149] +
//             mat_A[869] * mat_B[181] +
//             mat_A[870] * mat_B[213] +
//             mat_A[871] * mat_B[245] +
//             mat_A[872] * mat_B[277] +
//             mat_A[873] * mat_B[309] +
//             mat_A[874] * mat_B[341] +
//             mat_A[875] * mat_B[373] +
//             mat_A[876] * mat_B[405] +
//             mat_A[877] * mat_B[437] +
//             mat_A[878] * mat_B[469] +
//             mat_A[879] * mat_B[501] +
//             mat_A[880] * mat_B[533] +
//             mat_A[881] * mat_B[565] +
//             mat_A[882] * mat_B[597] +
//             mat_A[883] * mat_B[629] +
//             mat_A[884] * mat_B[661] +
//             mat_A[885] * mat_B[693] +
//             mat_A[886] * mat_B[725] +
//             mat_A[887] * mat_B[757] +
//             mat_A[888] * mat_B[789] +
//             mat_A[889] * mat_B[821] +
//             mat_A[890] * mat_B[853] +
//             mat_A[891] * mat_B[885] +
//             mat_A[892] * mat_B[917] +
//             mat_A[893] * mat_B[949] +
//             mat_A[894] * mat_B[981] +
//             mat_A[895] * mat_B[1013];
//  mat_C[886] <= 
//             mat_A[864] * mat_B[22] +
//             mat_A[865] * mat_B[54] +
//             mat_A[866] * mat_B[86] +
//             mat_A[867] * mat_B[118] +
//             mat_A[868] * mat_B[150] +
//             mat_A[869] * mat_B[182] +
//             mat_A[870] * mat_B[214] +
//             mat_A[871] * mat_B[246] +
//             mat_A[872] * mat_B[278] +
//             mat_A[873] * mat_B[310] +
//             mat_A[874] * mat_B[342] +
//             mat_A[875] * mat_B[374] +
//             mat_A[876] * mat_B[406] +
//             mat_A[877] * mat_B[438] +
//             mat_A[878] * mat_B[470] +
//             mat_A[879] * mat_B[502] +
//             mat_A[880] * mat_B[534] +
//             mat_A[881] * mat_B[566] +
//             mat_A[882] * mat_B[598] +
//             mat_A[883] * mat_B[630] +
//             mat_A[884] * mat_B[662] +
//             mat_A[885] * mat_B[694] +
//             mat_A[886] * mat_B[726] +
//             mat_A[887] * mat_B[758] +
//             mat_A[888] * mat_B[790] +
//             mat_A[889] * mat_B[822] +
//             mat_A[890] * mat_B[854] +
//             mat_A[891] * mat_B[886] +
//             mat_A[892] * mat_B[918] +
//             mat_A[893] * mat_B[950] +
//             mat_A[894] * mat_B[982] +
//             mat_A[895] * mat_B[1014];
//  mat_C[887] <= 
//             mat_A[864] * mat_B[23] +
//             mat_A[865] * mat_B[55] +
//             mat_A[866] * mat_B[87] +
//             mat_A[867] * mat_B[119] +
//             mat_A[868] * mat_B[151] +
//             mat_A[869] * mat_B[183] +
//             mat_A[870] * mat_B[215] +
//             mat_A[871] * mat_B[247] +
//             mat_A[872] * mat_B[279] +
//             mat_A[873] * mat_B[311] +
//             mat_A[874] * mat_B[343] +
//             mat_A[875] * mat_B[375] +
//             mat_A[876] * mat_B[407] +
//             mat_A[877] * mat_B[439] +
//             mat_A[878] * mat_B[471] +
//             mat_A[879] * mat_B[503] +
//             mat_A[880] * mat_B[535] +
//             mat_A[881] * mat_B[567] +
//             mat_A[882] * mat_B[599] +
//             mat_A[883] * mat_B[631] +
//             mat_A[884] * mat_B[663] +
//             mat_A[885] * mat_B[695] +
//             mat_A[886] * mat_B[727] +
//             mat_A[887] * mat_B[759] +
//             mat_A[888] * mat_B[791] +
//             mat_A[889] * mat_B[823] +
//             mat_A[890] * mat_B[855] +
//             mat_A[891] * mat_B[887] +
//             mat_A[892] * mat_B[919] +
//             mat_A[893] * mat_B[951] +
//             mat_A[894] * mat_B[983] +
//             mat_A[895] * mat_B[1015];
//  mat_C[888] <= 
//             mat_A[864] * mat_B[24] +
//             mat_A[865] * mat_B[56] +
//             mat_A[866] * mat_B[88] +
//             mat_A[867] * mat_B[120] +
//             mat_A[868] * mat_B[152] +
//             mat_A[869] * mat_B[184] +
//             mat_A[870] * mat_B[216] +
//             mat_A[871] * mat_B[248] +
//             mat_A[872] * mat_B[280] +
//             mat_A[873] * mat_B[312] +
//             mat_A[874] * mat_B[344] +
//             mat_A[875] * mat_B[376] +
//             mat_A[876] * mat_B[408] +
//             mat_A[877] * mat_B[440] +
//             mat_A[878] * mat_B[472] +
//             mat_A[879] * mat_B[504] +
//             mat_A[880] * mat_B[536] +
//             mat_A[881] * mat_B[568] +
//             mat_A[882] * mat_B[600] +
//             mat_A[883] * mat_B[632] +
//             mat_A[884] * mat_B[664] +
//             mat_A[885] * mat_B[696] +
//             mat_A[886] * mat_B[728] +
//             mat_A[887] * mat_B[760] +
//             mat_A[888] * mat_B[792] +
//             mat_A[889] * mat_B[824] +
//             mat_A[890] * mat_B[856] +
//             mat_A[891] * mat_B[888] +
//             mat_A[892] * mat_B[920] +
//             mat_A[893] * mat_B[952] +
//             mat_A[894] * mat_B[984] +
//             mat_A[895] * mat_B[1016];
//  mat_C[889] <= 
//             mat_A[864] * mat_B[25] +
//             mat_A[865] * mat_B[57] +
//             mat_A[866] * mat_B[89] +
//             mat_A[867] * mat_B[121] +
//             mat_A[868] * mat_B[153] +
//             mat_A[869] * mat_B[185] +
//             mat_A[870] * mat_B[217] +
//             mat_A[871] * mat_B[249] +
//             mat_A[872] * mat_B[281] +
//             mat_A[873] * mat_B[313] +
//             mat_A[874] * mat_B[345] +
//             mat_A[875] * mat_B[377] +
//             mat_A[876] * mat_B[409] +
//             mat_A[877] * mat_B[441] +
//             mat_A[878] * mat_B[473] +
//             mat_A[879] * mat_B[505] +
//             mat_A[880] * mat_B[537] +
//             mat_A[881] * mat_B[569] +
//             mat_A[882] * mat_B[601] +
//             mat_A[883] * mat_B[633] +
//             mat_A[884] * mat_B[665] +
//             mat_A[885] * mat_B[697] +
//             mat_A[886] * mat_B[729] +
//             mat_A[887] * mat_B[761] +
//             mat_A[888] * mat_B[793] +
//             mat_A[889] * mat_B[825] +
//             mat_A[890] * mat_B[857] +
//             mat_A[891] * mat_B[889] +
//             mat_A[892] * mat_B[921] +
//             mat_A[893] * mat_B[953] +
//             mat_A[894] * mat_B[985] +
//             mat_A[895] * mat_B[1017];
//  mat_C[890] <= 
//             mat_A[864] * mat_B[26] +
//             mat_A[865] * mat_B[58] +
//             mat_A[866] * mat_B[90] +
//             mat_A[867] * mat_B[122] +
//             mat_A[868] * mat_B[154] +
//             mat_A[869] * mat_B[186] +
//             mat_A[870] * mat_B[218] +
//             mat_A[871] * mat_B[250] +
//             mat_A[872] * mat_B[282] +
//             mat_A[873] * mat_B[314] +
//             mat_A[874] * mat_B[346] +
//             mat_A[875] * mat_B[378] +
//             mat_A[876] * mat_B[410] +
//             mat_A[877] * mat_B[442] +
//             mat_A[878] * mat_B[474] +
//             mat_A[879] * mat_B[506] +
//             mat_A[880] * mat_B[538] +
//             mat_A[881] * mat_B[570] +
//             mat_A[882] * mat_B[602] +
//             mat_A[883] * mat_B[634] +
//             mat_A[884] * mat_B[666] +
//             mat_A[885] * mat_B[698] +
//             mat_A[886] * mat_B[730] +
//             mat_A[887] * mat_B[762] +
//             mat_A[888] * mat_B[794] +
//             mat_A[889] * mat_B[826] +
//             mat_A[890] * mat_B[858] +
//             mat_A[891] * mat_B[890] +
//             mat_A[892] * mat_B[922] +
//             mat_A[893] * mat_B[954] +
//             mat_A[894] * mat_B[986] +
//             mat_A[895] * mat_B[1018];
//  mat_C[891] <= 
//             mat_A[864] * mat_B[27] +
//             mat_A[865] * mat_B[59] +
//             mat_A[866] * mat_B[91] +
//             mat_A[867] * mat_B[123] +
//             mat_A[868] * mat_B[155] +
//             mat_A[869] * mat_B[187] +
//             mat_A[870] * mat_B[219] +
//             mat_A[871] * mat_B[251] +
//             mat_A[872] * mat_B[283] +
//             mat_A[873] * mat_B[315] +
//             mat_A[874] * mat_B[347] +
//             mat_A[875] * mat_B[379] +
//             mat_A[876] * mat_B[411] +
//             mat_A[877] * mat_B[443] +
//             mat_A[878] * mat_B[475] +
//             mat_A[879] * mat_B[507] +
//             mat_A[880] * mat_B[539] +
//             mat_A[881] * mat_B[571] +
//             mat_A[882] * mat_B[603] +
//             mat_A[883] * mat_B[635] +
//             mat_A[884] * mat_B[667] +
//             mat_A[885] * mat_B[699] +
//             mat_A[886] * mat_B[731] +
//             mat_A[887] * mat_B[763] +
//             mat_A[888] * mat_B[795] +
//             mat_A[889] * mat_B[827] +
//             mat_A[890] * mat_B[859] +
//             mat_A[891] * mat_B[891] +
//             mat_A[892] * mat_B[923] +
//             mat_A[893] * mat_B[955] +
//             mat_A[894] * mat_B[987] +
//             mat_A[895] * mat_B[1019];
//  mat_C[892] <= 
//             mat_A[864] * mat_B[28] +
//             mat_A[865] * mat_B[60] +
//             mat_A[866] * mat_B[92] +
//             mat_A[867] * mat_B[124] +
//             mat_A[868] * mat_B[156] +
//             mat_A[869] * mat_B[188] +
//             mat_A[870] * mat_B[220] +
//             mat_A[871] * mat_B[252] +
//             mat_A[872] * mat_B[284] +
//             mat_A[873] * mat_B[316] +
//             mat_A[874] * mat_B[348] +
//             mat_A[875] * mat_B[380] +
//             mat_A[876] * mat_B[412] +
//             mat_A[877] * mat_B[444] +
//             mat_A[878] * mat_B[476] +
//             mat_A[879] * mat_B[508] +
//             mat_A[880] * mat_B[540] +
//             mat_A[881] * mat_B[572] +
//             mat_A[882] * mat_B[604] +
//             mat_A[883] * mat_B[636] +
//             mat_A[884] * mat_B[668] +
//             mat_A[885] * mat_B[700] +
//             mat_A[886] * mat_B[732] +
//             mat_A[887] * mat_B[764] +
//             mat_A[888] * mat_B[796] +
//             mat_A[889] * mat_B[828] +
//             mat_A[890] * mat_B[860] +
//             mat_A[891] * mat_B[892] +
//             mat_A[892] * mat_B[924] +
//             mat_A[893] * mat_B[956] +
//             mat_A[894] * mat_B[988] +
//             mat_A[895] * mat_B[1020];
//  mat_C[893] <= 
//             mat_A[864] * mat_B[29] +
//             mat_A[865] * mat_B[61] +
//             mat_A[866] * mat_B[93] +
//             mat_A[867] * mat_B[125] +
//             mat_A[868] * mat_B[157] +
//             mat_A[869] * mat_B[189] +
//             mat_A[870] * mat_B[221] +
//             mat_A[871] * mat_B[253] +
//             mat_A[872] * mat_B[285] +
//             mat_A[873] * mat_B[317] +
//             mat_A[874] * mat_B[349] +
//             mat_A[875] * mat_B[381] +
//             mat_A[876] * mat_B[413] +
//             mat_A[877] * mat_B[445] +
//             mat_A[878] * mat_B[477] +
//             mat_A[879] * mat_B[509] +
//             mat_A[880] * mat_B[541] +
//             mat_A[881] * mat_B[573] +
//             mat_A[882] * mat_B[605] +
//             mat_A[883] * mat_B[637] +
//             mat_A[884] * mat_B[669] +
//             mat_A[885] * mat_B[701] +
//             mat_A[886] * mat_B[733] +
//             mat_A[887] * mat_B[765] +
//             mat_A[888] * mat_B[797] +
//             mat_A[889] * mat_B[829] +
//             mat_A[890] * mat_B[861] +
//             mat_A[891] * mat_B[893] +
//             mat_A[892] * mat_B[925] +
//             mat_A[893] * mat_B[957] +
//             mat_A[894] * mat_B[989] +
//             mat_A[895] * mat_B[1021];
//  mat_C[894] <= 
//             mat_A[864] * mat_B[30] +
//             mat_A[865] * mat_B[62] +
//             mat_A[866] * mat_B[94] +
//             mat_A[867] * mat_B[126] +
//             mat_A[868] * mat_B[158] +
//             mat_A[869] * mat_B[190] +
//             mat_A[870] * mat_B[222] +
//             mat_A[871] * mat_B[254] +
//             mat_A[872] * mat_B[286] +
//             mat_A[873] * mat_B[318] +
//             mat_A[874] * mat_B[350] +
//             mat_A[875] * mat_B[382] +
//             mat_A[876] * mat_B[414] +
//             mat_A[877] * mat_B[446] +
//             mat_A[878] * mat_B[478] +
//             mat_A[879] * mat_B[510] +
//             mat_A[880] * mat_B[542] +
//             mat_A[881] * mat_B[574] +
//             mat_A[882] * mat_B[606] +
//             mat_A[883] * mat_B[638] +
//             mat_A[884] * mat_B[670] +
//             mat_A[885] * mat_B[702] +
//             mat_A[886] * mat_B[734] +
//             mat_A[887] * mat_B[766] +
//             mat_A[888] * mat_B[798] +
//             mat_A[889] * mat_B[830] +
//             mat_A[890] * mat_B[862] +
//             mat_A[891] * mat_B[894] +
//             mat_A[892] * mat_B[926] +
//             mat_A[893] * mat_B[958] +
//             mat_A[894] * mat_B[990] +
//             mat_A[895] * mat_B[1022];
//  mat_C[895] <= 
//             mat_A[864] * mat_B[31] +
//             mat_A[865] * mat_B[63] +
//             mat_A[866] * mat_B[95] +
//             mat_A[867] * mat_B[127] +
//             mat_A[868] * mat_B[159] +
//             mat_A[869] * mat_B[191] +
//             mat_A[870] * mat_B[223] +
//             mat_A[871] * mat_B[255] +
//             mat_A[872] * mat_B[287] +
//             mat_A[873] * mat_B[319] +
//             mat_A[874] * mat_B[351] +
//             mat_A[875] * mat_B[383] +
//             mat_A[876] * mat_B[415] +
//             mat_A[877] * mat_B[447] +
//             mat_A[878] * mat_B[479] +
//             mat_A[879] * mat_B[511] +
//             mat_A[880] * mat_B[543] +
//             mat_A[881] * mat_B[575] +
//             mat_A[882] * mat_B[607] +
//             mat_A[883] * mat_B[639] +
//             mat_A[884] * mat_B[671] +
//             mat_A[885] * mat_B[703] +
//             mat_A[886] * mat_B[735] +
//             mat_A[887] * mat_B[767] +
//             mat_A[888] * mat_B[799] +
//             mat_A[889] * mat_B[831] +
//             mat_A[890] * mat_B[863] +
//             mat_A[891] * mat_B[895] +
//             mat_A[892] * mat_B[927] +
//             mat_A[893] * mat_B[959] +
//             mat_A[894] * mat_B[991] +
//             mat_A[895] * mat_B[1023];
//  mat_C[896] <= 
//             mat_A[896] * mat_B[0] +
//             mat_A[897] * mat_B[32] +
//             mat_A[898] * mat_B[64] +
//             mat_A[899] * mat_B[96] +
//             mat_A[900] * mat_B[128] +
//             mat_A[901] * mat_B[160] +
//             mat_A[902] * mat_B[192] +
//             mat_A[903] * mat_B[224] +
//             mat_A[904] * mat_B[256] +
//             mat_A[905] * mat_B[288] +
//             mat_A[906] * mat_B[320] +
//             mat_A[907] * mat_B[352] +
//             mat_A[908] * mat_B[384] +
//             mat_A[909] * mat_B[416] +
//             mat_A[910] * mat_B[448] +
//             mat_A[911] * mat_B[480] +
//             mat_A[912] * mat_B[512] +
//             mat_A[913] * mat_B[544] +
//             mat_A[914] * mat_B[576] +
//             mat_A[915] * mat_B[608] +
//             mat_A[916] * mat_B[640] +
//             mat_A[917] * mat_B[672] +
//             mat_A[918] * mat_B[704] +
//             mat_A[919] * mat_B[736] +
//             mat_A[920] * mat_B[768] +
//             mat_A[921] * mat_B[800] +
//             mat_A[922] * mat_B[832] +
//             mat_A[923] * mat_B[864] +
//             mat_A[924] * mat_B[896] +
//             mat_A[925] * mat_B[928] +
//             mat_A[926] * mat_B[960] +
//             mat_A[927] * mat_B[992];
//  mat_C[897] <= 
//             mat_A[896] * mat_B[1] +
//             mat_A[897] * mat_B[33] +
//             mat_A[898] * mat_B[65] +
//             mat_A[899] * mat_B[97] +
//             mat_A[900] * mat_B[129] +
//             mat_A[901] * mat_B[161] +
//             mat_A[902] * mat_B[193] +
//             mat_A[903] * mat_B[225] +
//             mat_A[904] * mat_B[257] +
//             mat_A[905] * mat_B[289] +
//             mat_A[906] * mat_B[321] +
//             mat_A[907] * mat_B[353] +
//             mat_A[908] * mat_B[385] +
//             mat_A[909] * mat_B[417] +
//             mat_A[910] * mat_B[449] +
//             mat_A[911] * mat_B[481] +
//             mat_A[912] * mat_B[513] +
//             mat_A[913] * mat_B[545] +
//             mat_A[914] * mat_B[577] +
//             mat_A[915] * mat_B[609] +
//             mat_A[916] * mat_B[641] +
//             mat_A[917] * mat_B[673] +
//             mat_A[918] * mat_B[705] +
//             mat_A[919] * mat_B[737] +
//             mat_A[920] * mat_B[769] +
//             mat_A[921] * mat_B[801] +
//             mat_A[922] * mat_B[833] +
//             mat_A[923] * mat_B[865] +
//             mat_A[924] * mat_B[897] +
//             mat_A[925] * mat_B[929] +
//             mat_A[926] * mat_B[961] +
//             mat_A[927] * mat_B[993];
//  mat_C[898] <= 
//             mat_A[896] * mat_B[2] +
//             mat_A[897] * mat_B[34] +
//             mat_A[898] * mat_B[66] +
//             mat_A[899] * mat_B[98] +
//             mat_A[900] * mat_B[130] +
//             mat_A[901] * mat_B[162] +
//             mat_A[902] * mat_B[194] +
//             mat_A[903] * mat_B[226] +
//             mat_A[904] * mat_B[258] +
//             mat_A[905] * mat_B[290] +
//             mat_A[906] * mat_B[322] +
//             mat_A[907] * mat_B[354] +
//             mat_A[908] * mat_B[386] +
//             mat_A[909] * mat_B[418] +
//             mat_A[910] * mat_B[450] +
//             mat_A[911] * mat_B[482] +
//             mat_A[912] * mat_B[514] +
//             mat_A[913] * mat_B[546] +
//             mat_A[914] * mat_B[578] +
//             mat_A[915] * mat_B[610] +
//             mat_A[916] * mat_B[642] +
//             mat_A[917] * mat_B[674] +
//             mat_A[918] * mat_B[706] +
//             mat_A[919] * mat_B[738] +
//             mat_A[920] * mat_B[770] +
//             mat_A[921] * mat_B[802] +
//             mat_A[922] * mat_B[834] +
//             mat_A[923] * mat_B[866] +
//             mat_A[924] * mat_B[898] +
//             mat_A[925] * mat_B[930] +
//             mat_A[926] * mat_B[962] +
//             mat_A[927] * mat_B[994];
//  mat_C[899] <= 
//             mat_A[896] * mat_B[3] +
//             mat_A[897] * mat_B[35] +
//             mat_A[898] * mat_B[67] +
//             mat_A[899] * mat_B[99] +
//             mat_A[900] * mat_B[131] +
//             mat_A[901] * mat_B[163] +
//             mat_A[902] * mat_B[195] +
//             mat_A[903] * mat_B[227] +
//             mat_A[904] * mat_B[259] +
//             mat_A[905] * mat_B[291] +
//             mat_A[906] * mat_B[323] +
//             mat_A[907] * mat_B[355] +
//             mat_A[908] * mat_B[387] +
//             mat_A[909] * mat_B[419] +
//             mat_A[910] * mat_B[451] +
//             mat_A[911] * mat_B[483] +
//             mat_A[912] * mat_B[515] +
//             mat_A[913] * mat_B[547] +
//             mat_A[914] * mat_B[579] +
//             mat_A[915] * mat_B[611] +
//             mat_A[916] * mat_B[643] +
//             mat_A[917] * mat_B[675] +
//             mat_A[918] * mat_B[707] +
//             mat_A[919] * mat_B[739] +
//             mat_A[920] * mat_B[771] +
//             mat_A[921] * mat_B[803] +
//             mat_A[922] * mat_B[835] +
//             mat_A[923] * mat_B[867] +
//             mat_A[924] * mat_B[899] +
//             mat_A[925] * mat_B[931] +
//             mat_A[926] * mat_B[963] +
//             mat_A[927] * mat_B[995];
//  mat_C[900] <= 
//             mat_A[896] * mat_B[4] +
//             mat_A[897] * mat_B[36] +
//             mat_A[898] * mat_B[68] +
//             mat_A[899] * mat_B[100] +
//             mat_A[900] * mat_B[132] +
//             mat_A[901] * mat_B[164] +
//             mat_A[902] * mat_B[196] +
//             mat_A[903] * mat_B[228] +
//             mat_A[904] * mat_B[260] +
//             mat_A[905] * mat_B[292] +
//             mat_A[906] * mat_B[324] +
//             mat_A[907] * mat_B[356] +
//             mat_A[908] * mat_B[388] +
//             mat_A[909] * mat_B[420] +
//             mat_A[910] * mat_B[452] +
//             mat_A[911] * mat_B[484] +
//             mat_A[912] * mat_B[516] +
//             mat_A[913] * mat_B[548] +
//             mat_A[914] * mat_B[580] +
//             mat_A[915] * mat_B[612] +
//             mat_A[916] * mat_B[644] +
//             mat_A[917] * mat_B[676] +
//             mat_A[918] * mat_B[708] +
//             mat_A[919] * mat_B[740] +
//             mat_A[920] * mat_B[772] +
//             mat_A[921] * mat_B[804] +
//             mat_A[922] * mat_B[836] +
//             mat_A[923] * mat_B[868] +
//             mat_A[924] * mat_B[900] +
//             mat_A[925] * mat_B[932] +
//             mat_A[926] * mat_B[964] +
//             mat_A[927] * mat_B[996];
//  mat_C[901] <= 
//             mat_A[896] * mat_B[5] +
//             mat_A[897] * mat_B[37] +
//             mat_A[898] * mat_B[69] +
//             mat_A[899] * mat_B[101] +
//             mat_A[900] * mat_B[133] +
//             mat_A[901] * mat_B[165] +
//             mat_A[902] * mat_B[197] +
//             mat_A[903] * mat_B[229] +
//             mat_A[904] * mat_B[261] +
//             mat_A[905] * mat_B[293] +
//             mat_A[906] * mat_B[325] +
//             mat_A[907] * mat_B[357] +
//             mat_A[908] * mat_B[389] +
//             mat_A[909] * mat_B[421] +
//             mat_A[910] * mat_B[453] +
//             mat_A[911] * mat_B[485] +
//             mat_A[912] * mat_B[517] +
//             mat_A[913] * mat_B[549] +
//             mat_A[914] * mat_B[581] +
//             mat_A[915] * mat_B[613] +
//             mat_A[916] * mat_B[645] +
//             mat_A[917] * mat_B[677] +
//             mat_A[918] * mat_B[709] +
//             mat_A[919] * mat_B[741] +
//             mat_A[920] * mat_B[773] +
//             mat_A[921] * mat_B[805] +
//             mat_A[922] * mat_B[837] +
//             mat_A[923] * mat_B[869] +
//             mat_A[924] * mat_B[901] +
//             mat_A[925] * mat_B[933] +
//             mat_A[926] * mat_B[965] +
//             mat_A[927] * mat_B[997];
//  mat_C[902] <= 
//             mat_A[896] * mat_B[6] +
//             mat_A[897] * mat_B[38] +
//             mat_A[898] * mat_B[70] +
//             mat_A[899] * mat_B[102] +
//             mat_A[900] * mat_B[134] +
//             mat_A[901] * mat_B[166] +
//             mat_A[902] * mat_B[198] +
//             mat_A[903] * mat_B[230] +
//             mat_A[904] * mat_B[262] +
//             mat_A[905] * mat_B[294] +
//             mat_A[906] * mat_B[326] +
//             mat_A[907] * mat_B[358] +
//             mat_A[908] * mat_B[390] +
//             mat_A[909] * mat_B[422] +
//             mat_A[910] * mat_B[454] +
//             mat_A[911] * mat_B[486] +
//             mat_A[912] * mat_B[518] +
//             mat_A[913] * mat_B[550] +
//             mat_A[914] * mat_B[582] +
//             mat_A[915] * mat_B[614] +
//             mat_A[916] * mat_B[646] +
//             mat_A[917] * mat_B[678] +
//             mat_A[918] * mat_B[710] +
//             mat_A[919] * mat_B[742] +
//             mat_A[920] * mat_B[774] +
//             mat_A[921] * mat_B[806] +
//             mat_A[922] * mat_B[838] +
//             mat_A[923] * mat_B[870] +
//             mat_A[924] * mat_B[902] +
//             mat_A[925] * mat_B[934] +
//             mat_A[926] * mat_B[966] +
//             mat_A[927] * mat_B[998];
//  mat_C[903] <= 
//             mat_A[896] * mat_B[7] +
//             mat_A[897] * mat_B[39] +
//             mat_A[898] * mat_B[71] +
//             mat_A[899] * mat_B[103] +
//             mat_A[900] * mat_B[135] +
//             mat_A[901] * mat_B[167] +
//             mat_A[902] * mat_B[199] +
//             mat_A[903] * mat_B[231] +
//             mat_A[904] * mat_B[263] +
//             mat_A[905] * mat_B[295] +
//             mat_A[906] * mat_B[327] +
//             mat_A[907] * mat_B[359] +
//             mat_A[908] * mat_B[391] +
//             mat_A[909] * mat_B[423] +
//             mat_A[910] * mat_B[455] +
//             mat_A[911] * mat_B[487] +
//             mat_A[912] * mat_B[519] +
//             mat_A[913] * mat_B[551] +
//             mat_A[914] * mat_B[583] +
//             mat_A[915] * mat_B[615] +
//             mat_A[916] * mat_B[647] +
//             mat_A[917] * mat_B[679] +
//             mat_A[918] * mat_B[711] +
//             mat_A[919] * mat_B[743] +
//             mat_A[920] * mat_B[775] +
//             mat_A[921] * mat_B[807] +
//             mat_A[922] * mat_B[839] +
//             mat_A[923] * mat_B[871] +
//             mat_A[924] * mat_B[903] +
//             mat_A[925] * mat_B[935] +
//             mat_A[926] * mat_B[967] +
//             mat_A[927] * mat_B[999];
//  mat_C[904] <= 
//             mat_A[896] * mat_B[8] +
//             mat_A[897] * mat_B[40] +
//             mat_A[898] * mat_B[72] +
//             mat_A[899] * mat_B[104] +
//             mat_A[900] * mat_B[136] +
//             mat_A[901] * mat_B[168] +
//             mat_A[902] * mat_B[200] +
//             mat_A[903] * mat_B[232] +
//             mat_A[904] * mat_B[264] +
//             mat_A[905] * mat_B[296] +
//             mat_A[906] * mat_B[328] +
//             mat_A[907] * mat_B[360] +
//             mat_A[908] * mat_B[392] +
//             mat_A[909] * mat_B[424] +
//             mat_A[910] * mat_B[456] +
//             mat_A[911] * mat_B[488] +
//             mat_A[912] * mat_B[520] +
//             mat_A[913] * mat_B[552] +
//             mat_A[914] * mat_B[584] +
//             mat_A[915] * mat_B[616] +
//             mat_A[916] * mat_B[648] +
//             mat_A[917] * mat_B[680] +
//             mat_A[918] * mat_B[712] +
//             mat_A[919] * mat_B[744] +
//             mat_A[920] * mat_B[776] +
//             mat_A[921] * mat_B[808] +
//             mat_A[922] * mat_B[840] +
//             mat_A[923] * mat_B[872] +
//             mat_A[924] * mat_B[904] +
//             mat_A[925] * mat_B[936] +
//             mat_A[926] * mat_B[968] +
//             mat_A[927] * mat_B[1000];
//  mat_C[905] <= 
//             mat_A[896] * mat_B[9] +
//             mat_A[897] * mat_B[41] +
//             mat_A[898] * mat_B[73] +
//             mat_A[899] * mat_B[105] +
//             mat_A[900] * mat_B[137] +
//             mat_A[901] * mat_B[169] +
//             mat_A[902] * mat_B[201] +
//             mat_A[903] * mat_B[233] +
//             mat_A[904] * mat_B[265] +
//             mat_A[905] * mat_B[297] +
//             mat_A[906] * mat_B[329] +
//             mat_A[907] * mat_B[361] +
//             mat_A[908] * mat_B[393] +
//             mat_A[909] * mat_B[425] +
//             mat_A[910] * mat_B[457] +
//             mat_A[911] * mat_B[489] +
//             mat_A[912] * mat_B[521] +
//             mat_A[913] * mat_B[553] +
//             mat_A[914] * mat_B[585] +
//             mat_A[915] * mat_B[617] +
//             mat_A[916] * mat_B[649] +
//             mat_A[917] * mat_B[681] +
//             mat_A[918] * mat_B[713] +
//             mat_A[919] * mat_B[745] +
//             mat_A[920] * mat_B[777] +
//             mat_A[921] * mat_B[809] +
//             mat_A[922] * mat_B[841] +
//             mat_A[923] * mat_B[873] +
//             mat_A[924] * mat_B[905] +
//             mat_A[925] * mat_B[937] +
//             mat_A[926] * mat_B[969] +
//             mat_A[927] * mat_B[1001];
//  mat_C[906] <= 
//             mat_A[896] * mat_B[10] +
//             mat_A[897] * mat_B[42] +
//             mat_A[898] * mat_B[74] +
//             mat_A[899] * mat_B[106] +
//             mat_A[900] * mat_B[138] +
//             mat_A[901] * mat_B[170] +
//             mat_A[902] * mat_B[202] +
//             mat_A[903] * mat_B[234] +
//             mat_A[904] * mat_B[266] +
//             mat_A[905] * mat_B[298] +
//             mat_A[906] * mat_B[330] +
//             mat_A[907] * mat_B[362] +
//             mat_A[908] * mat_B[394] +
//             mat_A[909] * mat_B[426] +
//             mat_A[910] * mat_B[458] +
//             mat_A[911] * mat_B[490] +
//             mat_A[912] * mat_B[522] +
//             mat_A[913] * mat_B[554] +
//             mat_A[914] * mat_B[586] +
//             mat_A[915] * mat_B[618] +
//             mat_A[916] * mat_B[650] +
//             mat_A[917] * mat_B[682] +
//             mat_A[918] * mat_B[714] +
//             mat_A[919] * mat_B[746] +
//             mat_A[920] * mat_B[778] +
//             mat_A[921] * mat_B[810] +
//             mat_A[922] * mat_B[842] +
//             mat_A[923] * mat_B[874] +
//             mat_A[924] * mat_B[906] +
//             mat_A[925] * mat_B[938] +
//             mat_A[926] * mat_B[970] +
//             mat_A[927] * mat_B[1002];
//  mat_C[907] <= 
//             mat_A[896] * mat_B[11] +
//             mat_A[897] * mat_B[43] +
//             mat_A[898] * mat_B[75] +
//             mat_A[899] * mat_B[107] +
//             mat_A[900] * mat_B[139] +
//             mat_A[901] * mat_B[171] +
//             mat_A[902] * mat_B[203] +
//             mat_A[903] * mat_B[235] +
//             mat_A[904] * mat_B[267] +
//             mat_A[905] * mat_B[299] +
//             mat_A[906] * mat_B[331] +
//             mat_A[907] * mat_B[363] +
//             mat_A[908] * mat_B[395] +
//             mat_A[909] * mat_B[427] +
//             mat_A[910] * mat_B[459] +
//             mat_A[911] * mat_B[491] +
//             mat_A[912] * mat_B[523] +
//             mat_A[913] * mat_B[555] +
//             mat_A[914] * mat_B[587] +
//             mat_A[915] * mat_B[619] +
//             mat_A[916] * mat_B[651] +
//             mat_A[917] * mat_B[683] +
//             mat_A[918] * mat_B[715] +
//             mat_A[919] * mat_B[747] +
//             mat_A[920] * mat_B[779] +
//             mat_A[921] * mat_B[811] +
//             mat_A[922] * mat_B[843] +
//             mat_A[923] * mat_B[875] +
//             mat_A[924] * mat_B[907] +
//             mat_A[925] * mat_B[939] +
//             mat_A[926] * mat_B[971] +
//             mat_A[927] * mat_B[1003];
//  mat_C[908] <= 
//             mat_A[896] * mat_B[12] +
//             mat_A[897] * mat_B[44] +
//             mat_A[898] * mat_B[76] +
//             mat_A[899] * mat_B[108] +
//             mat_A[900] * mat_B[140] +
//             mat_A[901] * mat_B[172] +
//             mat_A[902] * mat_B[204] +
//             mat_A[903] * mat_B[236] +
//             mat_A[904] * mat_B[268] +
//             mat_A[905] * mat_B[300] +
//             mat_A[906] * mat_B[332] +
//             mat_A[907] * mat_B[364] +
//             mat_A[908] * mat_B[396] +
//             mat_A[909] * mat_B[428] +
//             mat_A[910] * mat_B[460] +
//             mat_A[911] * mat_B[492] +
//             mat_A[912] * mat_B[524] +
//             mat_A[913] * mat_B[556] +
//             mat_A[914] * mat_B[588] +
//             mat_A[915] * mat_B[620] +
//             mat_A[916] * mat_B[652] +
//             mat_A[917] * mat_B[684] +
//             mat_A[918] * mat_B[716] +
//             mat_A[919] * mat_B[748] +
//             mat_A[920] * mat_B[780] +
//             mat_A[921] * mat_B[812] +
//             mat_A[922] * mat_B[844] +
//             mat_A[923] * mat_B[876] +
//             mat_A[924] * mat_B[908] +
//             mat_A[925] * mat_B[940] +
//             mat_A[926] * mat_B[972] +
//             mat_A[927] * mat_B[1004];
//  mat_C[909] <= 
//             mat_A[896] * mat_B[13] +
//             mat_A[897] * mat_B[45] +
//             mat_A[898] * mat_B[77] +
//             mat_A[899] * mat_B[109] +
//             mat_A[900] * mat_B[141] +
//             mat_A[901] * mat_B[173] +
//             mat_A[902] * mat_B[205] +
//             mat_A[903] * mat_B[237] +
//             mat_A[904] * mat_B[269] +
//             mat_A[905] * mat_B[301] +
//             mat_A[906] * mat_B[333] +
//             mat_A[907] * mat_B[365] +
//             mat_A[908] * mat_B[397] +
//             mat_A[909] * mat_B[429] +
//             mat_A[910] * mat_B[461] +
//             mat_A[911] * mat_B[493] +
//             mat_A[912] * mat_B[525] +
//             mat_A[913] * mat_B[557] +
//             mat_A[914] * mat_B[589] +
//             mat_A[915] * mat_B[621] +
//             mat_A[916] * mat_B[653] +
//             mat_A[917] * mat_B[685] +
//             mat_A[918] * mat_B[717] +
//             mat_A[919] * mat_B[749] +
//             mat_A[920] * mat_B[781] +
//             mat_A[921] * mat_B[813] +
//             mat_A[922] * mat_B[845] +
//             mat_A[923] * mat_B[877] +
//             mat_A[924] * mat_B[909] +
//             mat_A[925] * mat_B[941] +
//             mat_A[926] * mat_B[973] +
//             mat_A[927] * mat_B[1005];
//  mat_C[910] <= 
//             mat_A[896] * mat_B[14] +
//             mat_A[897] * mat_B[46] +
//             mat_A[898] * mat_B[78] +
//             mat_A[899] * mat_B[110] +
//             mat_A[900] * mat_B[142] +
//             mat_A[901] * mat_B[174] +
//             mat_A[902] * mat_B[206] +
//             mat_A[903] * mat_B[238] +
//             mat_A[904] * mat_B[270] +
//             mat_A[905] * mat_B[302] +
//             mat_A[906] * mat_B[334] +
//             mat_A[907] * mat_B[366] +
//             mat_A[908] * mat_B[398] +
//             mat_A[909] * mat_B[430] +
//             mat_A[910] * mat_B[462] +
//             mat_A[911] * mat_B[494] +
//             mat_A[912] * mat_B[526] +
//             mat_A[913] * mat_B[558] +
//             mat_A[914] * mat_B[590] +
//             mat_A[915] * mat_B[622] +
//             mat_A[916] * mat_B[654] +
//             mat_A[917] * mat_B[686] +
//             mat_A[918] * mat_B[718] +
//             mat_A[919] * mat_B[750] +
//             mat_A[920] * mat_B[782] +
//             mat_A[921] * mat_B[814] +
//             mat_A[922] * mat_B[846] +
//             mat_A[923] * mat_B[878] +
//             mat_A[924] * mat_B[910] +
//             mat_A[925] * mat_B[942] +
//             mat_A[926] * mat_B[974] +
//             mat_A[927] * mat_B[1006];
//  mat_C[911] <= 
//             mat_A[896] * mat_B[15] +
//             mat_A[897] * mat_B[47] +
//             mat_A[898] * mat_B[79] +
//             mat_A[899] * mat_B[111] +
//             mat_A[900] * mat_B[143] +
//             mat_A[901] * mat_B[175] +
//             mat_A[902] * mat_B[207] +
//             mat_A[903] * mat_B[239] +
//             mat_A[904] * mat_B[271] +
//             mat_A[905] * mat_B[303] +
//             mat_A[906] * mat_B[335] +
//             mat_A[907] * mat_B[367] +
//             mat_A[908] * mat_B[399] +
//             mat_A[909] * mat_B[431] +
//             mat_A[910] * mat_B[463] +
//             mat_A[911] * mat_B[495] +
//             mat_A[912] * mat_B[527] +
//             mat_A[913] * mat_B[559] +
//             mat_A[914] * mat_B[591] +
//             mat_A[915] * mat_B[623] +
//             mat_A[916] * mat_B[655] +
//             mat_A[917] * mat_B[687] +
//             mat_A[918] * mat_B[719] +
//             mat_A[919] * mat_B[751] +
//             mat_A[920] * mat_B[783] +
//             mat_A[921] * mat_B[815] +
//             mat_A[922] * mat_B[847] +
//             mat_A[923] * mat_B[879] +
//             mat_A[924] * mat_B[911] +
//             mat_A[925] * mat_B[943] +
//             mat_A[926] * mat_B[975] +
//             mat_A[927] * mat_B[1007];
//  mat_C[912] <= 
//             mat_A[896] * mat_B[16] +
//             mat_A[897] * mat_B[48] +
//             mat_A[898] * mat_B[80] +
//             mat_A[899] * mat_B[112] +
//             mat_A[900] * mat_B[144] +
//             mat_A[901] * mat_B[176] +
//             mat_A[902] * mat_B[208] +
//             mat_A[903] * mat_B[240] +
//             mat_A[904] * mat_B[272] +
//             mat_A[905] * mat_B[304] +
//             mat_A[906] * mat_B[336] +
//             mat_A[907] * mat_B[368] +
//             mat_A[908] * mat_B[400] +
//             mat_A[909] * mat_B[432] +
//             mat_A[910] * mat_B[464] +
//             mat_A[911] * mat_B[496] +
//             mat_A[912] * mat_B[528] +
//             mat_A[913] * mat_B[560] +
//             mat_A[914] * mat_B[592] +
//             mat_A[915] * mat_B[624] +
//             mat_A[916] * mat_B[656] +
//             mat_A[917] * mat_B[688] +
//             mat_A[918] * mat_B[720] +
//             mat_A[919] * mat_B[752] +
//             mat_A[920] * mat_B[784] +
//             mat_A[921] * mat_B[816] +
//             mat_A[922] * mat_B[848] +
//             mat_A[923] * mat_B[880] +
//             mat_A[924] * mat_B[912] +
//             mat_A[925] * mat_B[944] +
//             mat_A[926] * mat_B[976] +
//             mat_A[927] * mat_B[1008];
//  mat_C[913] <= 
//             mat_A[896] * mat_B[17] +
//             mat_A[897] * mat_B[49] +
//             mat_A[898] * mat_B[81] +
//             mat_A[899] * mat_B[113] +
//             mat_A[900] * mat_B[145] +
//             mat_A[901] * mat_B[177] +
//             mat_A[902] * mat_B[209] +
//             mat_A[903] * mat_B[241] +
//             mat_A[904] * mat_B[273] +
//             mat_A[905] * mat_B[305] +
//             mat_A[906] * mat_B[337] +
//             mat_A[907] * mat_B[369] +
//             mat_A[908] * mat_B[401] +
//             mat_A[909] * mat_B[433] +
//             mat_A[910] * mat_B[465] +
//             mat_A[911] * mat_B[497] +
//             mat_A[912] * mat_B[529] +
//             mat_A[913] * mat_B[561] +
//             mat_A[914] * mat_B[593] +
//             mat_A[915] * mat_B[625] +
//             mat_A[916] * mat_B[657] +
//             mat_A[917] * mat_B[689] +
//             mat_A[918] * mat_B[721] +
//             mat_A[919] * mat_B[753] +
//             mat_A[920] * mat_B[785] +
//             mat_A[921] * mat_B[817] +
//             mat_A[922] * mat_B[849] +
//             mat_A[923] * mat_B[881] +
//             mat_A[924] * mat_B[913] +
//             mat_A[925] * mat_B[945] +
//             mat_A[926] * mat_B[977] +
//             mat_A[927] * mat_B[1009];
//  mat_C[914] <= 
//             mat_A[896] * mat_B[18] +
//             mat_A[897] * mat_B[50] +
//             mat_A[898] * mat_B[82] +
//             mat_A[899] * mat_B[114] +
//             mat_A[900] * mat_B[146] +
//             mat_A[901] * mat_B[178] +
//             mat_A[902] * mat_B[210] +
//             mat_A[903] * mat_B[242] +
//             mat_A[904] * mat_B[274] +
//             mat_A[905] * mat_B[306] +
//             mat_A[906] * mat_B[338] +
//             mat_A[907] * mat_B[370] +
//             mat_A[908] * mat_B[402] +
//             mat_A[909] * mat_B[434] +
//             mat_A[910] * mat_B[466] +
//             mat_A[911] * mat_B[498] +
//             mat_A[912] * mat_B[530] +
//             mat_A[913] * mat_B[562] +
//             mat_A[914] * mat_B[594] +
//             mat_A[915] * mat_B[626] +
//             mat_A[916] * mat_B[658] +
//             mat_A[917] * mat_B[690] +
//             mat_A[918] * mat_B[722] +
//             mat_A[919] * mat_B[754] +
//             mat_A[920] * mat_B[786] +
//             mat_A[921] * mat_B[818] +
//             mat_A[922] * mat_B[850] +
//             mat_A[923] * mat_B[882] +
//             mat_A[924] * mat_B[914] +
//             mat_A[925] * mat_B[946] +
//             mat_A[926] * mat_B[978] +
//             mat_A[927] * mat_B[1010];
//  mat_C[915] <= 
//             mat_A[896] * mat_B[19] +
//             mat_A[897] * mat_B[51] +
//             mat_A[898] * mat_B[83] +
//             mat_A[899] * mat_B[115] +
//             mat_A[900] * mat_B[147] +
//             mat_A[901] * mat_B[179] +
//             mat_A[902] * mat_B[211] +
//             mat_A[903] * mat_B[243] +
//             mat_A[904] * mat_B[275] +
//             mat_A[905] * mat_B[307] +
//             mat_A[906] * mat_B[339] +
//             mat_A[907] * mat_B[371] +
//             mat_A[908] * mat_B[403] +
//             mat_A[909] * mat_B[435] +
//             mat_A[910] * mat_B[467] +
//             mat_A[911] * mat_B[499] +
//             mat_A[912] * mat_B[531] +
//             mat_A[913] * mat_B[563] +
//             mat_A[914] * mat_B[595] +
//             mat_A[915] * mat_B[627] +
//             mat_A[916] * mat_B[659] +
//             mat_A[917] * mat_B[691] +
//             mat_A[918] * mat_B[723] +
//             mat_A[919] * mat_B[755] +
//             mat_A[920] * mat_B[787] +
//             mat_A[921] * mat_B[819] +
//             mat_A[922] * mat_B[851] +
//             mat_A[923] * mat_B[883] +
//             mat_A[924] * mat_B[915] +
//             mat_A[925] * mat_B[947] +
//             mat_A[926] * mat_B[979] +
//             mat_A[927] * mat_B[1011];
//  mat_C[916] <= 
//             mat_A[896] * mat_B[20] +
//             mat_A[897] * mat_B[52] +
//             mat_A[898] * mat_B[84] +
//             mat_A[899] * mat_B[116] +
//             mat_A[900] * mat_B[148] +
//             mat_A[901] * mat_B[180] +
//             mat_A[902] * mat_B[212] +
//             mat_A[903] * mat_B[244] +
//             mat_A[904] * mat_B[276] +
//             mat_A[905] * mat_B[308] +
//             mat_A[906] * mat_B[340] +
//             mat_A[907] * mat_B[372] +
//             mat_A[908] * mat_B[404] +
//             mat_A[909] * mat_B[436] +
//             mat_A[910] * mat_B[468] +
//             mat_A[911] * mat_B[500] +
//             mat_A[912] * mat_B[532] +
//             mat_A[913] * mat_B[564] +
//             mat_A[914] * mat_B[596] +
//             mat_A[915] * mat_B[628] +
//             mat_A[916] * mat_B[660] +
//             mat_A[917] * mat_B[692] +
//             mat_A[918] * mat_B[724] +
//             mat_A[919] * mat_B[756] +
//             mat_A[920] * mat_B[788] +
//             mat_A[921] * mat_B[820] +
//             mat_A[922] * mat_B[852] +
//             mat_A[923] * mat_B[884] +
//             mat_A[924] * mat_B[916] +
//             mat_A[925] * mat_B[948] +
//             mat_A[926] * mat_B[980] +
//             mat_A[927] * mat_B[1012];
//  mat_C[917] <= 
//             mat_A[896] * mat_B[21] +
//             mat_A[897] * mat_B[53] +
//             mat_A[898] * mat_B[85] +
//             mat_A[899] * mat_B[117] +
//             mat_A[900] * mat_B[149] +
//             mat_A[901] * mat_B[181] +
//             mat_A[902] * mat_B[213] +
//             mat_A[903] * mat_B[245] +
//             mat_A[904] * mat_B[277] +
//             mat_A[905] * mat_B[309] +
//             mat_A[906] * mat_B[341] +
//             mat_A[907] * mat_B[373] +
//             mat_A[908] * mat_B[405] +
//             mat_A[909] * mat_B[437] +
//             mat_A[910] * mat_B[469] +
//             mat_A[911] * mat_B[501] +
//             mat_A[912] * mat_B[533] +
//             mat_A[913] * mat_B[565] +
//             mat_A[914] * mat_B[597] +
//             mat_A[915] * mat_B[629] +
//             mat_A[916] * mat_B[661] +
//             mat_A[917] * mat_B[693] +
//             mat_A[918] * mat_B[725] +
//             mat_A[919] * mat_B[757] +
//             mat_A[920] * mat_B[789] +
//             mat_A[921] * mat_B[821] +
//             mat_A[922] * mat_B[853] +
//             mat_A[923] * mat_B[885] +
//             mat_A[924] * mat_B[917] +
//             mat_A[925] * mat_B[949] +
//             mat_A[926] * mat_B[981] +
//             mat_A[927] * mat_B[1013];
//  mat_C[918] <= 
//             mat_A[896] * mat_B[22] +
//             mat_A[897] * mat_B[54] +
//             mat_A[898] * mat_B[86] +
//             mat_A[899] * mat_B[118] +
//             mat_A[900] * mat_B[150] +
//             mat_A[901] * mat_B[182] +
//             mat_A[902] * mat_B[214] +
//             mat_A[903] * mat_B[246] +
//             mat_A[904] * mat_B[278] +
//             mat_A[905] * mat_B[310] +
//             mat_A[906] * mat_B[342] +
//             mat_A[907] * mat_B[374] +
//             mat_A[908] * mat_B[406] +
//             mat_A[909] * mat_B[438] +
//             mat_A[910] * mat_B[470] +
//             mat_A[911] * mat_B[502] +
//             mat_A[912] * mat_B[534] +
//             mat_A[913] * mat_B[566] +
//             mat_A[914] * mat_B[598] +
//             mat_A[915] * mat_B[630] +
//             mat_A[916] * mat_B[662] +
//             mat_A[917] * mat_B[694] +
//             mat_A[918] * mat_B[726] +
//             mat_A[919] * mat_B[758] +
//             mat_A[920] * mat_B[790] +
//             mat_A[921] * mat_B[822] +
//             mat_A[922] * mat_B[854] +
//             mat_A[923] * mat_B[886] +
//             mat_A[924] * mat_B[918] +
//             mat_A[925] * mat_B[950] +
//             mat_A[926] * mat_B[982] +
//             mat_A[927] * mat_B[1014];
//  mat_C[919] <= 
//             mat_A[896] * mat_B[23] +
//             mat_A[897] * mat_B[55] +
//             mat_A[898] * mat_B[87] +
//             mat_A[899] * mat_B[119] +
//             mat_A[900] * mat_B[151] +
//             mat_A[901] * mat_B[183] +
//             mat_A[902] * mat_B[215] +
//             mat_A[903] * mat_B[247] +
//             mat_A[904] * mat_B[279] +
//             mat_A[905] * mat_B[311] +
//             mat_A[906] * mat_B[343] +
//             mat_A[907] * mat_B[375] +
//             mat_A[908] * mat_B[407] +
//             mat_A[909] * mat_B[439] +
//             mat_A[910] * mat_B[471] +
//             mat_A[911] * mat_B[503] +
//             mat_A[912] * mat_B[535] +
//             mat_A[913] * mat_B[567] +
//             mat_A[914] * mat_B[599] +
//             mat_A[915] * mat_B[631] +
//             mat_A[916] * mat_B[663] +
//             mat_A[917] * mat_B[695] +
//             mat_A[918] * mat_B[727] +
//             mat_A[919] * mat_B[759] +
//             mat_A[920] * mat_B[791] +
//             mat_A[921] * mat_B[823] +
//             mat_A[922] * mat_B[855] +
//             mat_A[923] * mat_B[887] +
//             mat_A[924] * mat_B[919] +
//             mat_A[925] * mat_B[951] +
//             mat_A[926] * mat_B[983] +
//             mat_A[927] * mat_B[1015];
//  mat_C[920] <= 
//             mat_A[896] * mat_B[24] +
//             mat_A[897] * mat_B[56] +
//             mat_A[898] * mat_B[88] +
//             mat_A[899] * mat_B[120] +
//             mat_A[900] * mat_B[152] +
//             mat_A[901] * mat_B[184] +
//             mat_A[902] * mat_B[216] +
//             mat_A[903] * mat_B[248] +
//             mat_A[904] * mat_B[280] +
//             mat_A[905] * mat_B[312] +
//             mat_A[906] * mat_B[344] +
//             mat_A[907] * mat_B[376] +
//             mat_A[908] * mat_B[408] +
//             mat_A[909] * mat_B[440] +
//             mat_A[910] * mat_B[472] +
//             mat_A[911] * mat_B[504] +
//             mat_A[912] * mat_B[536] +
//             mat_A[913] * mat_B[568] +
//             mat_A[914] * mat_B[600] +
//             mat_A[915] * mat_B[632] +
//             mat_A[916] * mat_B[664] +
//             mat_A[917] * mat_B[696] +
//             mat_A[918] * mat_B[728] +
//             mat_A[919] * mat_B[760] +
//             mat_A[920] * mat_B[792] +
//             mat_A[921] * mat_B[824] +
//             mat_A[922] * mat_B[856] +
//             mat_A[923] * mat_B[888] +
//             mat_A[924] * mat_B[920] +
//             mat_A[925] * mat_B[952] +
//             mat_A[926] * mat_B[984] +
//             mat_A[927] * mat_B[1016];
//  mat_C[921] <= 
//             mat_A[896] * mat_B[25] +
//             mat_A[897] * mat_B[57] +
//             mat_A[898] * mat_B[89] +
//             mat_A[899] * mat_B[121] +
//             mat_A[900] * mat_B[153] +
//             mat_A[901] * mat_B[185] +
//             mat_A[902] * mat_B[217] +
//             mat_A[903] * mat_B[249] +
//             mat_A[904] * mat_B[281] +
//             mat_A[905] * mat_B[313] +
//             mat_A[906] * mat_B[345] +
//             mat_A[907] * mat_B[377] +
//             mat_A[908] * mat_B[409] +
//             mat_A[909] * mat_B[441] +
//             mat_A[910] * mat_B[473] +
//             mat_A[911] * mat_B[505] +
//             mat_A[912] * mat_B[537] +
//             mat_A[913] * mat_B[569] +
//             mat_A[914] * mat_B[601] +
//             mat_A[915] * mat_B[633] +
//             mat_A[916] * mat_B[665] +
//             mat_A[917] * mat_B[697] +
//             mat_A[918] * mat_B[729] +
//             mat_A[919] * mat_B[761] +
//             mat_A[920] * mat_B[793] +
//             mat_A[921] * mat_B[825] +
//             mat_A[922] * mat_B[857] +
//             mat_A[923] * mat_B[889] +
//             mat_A[924] * mat_B[921] +
//             mat_A[925] * mat_B[953] +
//             mat_A[926] * mat_B[985] +
//             mat_A[927] * mat_B[1017];
//  mat_C[922] <= 
//             mat_A[896] * mat_B[26] +
//             mat_A[897] * mat_B[58] +
//             mat_A[898] * mat_B[90] +
//             mat_A[899] * mat_B[122] +
//             mat_A[900] * mat_B[154] +
//             mat_A[901] * mat_B[186] +
//             mat_A[902] * mat_B[218] +
//             mat_A[903] * mat_B[250] +
//             mat_A[904] * mat_B[282] +
//             mat_A[905] * mat_B[314] +
//             mat_A[906] * mat_B[346] +
//             mat_A[907] * mat_B[378] +
//             mat_A[908] * mat_B[410] +
//             mat_A[909] * mat_B[442] +
//             mat_A[910] * mat_B[474] +
//             mat_A[911] * mat_B[506] +
//             mat_A[912] * mat_B[538] +
//             mat_A[913] * mat_B[570] +
//             mat_A[914] * mat_B[602] +
//             mat_A[915] * mat_B[634] +
//             mat_A[916] * mat_B[666] +
//             mat_A[917] * mat_B[698] +
//             mat_A[918] * mat_B[730] +
//             mat_A[919] * mat_B[762] +
//             mat_A[920] * mat_B[794] +
//             mat_A[921] * mat_B[826] +
//             mat_A[922] * mat_B[858] +
//             mat_A[923] * mat_B[890] +
//             mat_A[924] * mat_B[922] +
//             mat_A[925] * mat_B[954] +
//             mat_A[926] * mat_B[986] +
//             mat_A[927] * mat_B[1018];
//  mat_C[923] <= 
//             mat_A[896] * mat_B[27] +
//             mat_A[897] * mat_B[59] +
//             mat_A[898] * mat_B[91] +
//             mat_A[899] * mat_B[123] +
//             mat_A[900] * mat_B[155] +
//             mat_A[901] * mat_B[187] +
//             mat_A[902] * mat_B[219] +
//             mat_A[903] * mat_B[251] +
//             mat_A[904] * mat_B[283] +
//             mat_A[905] * mat_B[315] +
//             mat_A[906] * mat_B[347] +
//             mat_A[907] * mat_B[379] +
//             mat_A[908] * mat_B[411] +
//             mat_A[909] * mat_B[443] +
//             mat_A[910] * mat_B[475] +
//             mat_A[911] * mat_B[507] +
//             mat_A[912] * mat_B[539] +
//             mat_A[913] * mat_B[571] +
//             mat_A[914] * mat_B[603] +
//             mat_A[915] * mat_B[635] +
//             mat_A[916] * mat_B[667] +
//             mat_A[917] * mat_B[699] +
//             mat_A[918] * mat_B[731] +
//             mat_A[919] * mat_B[763] +
//             mat_A[920] * mat_B[795] +
//             mat_A[921] * mat_B[827] +
//             mat_A[922] * mat_B[859] +
//             mat_A[923] * mat_B[891] +
//             mat_A[924] * mat_B[923] +
//             mat_A[925] * mat_B[955] +
//             mat_A[926] * mat_B[987] +
//             mat_A[927] * mat_B[1019];
//  mat_C[924] <= 
//             mat_A[896] * mat_B[28] +
//             mat_A[897] * mat_B[60] +
//             mat_A[898] * mat_B[92] +
//             mat_A[899] * mat_B[124] +
//             mat_A[900] * mat_B[156] +
//             mat_A[901] * mat_B[188] +
//             mat_A[902] * mat_B[220] +
//             mat_A[903] * mat_B[252] +
//             mat_A[904] * mat_B[284] +
//             mat_A[905] * mat_B[316] +
//             mat_A[906] * mat_B[348] +
//             mat_A[907] * mat_B[380] +
//             mat_A[908] * mat_B[412] +
//             mat_A[909] * mat_B[444] +
//             mat_A[910] * mat_B[476] +
//             mat_A[911] * mat_B[508] +
//             mat_A[912] * mat_B[540] +
//             mat_A[913] * mat_B[572] +
//             mat_A[914] * mat_B[604] +
//             mat_A[915] * mat_B[636] +
//             mat_A[916] * mat_B[668] +
//             mat_A[917] * mat_B[700] +
//             mat_A[918] * mat_B[732] +
//             mat_A[919] * mat_B[764] +
//             mat_A[920] * mat_B[796] +
//             mat_A[921] * mat_B[828] +
//             mat_A[922] * mat_B[860] +
//             mat_A[923] * mat_B[892] +
//             mat_A[924] * mat_B[924] +
//             mat_A[925] * mat_B[956] +
//             mat_A[926] * mat_B[988] +
//             mat_A[927] * mat_B[1020];
//  mat_C[925] <= 
//             mat_A[896] * mat_B[29] +
//             mat_A[897] * mat_B[61] +
//             mat_A[898] * mat_B[93] +
//             mat_A[899] * mat_B[125] +
//             mat_A[900] * mat_B[157] +
//             mat_A[901] * mat_B[189] +
//             mat_A[902] * mat_B[221] +
//             mat_A[903] * mat_B[253] +
//             mat_A[904] * mat_B[285] +
//             mat_A[905] * mat_B[317] +
//             mat_A[906] * mat_B[349] +
//             mat_A[907] * mat_B[381] +
//             mat_A[908] * mat_B[413] +
//             mat_A[909] * mat_B[445] +
//             mat_A[910] * mat_B[477] +
//             mat_A[911] * mat_B[509] +
//             mat_A[912] * mat_B[541] +
//             mat_A[913] * mat_B[573] +
//             mat_A[914] * mat_B[605] +
//             mat_A[915] * mat_B[637] +
//             mat_A[916] * mat_B[669] +
//             mat_A[917] * mat_B[701] +
//             mat_A[918] * mat_B[733] +
//             mat_A[919] * mat_B[765] +
//             mat_A[920] * mat_B[797] +
//             mat_A[921] * mat_B[829] +
//             mat_A[922] * mat_B[861] +
//             mat_A[923] * mat_B[893] +
//             mat_A[924] * mat_B[925] +
//             mat_A[925] * mat_B[957] +
//             mat_A[926] * mat_B[989] +
//             mat_A[927] * mat_B[1021];
//  mat_C[926] <= 
//             mat_A[896] * mat_B[30] +
//             mat_A[897] * mat_B[62] +
//             mat_A[898] * mat_B[94] +
//             mat_A[899] * mat_B[126] +
//             mat_A[900] * mat_B[158] +
//             mat_A[901] * mat_B[190] +
//             mat_A[902] * mat_B[222] +
//             mat_A[903] * mat_B[254] +
//             mat_A[904] * mat_B[286] +
//             mat_A[905] * mat_B[318] +
//             mat_A[906] * mat_B[350] +
//             mat_A[907] * mat_B[382] +
//             mat_A[908] * mat_B[414] +
//             mat_A[909] * mat_B[446] +
//             mat_A[910] * mat_B[478] +
//             mat_A[911] * mat_B[510] +
//             mat_A[912] * mat_B[542] +
//             mat_A[913] * mat_B[574] +
//             mat_A[914] * mat_B[606] +
//             mat_A[915] * mat_B[638] +
//             mat_A[916] * mat_B[670] +
//             mat_A[917] * mat_B[702] +
//             mat_A[918] * mat_B[734] +
//             mat_A[919] * mat_B[766] +
//             mat_A[920] * mat_B[798] +
//             mat_A[921] * mat_B[830] +
//             mat_A[922] * mat_B[862] +
//             mat_A[923] * mat_B[894] +
//             mat_A[924] * mat_B[926] +
//             mat_A[925] * mat_B[958] +
//             mat_A[926] * mat_B[990] +
//             mat_A[927] * mat_B[1022];
//  mat_C[927] <= 
//             mat_A[896] * mat_B[31] +
//             mat_A[897] * mat_B[63] +
//             mat_A[898] * mat_B[95] +
//             mat_A[899] * mat_B[127] +
//             mat_A[900] * mat_B[159] +
//             mat_A[901] * mat_B[191] +
//             mat_A[902] * mat_B[223] +
//             mat_A[903] * mat_B[255] +
//             mat_A[904] * mat_B[287] +
//             mat_A[905] * mat_B[319] +
//             mat_A[906] * mat_B[351] +
//             mat_A[907] * mat_B[383] +
//             mat_A[908] * mat_B[415] +
//             mat_A[909] * mat_B[447] +
//             mat_A[910] * mat_B[479] +
//             mat_A[911] * mat_B[511] +
//             mat_A[912] * mat_B[543] +
//             mat_A[913] * mat_B[575] +
//             mat_A[914] * mat_B[607] +
//             mat_A[915] * mat_B[639] +
//             mat_A[916] * mat_B[671] +
//             mat_A[917] * mat_B[703] +
//             mat_A[918] * mat_B[735] +
//             mat_A[919] * mat_B[767] +
//             mat_A[920] * mat_B[799] +
//             mat_A[921] * mat_B[831] +
//             mat_A[922] * mat_B[863] +
//             mat_A[923] * mat_B[895] +
//             mat_A[924] * mat_B[927] +
//             mat_A[925] * mat_B[959] +
//             mat_A[926] * mat_B[991] +
//             mat_A[927] * mat_B[1023];
//  mat_C[928] <= 
//             mat_A[928] * mat_B[0] +
//             mat_A[929] * mat_B[32] +
//             mat_A[930] * mat_B[64] +
//             mat_A[931] * mat_B[96] +
//             mat_A[932] * mat_B[128] +
//             mat_A[933] * mat_B[160] +
//             mat_A[934] * mat_B[192] +
//             mat_A[935] * mat_B[224] +
//             mat_A[936] * mat_B[256] +
//             mat_A[937] * mat_B[288] +
//             mat_A[938] * mat_B[320] +
//             mat_A[939] * mat_B[352] +
//             mat_A[940] * mat_B[384] +
//             mat_A[941] * mat_B[416] +
//             mat_A[942] * mat_B[448] +
//             mat_A[943] * mat_B[480] +
//             mat_A[944] * mat_B[512] +
//             mat_A[945] * mat_B[544] +
//             mat_A[946] * mat_B[576] +
//             mat_A[947] * mat_B[608] +
//             mat_A[948] * mat_B[640] +
//             mat_A[949] * mat_B[672] +
//             mat_A[950] * mat_B[704] +
//             mat_A[951] * mat_B[736] +
//             mat_A[952] * mat_B[768] +
//             mat_A[953] * mat_B[800] +
//             mat_A[954] * mat_B[832] +
//             mat_A[955] * mat_B[864] +
//             mat_A[956] * mat_B[896] +
//             mat_A[957] * mat_B[928] +
//             mat_A[958] * mat_B[960] +
//             mat_A[959] * mat_B[992];
//  mat_C[929] <= 
//             mat_A[928] * mat_B[1] +
//             mat_A[929] * mat_B[33] +
//             mat_A[930] * mat_B[65] +
//             mat_A[931] * mat_B[97] +
//             mat_A[932] * mat_B[129] +
//             mat_A[933] * mat_B[161] +
//             mat_A[934] * mat_B[193] +
//             mat_A[935] * mat_B[225] +
//             mat_A[936] * mat_B[257] +
//             mat_A[937] * mat_B[289] +
//             mat_A[938] * mat_B[321] +
//             mat_A[939] * mat_B[353] +
//             mat_A[940] * mat_B[385] +
//             mat_A[941] * mat_B[417] +
//             mat_A[942] * mat_B[449] +
//             mat_A[943] * mat_B[481] +
//             mat_A[944] * mat_B[513] +
//             mat_A[945] * mat_B[545] +
//             mat_A[946] * mat_B[577] +
//             mat_A[947] * mat_B[609] +
//             mat_A[948] * mat_B[641] +
//             mat_A[949] * mat_B[673] +
//             mat_A[950] * mat_B[705] +
//             mat_A[951] * mat_B[737] +
//             mat_A[952] * mat_B[769] +
//             mat_A[953] * mat_B[801] +
//             mat_A[954] * mat_B[833] +
//             mat_A[955] * mat_B[865] +
//             mat_A[956] * mat_B[897] +
//             mat_A[957] * mat_B[929] +
//             mat_A[958] * mat_B[961] +
//             mat_A[959] * mat_B[993];
//  mat_C[930] <= 
//             mat_A[928] * mat_B[2] +
//             mat_A[929] * mat_B[34] +
//             mat_A[930] * mat_B[66] +
//             mat_A[931] * mat_B[98] +
//             mat_A[932] * mat_B[130] +
//             mat_A[933] * mat_B[162] +
//             mat_A[934] * mat_B[194] +
//             mat_A[935] * mat_B[226] +
//             mat_A[936] * mat_B[258] +
//             mat_A[937] * mat_B[290] +
//             mat_A[938] * mat_B[322] +
//             mat_A[939] * mat_B[354] +
//             mat_A[940] * mat_B[386] +
//             mat_A[941] * mat_B[418] +
//             mat_A[942] * mat_B[450] +
//             mat_A[943] * mat_B[482] +
//             mat_A[944] * mat_B[514] +
//             mat_A[945] * mat_B[546] +
//             mat_A[946] * mat_B[578] +
//             mat_A[947] * mat_B[610] +
//             mat_A[948] * mat_B[642] +
//             mat_A[949] * mat_B[674] +
//             mat_A[950] * mat_B[706] +
//             mat_A[951] * mat_B[738] +
//             mat_A[952] * mat_B[770] +
//             mat_A[953] * mat_B[802] +
//             mat_A[954] * mat_B[834] +
//             mat_A[955] * mat_B[866] +
//             mat_A[956] * mat_B[898] +
//             mat_A[957] * mat_B[930] +
//             mat_A[958] * mat_B[962] +
//             mat_A[959] * mat_B[994];
//  mat_C[931] <= 
//             mat_A[928] * mat_B[3] +
//             mat_A[929] * mat_B[35] +
//             mat_A[930] * mat_B[67] +
//             mat_A[931] * mat_B[99] +
//             mat_A[932] * mat_B[131] +
//             mat_A[933] * mat_B[163] +
//             mat_A[934] * mat_B[195] +
//             mat_A[935] * mat_B[227] +
//             mat_A[936] * mat_B[259] +
//             mat_A[937] * mat_B[291] +
//             mat_A[938] * mat_B[323] +
//             mat_A[939] * mat_B[355] +
//             mat_A[940] * mat_B[387] +
//             mat_A[941] * mat_B[419] +
//             mat_A[942] * mat_B[451] +
//             mat_A[943] * mat_B[483] +
//             mat_A[944] * mat_B[515] +
//             mat_A[945] * mat_B[547] +
//             mat_A[946] * mat_B[579] +
//             mat_A[947] * mat_B[611] +
//             mat_A[948] * mat_B[643] +
//             mat_A[949] * mat_B[675] +
//             mat_A[950] * mat_B[707] +
//             mat_A[951] * mat_B[739] +
//             mat_A[952] * mat_B[771] +
//             mat_A[953] * mat_B[803] +
//             mat_A[954] * mat_B[835] +
//             mat_A[955] * mat_B[867] +
//             mat_A[956] * mat_B[899] +
//             mat_A[957] * mat_B[931] +
//             mat_A[958] * mat_B[963] +
//             mat_A[959] * mat_B[995];
//  mat_C[932] <= 
//             mat_A[928] * mat_B[4] +
//             mat_A[929] * mat_B[36] +
//             mat_A[930] * mat_B[68] +
//             mat_A[931] * mat_B[100] +
//             mat_A[932] * mat_B[132] +
//             mat_A[933] * mat_B[164] +
//             mat_A[934] * mat_B[196] +
//             mat_A[935] * mat_B[228] +
//             mat_A[936] * mat_B[260] +
//             mat_A[937] * mat_B[292] +
//             mat_A[938] * mat_B[324] +
//             mat_A[939] * mat_B[356] +
//             mat_A[940] * mat_B[388] +
//             mat_A[941] * mat_B[420] +
//             mat_A[942] * mat_B[452] +
//             mat_A[943] * mat_B[484] +
//             mat_A[944] * mat_B[516] +
//             mat_A[945] * mat_B[548] +
//             mat_A[946] * mat_B[580] +
//             mat_A[947] * mat_B[612] +
//             mat_A[948] * mat_B[644] +
//             mat_A[949] * mat_B[676] +
//             mat_A[950] * mat_B[708] +
//             mat_A[951] * mat_B[740] +
//             mat_A[952] * mat_B[772] +
//             mat_A[953] * mat_B[804] +
//             mat_A[954] * mat_B[836] +
//             mat_A[955] * mat_B[868] +
//             mat_A[956] * mat_B[900] +
//             mat_A[957] * mat_B[932] +
//             mat_A[958] * mat_B[964] +
//             mat_A[959] * mat_B[996];
//  mat_C[933] <= 
//             mat_A[928] * mat_B[5] +
//             mat_A[929] * mat_B[37] +
//             mat_A[930] * mat_B[69] +
//             mat_A[931] * mat_B[101] +
//             mat_A[932] * mat_B[133] +
//             mat_A[933] * mat_B[165] +
//             mat_A[934] * mat_B[197] +
//             mat_A[935] * mat_B[229] +
//             mat_A[936] * mat_B[261] +
//             mat_A[937] * mat_B[293] +
//             mat_A[938] * mat_B[325] +
//             mat_A[939] * mat_B[357] +
//             mat_A[940] * mat_B[389] +
//             mat_A[941] * mat_B[421] +
//             mat_A[942] * mat_B[453] +
//             mat_A[943] * mat_B[485] +
//             mat_A[944] * mat_B[517] +
//             mat_A[945] * mat_B[549] +
//             mat_A[946] * mat_B[581] +
//             mat_A[947] * mat_B[613] +
//             mat_A[948] * mat_B[645] +
//             mat_A[949] * mat_B[677] +
//             mat_A[950] * mat_B[709] +
//             mat_A[951] * mat_B[741] +
//             mat_A[952] * mat_B[773] +
//             mat_A[953] * mat_B[805] +
//             mat_A[954] * mat_B[837] +
//             mat_A[955] * mat_B[869] +
//             mat_A[956] * mat_B[901] +
//             mat_A[957] * mat_B[933] +
//             mat_A[958] * mat_B[965] +
//             mat_A[959] * mat_B[997];
//  mat_C[934] <= 
//             mat_A[928] * mat_B[6] +
//             mat_A[929] * mat_B[38] +
//             mat_A[930] * mat_B[70] +
//             mat_A[931] * mat_B[102] +
//             mat_A[932] * mat_B[134] +
//             mat_A[933] * mat_B[166] +
//             mat_A[934] * mat_B[198] +
//             mat_A[935] * mat_B[230] +
//             mat_A[936] * mat_B[262] +
//             mat_A[937] * mat_B[294] +
//             mat_A[938] * mat_B[326] +
//             mat_A[939] * mat_B[358] +
//             mat_A[940] * mat_B[390] +
//             mat_A[941] * mat_B[422] +
//             mat_A[942] * mat_B[454] +
//             mat_A[943] * mat_B[486] +
//             mat_A[944] * mat_B[518] +
//             mat_A[945] * mat_B[550] +
//             mat_A[946] * mat_B[582] +
//             mat_A[947] * mat_B[614] +
//             mat_A[948] * mat_B[646] +
//             mat_A[949] * mat_B[678] +
//             mat_A[950] * mat_B[710] +
//             mat_A[951] * mat_B[742] +
//             mat_A[952] * mat_B[774] +
//             mat_A[953] * mat_B[806] +
//             mat_A[954] * mat_B[838] +
//             mat_A[955] * mat_B[870] +
//             mat_A[956] * mat_B[902] +
//             mat_A[957] * mat_B[934] +
//             mat_A[958] * mat_B[966] +
//             mat_A[959] * mat_B[998];
//  mat_C[935] <= 
//             mat_A[928] * mat_B[7] +
//             mat_A[929] * mat_B[39] +
//             mat_A[930] * mat_B[71] +
//             mat_A[931] * mat_B[103] +
//             mat_A[932] * mat_B[135] +
//             mat_A[933] * mat_B[167] +
//             mat_A[934] * mat_B[199] +
//             mat_A[935] * mat_B[231] +
//             mat_A[936] * mat_B[263] +
//             mat_A[937] * mat_B[295] +
//             mat_A[938] * mat_B[327] +
//             mat_A[939] * mat_B[359] +
//             mat_A[940] * mat_B[391] +
//             mat_A[941] * mat_B[423] +
//             mat_A[942] * mat_B[455] +
//             mat_A[943] * mat_B[487] +
//             mat_A[944] * mat_B[519] +
//             mat_A[945] * mat_B[551] +
//             mat_A[946] * mat_B[583] +
//             mat_A[947] * mat_B[615] +
//             mat_A[948] * mat_B[647] +
//             mat_A[949] * mat_B[679] +
//             mat_A[950] * mat_B[711] +
//             mat_A[951] * mat_B[743] +
//             mat_A[952] * mat_B[775] +
//             mat_A[953] * mat_B[807] +
//             mat_A[954] * mat_B[839] +
//             mat_A[955] * mat_B[871] +
//             mat_A[956] * mat_B[903] +
//             mat_A[957] * mat_B[935] +
//             mat_A[958] * mat_B[967] +
//             mat_A[959] * mat_B[999];
//  mat_C[936] <= 
//             mat_A[928] * mat_B[8] +
//             mat_A[929] * mat_B[40] +
//             mat_A[930] * mat_B[72] +
//             mat_A[931] * mat_B[104] +
//             mat_A[932] * mat_B[136] +
//             mat_A[933] * mat_B[168] +
//             mat_A[934] * mat_B[200] +
//             mat_A[935] * mat_B[232] +
//             mat_A[936] * mat_B[264] +
//             mat_A[937] * mat_B[296] +
//             mat_A[938] * mat_B[328] +
//             mat_A[939] * mat_B[360] +
//             mat_A[940] * mat_B[392] +
//             mat_A[941] * mat_B[424] +
//             mat_A[942] * mat_B[456] +
//             mat_A[943] * mat_B[488] +
//             mat_A[944] * mat_B[520] +
//             mat_A[945] * mat_B[552] +
//             mat_A[946] * mat_B[584] +
//             mat_A[947] * mat_B[616] +
//             mat_A[948] * mat_B[648] +
//             mat_A[949] * mat_B[680] +
//             mat_A[950] * mat_B[712] +
//             mat_A[951] * mat_B[744] +
//             mat_A[952] * mat_B[776] +
//             mat_A[953] * mat_B[808] +
//             mat_A[954] * mat_B[840] +
//             mat_A[955] * mat_B[872] +
//             mat_A[956] * mat_B[904] +
//             mat_A[957] * mat_B[936] +
//             mat_A[958] * mat_B[968] +
//             mat_A[959] * mat_B[1000];
//  mat_C[937] <= 
//             mat_A[928] * mat_B[9] +
//             mat_A[929] * mat_B[41] +
//             mat_A[930] * mat_B[73] +
//             mat_A[931] * mat_B[105] +
//             mat_A[932] * mat_B[137] +
//             mat_A[933] * mat_B[169] +
//             mat_A[934] * mat_B[201] +
//             mat_A[935] * mat_B[233] +
//             mat_A[936] * mat_B[265] +
//             mat_A[937] * mat_B[297] +
//             mat_A[938] * mat_B[329] +
//             mat_A[939] * mat_B[361] +
//             mat_A[940] * mat_B[393] +
//             mat_A[941] * mat_B[425] +
//             mat_A[942] * mat_B[457] +
//             mat_A[943] * mat_B[489] +
//             mat_A[944] * mat_B[521] +
//             mat_A[945] * mat_B[553] +
//             mat_A[946] * mat_B[585] +
//             mat_A[947] * mat_B[617] +
//             mat_A[948] * mat_B[649] +
//             mat_A[949] * mat_B[681] +
//             mat_A[950] * mat_B[713] +
//             mat_A[951] * mat_B[745] +
//             mat_A[952] * mat_B[777] +
//             mat_A[953] * mat_B[809] +
//             mat_A[954] * mat_B[841] +
//             mat_A[955] * mat_B[873] +
//             mat_A[956] * mat_B[905] +
//             mat_A[957] * mat_B[937] +
//             mat_A[958] * mat_B[969] +
//             mat_A[959] * mat_B[1001];
//  mat_C[938] <= 
//             mat_A[928] * mat_B[10] +
//             mat_A[929] * mat_B[42] +
//             mat_A[930] * mat_B[74] +
//             mat_A[931] * mat_B[106] +
//             mat_A[932] * mat_B[138] +
//             mat_A[933] * mat_B[170] +
//             mat_A[934] * mat_B[202] +
//             mat_A[935] * mat_B[234] +
//             mat_A[936] * mat_B[266] +
//             mat_A[937] * mat_B[298] +
//             mat_A[938] * mat_B[330] +
//             mat_A[939] * mat_B[362] +
//             mat_A[940] * mat_B[394] +
//             mat_A[941] * mat_B[426] +
//             mat_A[942] * mat_B[458] +
//             mat_A[943] * mat_B[490] +
//             mat_A[944] * mat_B[522] +
//             mat_A[945] * mat_B[554] +
//             mat_A[946] * mat_B[586] +
//             mat_A[947] * mat_B[618] +
//             mat_A[948] * mat_B[650] +
//             mat_A[949] * mat_B[682] +
//             mat_A[950] * mat_B[714] +
//             mat_A[951] * mat_B[746] +
//             mat_A[952] * mat_B[778] +
//             mat_A[953] * mat_B[810] +
//             mat_A[954] * mat_B[842] +
//             mat_A[955] * mat_B[874] +
//             mat_A[956] * mat_B[906] +
//             mat_A[957] * mat_B[938] +
//             mat_A[958] * mat_B[970] +
//             mat_A[959] * mat_B[1002];
//  mat_C[939] <= 
//             mat_A[928] * mat_B[11] +
//             mat_A[929] * mat_B[43] +
//             mat_A[930] * mat_B[75] +
//             mat_A[931] * mat_B[107] +
//             mat_A[932] * mat_B[139] +
//             mat_A[933] * mat_B[171] +
//             mat_A[934] * mat_B[203] +
//             mat_A[935] * mat_B[235] +
//             mat_A[936] * mat_B[267] +
//             mat_A[937] * mat_B[299] +
//             mat_A[938] * mat_B[331] +
//             mat_A[939] * mat_B[363] +
//             mat_A[940] * mat_B[395] +
//             mat_A[941] * mat_B[427] +
//             mat_A[942] * mat_B[459] +
//             mat_A[943] * mat_B[491] +
//             mat_A[944] * mat_B[523] +
//             mat_A[945] * mat_B[555] +
//             mat_A[946] * mat_B[587] +
//             mat_A[947] * mat_B[619] +
//             mat_A[948] * mat_B[651] +
//             mat_A[949] * mat_B[683] +
//             mat_A[950] * mat_B[715] +
//             mat_A[951] * mat_B[747] +
//             mat_A[952] * mat_B[779] +
//             mat_A[953] * mat_B[811] +
//             mat_A[954] * mat_B[843] +
//             mat_A[955] * mat_B[875] +
//             mat_A[956] * mat_B[907] +
//             mat_A[957] * mat_B[939] +
//             mat_A[958] * mat_B[971] +
//             mat_A[959] * mat_B[1003];
//  mat_C[940] <= 
//             mat_A[928] * mat_B[12] +
//             mat_A[929] * mat_B[44] +
//             mat_A[930] * mat_B[76] +
//             mat_A[931] * mat_B[108] +
//             mat_A[932] * mat_B[140] +
//             mat_A[933] * mat_B[172] +
//             mat_A[934] * mat_B[204] +
//             mat_A[935] * mat_B[236] +
//             mat_A[936] * mat_B[268] +
//             mat_A[937] * mat_B[300] +
//             mat_A[938] * mat_B[332] +
//             mat_A[939] * mat_B[364] +
//             mat_A[940] * mat_B[396] +
//             mat_A[941] * mat_B[428] +
//             mat_A[942] * mat_B[460] +
//             mat_A[943] * mat_B[492] +
//             mat_A[944] * mat_B[524] +
//             mat_A[945] * mat_B[556] +
//             mat_A[946] * mat_B[588] +
//             mat_A[947] * mat_B[620] +
//             mat_A[948] * mat_B[652] +
//             mat_A[949] * mat_B[684] +
//             mat_A[950] * mat_B[716] +
//             mat_A[951] * mat_B[748] +
//             mat_A[952] * mat_B[780] +
//             mat_A[953] * mat_B[812] +
//             mat_A[954] * mat_B[844] +
//             mat_A[955] * mat_B[876] +
//             mat_A[956] * mat_B[908] +
//             mat_A[957] * mat_B[940] +
//             mat_A[958] * mat_B[972] +
//             mat_A[959] * mat_B[1004];
//  mat_C[941] <= 
//             mat_A[928] * mat_B[13] +
//             mat_A[929] * mat_B[45] +
//             mat_A[930] * mat_B[77] +
//             mat_A[931] * mat_B[109] +
//             mat_A[932] * mat_B[141] +
//             mat_A[933] * mat_B[173] +
//             mat_A[934] * mat_B[205] +
//             mat_A[935] * mat_B[237] +
//             mat_A[936] * mat_B[269] +
//             mat_A[937] * mat_B[301] +
//             mat_A[938] * mat_B[333] +
//             mat_A[939] * mat_B[365] +
//             mat_A[940] * mat_B[397] +
//             mat_A[941] * mat_B[429] +
//             mat_A[942] * mat_B[461] +
//             mat_A[943] * mat_B[493] +
//             mat_A[944] * mat_B[525] +
//             mat_A[945] * mat_B[557] +
//             mat_A[946] * mat_B[589] +
//             mat_A[947] * mat_B[621] +
//             mat_A[948] * mat_B[653] +
//             mat_A[949] * mat_B[685] +
//             mat_A[950] * mat_B[717] +
//             mat_A[951] * mat_B[749] +
//             mat_A[952] * mat_B[781] +
//             mat_A[953] * mat_B[813] +
//             mat_A[954] * mat_B[845] +
//             mat_A[955] * mat_B[877] +
//             mat_A[956] * mat_B[909] +
//             mat_A[957] * mat_B[941] +
//             mat_A[958] * mat_B[973] +
//             mat_A[959] * mat_B[1005];
//  mat_C[942] <= 
//             mat_A[928] * mat_B[14] +
//             mat_A[929] * mat_B[46] +
//             mat_A[930] * mat_B[78] +
//             mat_A[931] * mat_B[110] +
//             mat_A[932] * mat_B[142] +
//             mat_A[933] * mat_B[174] +
//             mat_A[934] * mat_B[206] +
//             mat_A[935] * mat_B[238] +
//             mat_A[936] * mat_B[270] +
//             mat_A[937] * mat_B[302] +
//             mat_A[938] * mat_B[334] +
//             mat_A[939] * mat_B[366] +
//             mat_A[940] * mat_B[398] +
//             mat_A[941] * mat_B[430] +
//             mat_A[942] * mat_B[462] +
//             mat_A[943] * mat_B[494] +
//             mat_A[944] * mat_B[526] +
//             mat_A[945] * mat_B[558] +
//             mat_A[946] * mat_B[590] +
//             mat_A[947] * mat_B[622] +
//             mat_A[948] * mat_B[654] +
//             mat_A[949] * mat_B[686] +
//             mat_A[950] * mat_B[718] +
//             mat_A[951] * mat_B[750] +
//             mat_A[952] * mat_B[782] +
//             mat_A[953] * mat_B[814] +
//             mat_A[954] * mat_B[846] +
//             mat_A[955] * mat_B[878] +
//             mat_A[956] * mat_B[910] +
//             mat_A[957] * mat_B[942] +
//             mat_A[958] * mat_B[974] +
//             mat_A[959] * mat_B[1006];
//  mat_C[943] <= 
//             mat_A[928] * mat_B[15] +
//             mat_A[929] * mat_B[47] +
//             mat_A[930] * mat_B[79] +
//             mat_A[931] * mat_B[111] +
//             mat_A[932] * mat_B[143] +
//             mat_A[933] * mat_B[175] +
//             mat_A[934] * mat_B[207] +
//             mat_A[935] * mat_B[239] +
//             mat_A[936] * mat_B[271] +
//             mat_A[937] * mat_B[303] +
//             mat_A[938] * mat_B[335] +
//             mat_A[939] * mat_B[367] +
//             mat_A[940] * mat_B[399] +
//             mat_A[941] * mat_B[431] +
//             mat_A[942] * mat_B[463] +
//             mat_A[943] * mat_B[495] +
//             mat_A[944] * mat_B[527] +
//             mat_A[945] * mat_B[559] +
//             mat_A[946] * mat_B[591] +
//             mat_A[947] * mat_B[623] +
//             mat_A[948] * mat_B[655] +
//             mat_A[949] * mat_B[687] +
//             mat_A[950] * mat_B[719] +
//             mat_A[951] * mat_B[751] +
//             mat_A[952] * mat_B[783] +
//             mat_A[953] * mat_B[815] +
//             mat_A[954] * mat_B[847] +
//             mat_A[955] * mat_B[879] +
//             mat_A[956] * mat_B[911] +
//             mat_A[957] * mat_B[943] +
//             mat_A[958] * mat_B[975] +
//             mat_A[959] * mat_B[1007];
//  mat_C[944] <= 
//             mat_A[928] * mat_B[16] +
//             mat_A[929] * mat_B[48] +
//             mat_A[930] * mat_B[80] +
//             mat_A[931] * mat_B[112] +
//             mat_A[932] * mat_B[144] +
//             mat_A[933] * mat_B[176] +
//             mat_A[934] * mat_B[208] +
//             mat_A[935] * mat_B[240] +
//             mat_A[936] * mat_B[272] +
//             mat_A[937] * mat_B[304] +
//             mat_A[938] * mat_B[336] +
//             mat_A[939] * mat_B[368] +
//             mat_A[940] * mat_B[400] +
//             mat_A[941] * mat_B[432] +
//             mat_A[942] * mat_B[464] +
//             mat_A[943] * mat_B[496] +
//             mat_A[944] * mat_B[528] +
//             mat_A[945] * mat_B[560] +
//             mat_A[946] * mat_B[592] +
//             mat_A[947] * mat_B[624] +
//             mat_A[948] * mat_B[656] +
//             mat_A[949] * mat_B[688] +
//             mat_A[950] * mat_B[720] +
//             mat_A[951] * mat_B[752] +
//             mat_A[952] * mat_B[784] +
//             mat_A[953] * mat_B[816] +
//             mat_A[954] * mat_B[848] +
//             mat_A[955] * mat_B[880] +
//             mat_A[956] * mat_B[912] +
//             mat_A[957] * mat_B[944] +
//             mat_A[958] * mat_B[976] +
//             mat_A[959] * mat_B[1008];
//  mat_C[945] <= 
//             mat_A[928] * mat_B[17] +
//             mat_A[929] * mat_B[49] +
//             mat_A[930] * mat_B[81] +
//             mat_A[931] * mat_B[113] +
//             mat_A[932] * mat_B[145] +
//             mat_A[933] * mat_B[177] +
//             mat_A[934] * mat_B[209] +
//             mat_A[935] * mat_B[241] +
//             mat_A[936] * mat_B[273] +
//             mat_A[937] * mat_B[305] +
//             mat_A[938] * mat_B[337] +
//             mat_A[939] * mat_B[369] +
//             mat_A[940] * mat_B[401] +
//             mat_A[941] * mat_B[433] +
//             mat_A[942] * mat_B[465] +
//             mat_A[943] * mat_B[497] +
//             mat_A[944] * mat_B[529] +
//             mat_A[945] * mat_B[561] +
//             mat_A[946] * mat_B[593] +
//             mat_A[947] * mat_B[625] +
//             mat_A[948] * mat_B[657] +
//             mat_A[949] * mat_B[689] +
//             mat_A[950] * mat_B[721] +
//             mat_A[951] * mat_B[753] +
//             mat_A[952] * mat_B[785] +
//             mat_A[953] * mat_B[817] +
//             mat_A[954] * mat_B[849] +
//             mat_A[955] * mat_B[881] +
//             mat_A[956] * mat_B[913] +
//             mat_A[957] * mat_B[945] +
//             mat_A[958] * mat_B[977] +
//             mat_A[959] * mat_B[1009];
//  mat_C[946] <= 
//             mat_A[928] * mat_B[18] +
//             mat_A[929] * mat_B[50] +
//             mat_A[930] * mat_B[82] +
//             mat_A[931] * mat_B[114] +
//             mat_A[932] * mat_B[146] +
//             mat_A[933] * mat_B[178] +
//             mat_A[934] * mat_B[210] +
//             mat_A[935] * mat_B[242] +
//             mat_A[936] * mat_B[274] +
//             mat_A[937] * mat_B[306] +
//             mat_A[938] * mat_B[338] +
//             mat_A[939] * mat_B[370] +
//             mat_A[940] * mat_B[402] +
//             mat_A[941] * mat_B[434] +
//             mat_A[942] * mat_B[466] +
//             mat_A[943] * mat_B[498] +
//             mat_A[944] * mat_B[530] +
//             mat_A[945] * mat_B[562] +
//             mat_A[946] * mat_B[594] +
//             mat_A[947] * mat_B[626] +
//             mat_A[948] * mat_B[658] +
//             mat_A[949] * mat_B[690] +
//             mat_A[950] * mat_B[722] +
//             mat_A[951] * mat_B[754] +
//             mat_A[952] * mat_B[786] +
//             mat_A[953] * mat_B[818] +
//             mat_A[954] * mat_B[850] +
//             mat_A[955] * mat_B[882] +
//             mat_A[956] * mat_B[914] +
//             mat_A[957] * mat_B[946] +
//             mat_A[958] * mat_B[978] +
//             mat_A[959] * mat_B[1010];
//  mat_C[947] <= 
//             mat_A[928] * mat_B[19] +
//             mat_A[929] * mat_B[51] +
//             mat_A[930] * mat_B[83] +
//             mat_A[931] * mat_B[115] +
//             mat_A[932] * mat_B[147] +
//             mat_A[933] * mat_B[179] +
//             mat_A[934] * mat_B[211] +
//             mat_A[935] * mat_B[243] +
//             mat_A[936] * mat_B[275] +
//             mat_A[937] * mat_B[307] +
//             mat_A[938] * mat_B[339] +
//             mat_A[939] * mat_B[371] +
//             mat_A[940] * mat_B[403] +
//             mat_A[941] * mat_B[435] +
//             mat_A[942] * mat_B[467] +
//             mat_A[943] * mat_B[499] +
//             mat_A[944] * mat_B[531] +
//             mat_A[945] * mat_B[563] +
//             mat_A[946] * mat_B[595] +
//             mat_A[947] * mat_B[627] +
//             mat_A[948] * mat_B[659] +
//             mat_A[949] * mat_B[691] +
//             mat_A[950] * mat_B[723] +
//             mat_A[951] * mat_B[755] +
//             mat_A[952] * mat_B[787] +
//             mat_A[953] * mat_B[819] +
//             mat_A[954] * mat_B[851] +
//             mat_A[955] * mat_B[883] +
//             mat_A[956] * mat_B[915] +
//             mat_A[957] * mat_B[947] +
//             mat_A[958] * mat_B[979] +
//             mat_A[959] * mat_B[1011];
//  mat_C[948] <= 
//             mat_A[928] * mat_B[20] +
//             mat_A[929] * mat_B[52] +
//             mat_A[930] * mat_B[84] +
//             mat_A[931] * mat_B[116] +
//             mat_A[932] * mat_B[148] +
//             mat_A[933] * mat_B[180] +
//             mat_A[934] * mat_B[212] +
//             mat_A[935] * mat_B[244] +
//             mat_A[936] * mat_B[276] +
//             mat_A[937] * mat_B[308] +
//             mat_A[938] * mat_B[340] +
//             mat_A[939] * mat_B[372] +
//             mat_A[940] * mat_B[404] +
//             mat_A[941] * mat_B[436] +
//             mat_A[942] * mat_B[468] +
//             mat_A[943] * mat_B[500] +
//             mat_A[944] * mat_B[532] +
//             mat_A[945] * mat_B[564] +
//             mat_A[946] * mat_B[596] +
//             mat_A[947] * mat_B[628] +
//             mat_A[948] * mat_B[660] +
//             mat_A[949] * mat_B[692] +
//             mat_A[950] * mat_B[724] +
//             mat_A[951] * mat_B[756] +
//             mat_A[952] * mat_B[788] +
//             mat_A[953] * mat_B[820] +
//             mat_A[954] * mat_B[852] +
//             mat_A[955] * mat_B[884] +
//             mat_A[956] * mat_B[916] +
//             mat_A[957] * mat_B[948] +
//             mat_A[958] * mat_B[980] +
//             mat_A[959] * mat_B[1012];
//  mat_C[949] <= 
//             mat_A[928] * mat_B[21] +
//             mat_A[929] * mat_B[53] +
//             mat_A[930] * mat_B[85] +
//             mat_A[931] * mat_B[117] +
//             mat_A[932] * mat_B[149] +
//             mat_A[933] * mat_B[181] +
//             mat_A[934] * mat_B[213] +
//             mat_A[935] * mat_B[245] +
//             mat_A[936] * mat_B[277] +
//             mat_A[937] * mat_B[309] +
//             mat_A[938] * mat_B[341] +
//             mat_A[939] * mat_B[373] +
//             mat_A[940] * mat_B[405] +
//             mat_A[941] * mat_B[437] +
//             mat_A[942] * mat_B[469] +
//             mat_A[943] * mat_B[501] +
//             mat_A[944] * mat_B[533] +
//             mat_A[945] * mat_B[565] +
//             mat_A[946] * mat_B[597] +
//             mat_A[947] * mat_B[629] +
//             mat_A[948] * mat_B[661] +
//             mat_A[949] * mat_B[693] +
//             mat_A[950] * mat_B[725] +
//             mat_A[951] * mat_B[757] +
//             mat_A[952] * mat_B[789] +
//             mat_A[953] * mat_B[821] +
//             mat_A[954] * mat_B[853] +
//             mat_A[955] * mat_B[885] +
//             mat_A[956] * mat_B[917] +
//             mat_A[957] * mat_B[949] +
//             mat_A[958] * mat_B[981] +
//             mat_A[959] * mat_B[1013];
//  mat_C[950] <= 
//             mat_A[928] * mat_B[22] +
//             mat_A[929] * mat_B[54] +
//             mat_A[930] * mat_B[86] +
//             mat_A[931] * mat_B[118] +
//             mat_A[932] * mat_B[150] +
//             mat_A[933] * mat_B[182] +
//             mat_A[934] * mat_B[214] +
//             mat_A[935] * mat_B[246] +
//             mat_A[936] * mat_B[278] +
//             mat_A[937] * mat_B[310] +
//             mat_A[938] * mat_B[342] +
//             mat_A[939] * mat_B[374] +
//             mat_A[940] * mat_B[406] +
//             mat_A[941] * mat_B[438] +
//             mat_A[942] * mat_B[470] +
//             mat_A[943] * mat_B[502] +
//             mat_A[944] * mat_B[534] +
//             mat_A[945] * mat_B[566] +
//             mat_A[946] * mat_B[598] +
//             mat_A[947] * mat_B[630] +
//             mat_A[948] * mat_B[662] +
//             mat_A[949] * mat_B[694] +
//             mat_A[950] * mat_B[726] +
//             mat_A[951] * mat_B[758] +
//             mat_A[952] * mat_B[790] +
//             mat_A[953] * mat_B[822] +
//             mat_A[954] * mat_B[854] +
//             mat_A[955] * mat_B[886] +
//             mat_A[956] * mat_B[918] +
//             mat_A[957] * mat_B[950] +
//             mat_A[958] * mat_B[982] +
//             mat_A[959] * mat_B[1014];
//  mat_C[951] <= 
//             mat_A[928] * mat_B[23] +
//             mat_A[929] * mat_B[55] +
//             mat_A[930] * mat_B[87] +
//             mat_A[931] * mat_B[119] +
//             mat_A[932] * mat_B[151] +
//             mat_A[933] * mat_B[183] +
//             mat_A[934] * mat_B[215] +
//             mat_A[935] * mat_B[247] +
//             mat_A[936] * mat_B[279] +
//             mat_A[937] * mat_B[311] +
//             mat_A[938] * mat_B[343] +
//             mat_A[939] * mat_B[375] +
//             mat_A[940] * mat_B[407] +
//             mat_A[941] * mat_B[439] +
//             mat_A[942] * mat_B[471] +
//             mat_A[943] * mat_B[503] +
//             mat_A[944] * mat_B[535] +
//             mat_A[945] * mat_B[567] +
//             mat_A[946] * mat_B[599] +
//             mat_A[947] * mat_B[631] +
//             mat_A[948] * mat_B[663] +
//             mat_A[949] * mat_B[695] +
//             mat_A[950] * mat_B[727] +
//             mat_A[951] * mat_B[759] +
//             mat_A[952] * mat_B[791] +
//             mat_A[953] * mat_B[823] +
//             mat_A[954] * mat_B[855] +
//             mat_A[955] * mat_B[887] +
//             mat_A[956] * mat_B[919] +
//             mat_A[957] * mat_B[951] +
//             mat_A[958] * mat_B[983] +
//             mat_A[959] * mat_B[1015];
//  mat_C[952] <= 
//             mat_A[928] * mat_B[24] +
//             mat_A[929] * mat_B[56] +
//             mat_A[930] * mat_B[88] +
//             mat_A[931] * mat_B[120] +
//             mat_A[932] * mat_B[152] +
//             mat_A[933] * mat_B[184] +
//             mat_A[934] * mat_B[216] +
//             mat_A[935] * mat_B[248] +
//             mat_A[936] * mat_B[280] +
//             mat_A[937] * mat_B[312] +
//             mat_A[938] * mat_B[344] +
//             mat_A[939] * mat_B[376] +
//             mat_A[940] * mat_B[408] +
//             mat_A[941] * mat_B[440] +
//             mat_A[942] * mat_B[472] +
//             mat_A[943] * mat_B[504] +
//             mat_A[944] * mat_B[536] +
//             mat_A[945] * mat_B[568] +
//             mat_A[946] * mat_B[600] +
//             mat_A[947] * mat_B[632] +
//             mat_A[948] * mat_B[664] +
//             mat_A[949] * mat_B[696] +
//             mat_A[950] * mat_B[728] +
//             mat_A[951] * mat_B[760] +
//             mat_A[952] * mat_B[792] +
//             mat_A[953] * mat_B[824] +
//             mat_A[954] * mat_B[856] +
//             mat_A[955] * mat_B[888] +
//             mat_A[956] * mat_B[920] +
//             mat_A[957] * mat_B[952] +
//             mat_A[958] * mat_B[984] +
//             mat_A[959] * mat_B[1016];
//  mat_C[953] <= 
//             mat_A[928] * mat_B[25] +
//             mat_A[929] * mat_B[57] +
//             mat_A[930] * mat_B[89] +
//             mat_A[931] * mat_B[121] +
//             mat_A[932] * mat_B[153] +
//             mat_A[933] * mat_B[185] +
//             mat_A[934] * mat_B[217] +
//             mat_A[935] * mat_B[249] +
//             mat_A[936] * mat_B[281] +
//             mat_A[937] * mat_B[313] +
//             mat_A[938] * mat_B[345] +
//             mat_A[939] * mat_B[377] +
//             mat_A[940] * mat_B[409] +
//             mat_A[941] * mat_B[441] +
//             mat_A[942] * mat_B[473] +
//             mat_A[943] * mat_B[505] +
//             mat_A[944] * mat_B[537] +
//             mat_A[945] * mat_B[569] +
//             mat_A[946] * mat_B[601] +
//             mat_A[947] * mat_B[633] +
//             mat_A[948] * mat_B[665] +
//             mat_A[949] * mat_B[697] +
//             mat_A[950] * mat_B[729] +
//             mat_A[951] * mat_B[761] +
//             mat_A[952] * mat_B[793] +
//             mat_A[953] * mat_B[825] +
//             mat_A[954] * mat_B[857] +
//             mat_A[955] * mat_B[889] +
//             mat_A[956] * mat_B[921] +
//             mat_A[957] * mat_B[953] +
//             mat_A[958] * mat_B[985] +
//             mat_A[959] * mat_B[1017];
//  mat_C[954] <= 
//             mat_A[928] * mat_B[26] +
//             mat_A[929] * mat_B[58] +
//             mat_A[930] * mat_B[90] +
//             mat_A[931] * mat_B[122] +
//             mat_A[932] * mat_B[154] +
//             mat_A[933] * mat_B[186] +
//             mat_A[934] * mat_B[218] +
//             mat_A[935] * mat_B[250] +
//             mat_A[936] * mat_B[282] +
//             mat_A[937] * mat_B[314] +
//             mat_A[938] * mat_B[346] +
//             mat_A[939] * mat_B[378] +
//             mat_A[940] * mat_B[410] +
//             mat_A[941] * mat_B[442] +
//             mat_A[942] * mat_B[474] +
//             mat_A[943] * mat_B[506] +
//             mat_A[944] * mat_B[538] +
//             mat_A[945] * mat_B[570] +
//             mat_A[946] * mat_B[602] +
//             mat_A[947] * mat_B[634] +
//             mat_A[948] * mat_B[666] +
//             mat_A[949] * mat_B[698] +
//             mat_A[950] * mat_B[730] +
//             mat_A[951] * mat_B[762] +
//             mat_A[952] * mat_B[794] +
//             mat_A[953] * mat_B[826] +
//             mat_A[954] * mat_B[858] +
//             mat_A[955] * mat_B[890] +
//             mat_A[956] * mat_B[922] +
//             mat_A[957] * mat_B[954] +
//             mat_A[958] * mat_B[986] +
//             mat_A[959] * mat_B[1018];
//  mat_C[955] <= 
//             mat_A[928] * mat_B[27] +
//             mat_A[929] * mat_B[59] +
//             mat_A[930] * mat_B[91] +
//             mat_A[931] * mat_B[123] +
//             mat_A[932] * mat_B[155] +
//             mat_A[933] * mat_B[187] +
//             mat_A[934] * mat_B[219] +
//             mat_A[935] * mat_B[251] +
//             mat_A[936] * mat_B[283] +
//             mat_A[937] * mat_B[315] +
//             mat_A[938] * mat_B[347] +
//             mat_A[939] * mat_B[379] +
//             mat_A[940] * mat_B[411] +
//             mat_A[941] * mat_B[443] +
//             mat_A[942] * mat_B[475] +
//             mat_A[943] * mat_B[507] +
//             mat_A[944] * mat_B[539] +
//             mat_A[945] * mat_B[571] +
//             mat_A[946] * mat_B[603] +
//             mat_A[947] * mat_B[635] +
//             mat_A[948] * mat_B[667] +
//             mat_A[949] * mat_B[699] +
//             mat_A[950] * mat_B[731] +
//             mat_A[951] * mat_B[763] +
//             mat_A[952] * mat_B[795] +
//             mat_A[953] * mat_B[827] +
//             mat_A[954] * mat_B[859] +
//             mat_A[955] * mat_B[891] +
//             mat_A[956] * mat_B[923] +
//             mat_A[957] * mat_B[955] +
//             mat_A[958] * mat_B[987] +
//             mat_A[959] * mat_B[1019];
//  mat_C[956] <= 
//             mat_A[928] * mat_B[28] +
//             mat_A[929] * mat_B[60] +
//             mat_A[930] * mat_B[92] +
//             mat_A[931] * mat_B[124] +
//             mat_A[932] * mat_B[156] +
//             mat_A[933] * mat_B[188] +
//             mat_A[934] * mat_B[220] +
//             mat_A[935] * mat_B[252] +
//             mat_A[936] * mat_B[284] +
//             mat_A[937] * mat_B[316] +
//             mat_A[938] * mat_B[348] +
//             mat_A[939] * mat_B[380] +
//             mat_A[940] * mat_B[412] +
//             mat_A[941] * mat_B[444] +
//             mat_A[942] * mat_B[476] +
//             mat_A[943] * mat_B[508] +
//             mat_A[944] * mat_B[540] +
//             mat_A[945] * mat_B[572] +
//             mat_A[946] * mat_B[604] +
//             mat_A[947] * mat_B[636] +
//             mat_A[948] * mat_B[668] +
//             mat_A[949] * mat_B[700] +
//             mat_A[950] * mat_B[732] +
//             mat_A[951] * mat_B[764] +
//             mat_A[952] * mat_B[796] +
//             mat_A[953] * mat_B[828] +
//             mat_A[954] * mat_B[860] +
//             mat_A[955] * mat_B[892] +
//             mat_A[956] * mat_B[924] +
//             mat_A[957] * mat_B[956] +
//             mat_A[958] * mat_B[988] +
//             mat_A[959] * mat_B[1020];
//  mat_C[957] <= 
//             mat_A[928] * mat_B[29] +
//             mat_A[929] * mat_B[61] +
//             mat_A[930] * mat_B[93] +
//             mat_A[931] * mat_B[125] +
//             mat_A[932] * mat_B[157] +
//             mat_A[933] * mat_B[189] +
//             mat_A[934] * mat_B[221] +
//             mat_A[935] * mat_B[253] +
//             mat_A[936] * mat_B[285] +
//             mat_A[937] * mat_B[317] +
//             mat_A[938] * mat_B[349] +
//             mat_A[939] * mat_B[381] +
//             mat_A[940] * mat_B[413] +
//             mat_A[941] * mat_B[445] +
//             mat_A[942] * mat_B[477] +
//             mat_A[943] * mat_B[509] +
//             mat_A[944] * mat_B[541] +
//             mat_A[945] * mat_B[573] +
//             mat_A[946] * mat_B[605] +
//             mat_A[947] * mat_B[637] +
//             mat_A[948] * mat_B[669] +
//             mat_A[949] * mat_B[701] +
//             mat_A[950] * mat_B[733] +
//             mat_A[951] * mat_B[765] +
//             mat_A[952] * mat_B[797] +
//             mat_A[953] * mat_B[829] +
//             mat_A[954] * mat_B[861] +
//             mat_A[955] * mat_B[893] +
//             mat_A[956] * mat_B[925] +
//             mat_A[957] * mat_B[957] +
//             mat_A[958] * mat_B[989] +
//             mat_A[959] * mat_B[1021];
//  mat_C[958] <= 
//             mat_A[928] * mat_B[30] +
//             mat_A[929] * mat_B[62] +
//             mat_A[930] * mat_B[94] +
//             mat_A[931] * mat_B[126] +
//             mat_A[932] * mat_B[158] +
//             mat_A[933] * mat_B[190] +
//             mat_A[934] * mat_B[222] +
//             mat_A[935] * mat_B[254] +
//             mat_A[936] * mat_B[286] +
//             mat_A[937] * mat_B[318] +
//             mat_A[938] * mat_B[350] +
//             mat_A[939] * mat_B[382] +
//             mat_A[940] * mat_B[414] +
//             mat_A[941] * mat_B[446] +
//             mat_A[942] * mat_B[478] +
//             mat_A[943] * mat_B[510] +
//             mat_A[944] * mat_B[542] +
//             mat_A[945] * mat_B[574] +
//             mat_A[946] * mat_B[606] +
//             mat_A[947] * mat_B[638] +
//             mat_A[948] * mat_B[670] +
//             mat_A[949] * mat_B[702] +
//             mat_A[950] * mat_B[734] +
//             mat_A[951] * mat_B[766] +
//             mat_A[952] * mat_B[798] +
//             mat_A[953] * mat_B[830] +
//             mat_A[954] * mat_B[862] +
//             mat_A[955] * mat_B[894] +
//             mat_A[956] * mat_B[926] +
//             mat_A[957] * mat_B[958] +
//             mat_A[958] * mat_B[990] +
//             mat_A[959] * mat_B[1022];
//  mat_C[959] <= 
//             mat_A[928] * mat_B[31] +
//             mat_A[929] * mat_B[63] +
//             mat_A[930] * mat_B[95] +
//             mat_A[931] * mat_B[127] +
//             mat_A[932] * mat_B[159] +
//             mat_A[933] * mat_B[191] +
//             mat_A[934] * mat_B[223] +
//             mat_A[935] * mat_B[255] +
//             mat_A[936] * mat_B[287] +
//             mat_A[937] * mat_B[319] +
//             mat_A[938] * mat_B[351] +
//             mat_A[939] * mat_B[383] +
//             mat_A[940] * mat_B[415] +
//             mat_A[941] * mat_B[447] +
//             mat_A[942] * mat_B[479] +
//             mat_A[943] * mat_B[511] +
//             mat_A[944] * mat_B[543] +
//             mat_A[945] * mat_B[575] +
//             mat_A[946] * mat_B[607] +
//             mat_A[947] * mat_B[639] +
//             mat_A[948] * mat_B[671] +
//             mat_A[949] * mat_B[703] +
//             mat_A[950] * mat_B[735] +
//             mat_A[951] * mat_B[767] +
//             mat_A[952] * mat_B[799] +
//             mat_A[953] * mat_B[831] +
//             mat_A[954] * mat_B[863] +
//             mat_A[955] * mat_B[895] +
//             mat_A[956] * mat_B[927] +
//             mat_A[957] * mat_B[959] +
//             mat_A[958] * mat_B[991] +
//             mat_A[959] * mat_B[1023];
//  mat_C[960] <= 
//             mat_A[960] * mat_B[0] +
//             mat_A[961] * mat_B[32] +
//             mat_A[962] * mat_B[64] +
//             mat_A[963] * mat_B[96] +
//             mat_A[964] * mat_B[128] +
//             mat_A[965] * mat_B[160] +
//             mat_A[966] * mat_B[192] +
//             mat_A[967] * mat_B[224] +
//             mat_A[968] * mat_B[256] +
//             mat_A[969] * mat_B[288] +
//             mat_A[970] * mat_B[320] +
//             mat_A[971] * mat_B[352] +
//             mat_A[972] * mat_B[384] +
//             mat_A[973] * mat_B[416] +
//             mat_A[974] * mat_B[448] +
//             mat_A[975] * mat_B[480] +
//             mat_A[976] * mat_B[512] +
//             mat_A[977] * mat_B[544] +
//             mat_A[978] * mat_B[576] +
//             mat_A[979] * mat_B[608] +
//             mat_A[980] * mat_B[640] +
//             mat_A[981] * mat_B[672] +
//             mat_A[982] * mat_B[704] +
//             mat_A[983] * mat_B[736] +
//             mat_A[984] * mat_B[768] +
//             mat_A[985] * mat_B[800] +
//             mat_A[986] * mat_B[832] +
//             mat_A[987] * mat_B[864] +
//             mat_A[988] * mat_B[896] +
//             mat_A[989] * mat_B[928] +
//             mat_A[990] * mat_B[960] +
//             mat_A[991] * mat_B[992];
//  mat_C[961] <= 
//             mat_A[960] * mat_B[1] +
//             mat_A[961] * mat_B[33] +
//             mat_A[962] * mat_B[65] +
//             mat_A[963] * mat_B[97] +
//             mat_A[964] * mat_B[129] +
//             mat_A[965] * mat_B[161] +
//             mat_A[966] * mat_B[193] +
//             mat_A[967] * mat_B[225] +
//             mat_A[968] * mat_B[257] +
//             mat_A[969] * mat_B[289] +
//             mat_A[970] * mat_B[321] +
//             mat_A[971] * mat_B[353] +
//             mat_A[972] * mat_B[385] +
//             mat_A[973] * mat_B[417] +
//             mat_A[974] * mat_B[449] +
//             mat_A[975] * mat_B[481] +
//             mat_A[976] * mat_B[513] +
//             mat_A[977] * mat_B[545] +
//             mat_A[978] * mat_B[577] +
//             mat_A[979] * mat_B[609] +
//             mat_A[980] * mat_B[641] +
//             mat_A[981] * mat_B[673] +
//             mat_A[982] * mat_B[705] +
//             mat_A[983] * mat_B[737] +
//             mat_A[984] * mat_B[769] +
//             mat_A[985] * mat_B[801] +
//             mat_A[986] * mat_B[833] +
//             mat_A[987] * mat_B[865] +
//             mat_A[988] * mat_B[897] +
//             mat_A[989] * mat_B[929] +
//             mat_A[990] * mat_B[961] +
//             mat_A[991] * mat_B[993];
//  mat_C[962] <= 
//             mat_A[960] * mat_B[2] +
//             mat_A[961] * mat_B[34] +
//             mat_A[962] * mat_B[66] +
//             mat_A[963] * mat_B[98] +
//             mat_A[964] * mat_B[130] +
//             mat_A[965] * mat_B[162] +
//             mat_A[966] * mat_B[194] +
//             mat_A[967] * mat_B[226] +
//             mat_A[968] * mat_B[258] +
//             mat_A[969] * mat_B[290] +
//             mat_A[970] * mat_B[322] +
//             mat_A[971] * mat_B[354] +
//             mat_A[972] * mat_B[386] +
//             mat_A[973] * mat_B[418] +
//             mat_A[974] * mat_B[450] +
//             mat_A[975] * mat_B[482] +
//             mat_A[976] * mat_B[514] +
//             mat_A[977] * mat_B[546] +
//             mat_A[978] * mat_B[578] +
//             mat_A[979] * mat_B[610] +
//             mat_A[980] * mat_B[642] +
//             mat_A[981] * mat_B[674] +
//             mat_A[982] * mat_B[706] +
//             mat_A[983] * mat_B[738] +
//             mat_A[984] * mat_B[770] +
//             mat_A[985] * mat_B[802] +
//             mat_A[986] * mat_B[834] +
//             mat_A[987] * mat_B[866] +
//             mat_A[988] * mat_B[898] +
//             mat_A[989] * mat_B[930] +
//             mat_A[990] * mat_B[962] +
//             mat_A[991] * mat_B[994];
//  mat_C[963] <= 
//             mat_A[960] * mat_B[3] +
//             mat_A[961] * mat_B[35] +
//             mat_A[962] * mat_B[67] +
//             mat_A[963] * mat_B[99] +
//             mat_A[964] * mat_B[131] +
//             mat_A[965] * mat_B[163] +
//             mat_A[966] * mat_B[195] +
//             mat_A[967] * mat_B[227] +
//             mat_A[968] * mat_B[259] +
//             mat_A[969] * mat_B[291] +
//             mat_A[970] * mat_B[323] +
//             mat_A[971] * mat_B[355] +
//             mat_A[972] * mat_B[387] +
//             mat_A[973] * mat_B[419] +
//             mat_A[974] * mat_B[451] +
//             mat_A[975] * mat_B[483] +
//             mat_A[976] * mat_B[515] +
//             mat_A[977] * mat_B[547] +
//             mat_A[978] * mat_B[579] +
//             mat_A[979] * mat_B[611] +
//             mat_A[980] * mat_B[643] +
//             mat_A[981] * mat_B[675] +
//             mat_A[982] * mat_B[707] +
//             mat_A[983] * mat_B[739] +
//             mat_A[984] * mat_B[771] +
//             mat_A[985] * mat_B[803] +
//             mat_A[986] * mat_B[835] +
//             mat_A[987] * mat_B[867] +
//             mat_A[988] * mat_B[899] +
//             mat_A[989] * mat_B[931] +
//             mat_A[990] * mat_B[963] +
//             mat_A[991] * mat_B[995];
//  mat_C[964] <= 
//             mat_A[960] * mat_B[4] +
//             mat_A[961] * mat_B[36] +
//             mat_A[962] * mat_B[68] +
//             mat_A[963] * mat_B[100] +
//             mat_A[964] * mat_B[132] +
//             mat_A[965] * mat_B[164] +
//             mat_A[966] * mat_B[196] +
//             mat_A[967] * mat_B[228] +
//             mat_A[968] * mat_B[260] +
//             mat_A[969] * mat_B[292] +
//             mat_A[970] * mat_B[324] +
//             mat_A[971] * mat_B[356] +
//             mat_A[972] * mat_B[388] +
//             mat_A[973] * mat_B[420] +
//             mat_A[974] * mat_B[452] +
//             mat_A[975] * mat_B[484] +
//             mat_A[976] * mat_B[516] +
//             mat_A[977] * mat_B[548] +
//             mat_A[978] * mat_B[580] +
//             mat_A[979] * mat_B[612] +
//             mat_A[980] * mat_B[644] +
//             mat_A[981] * mat_B[676] +
//             mat_A[982] * mat_B[708] +
//             mat_A[983] * mat_B[740] +
//             mat_A[984] * mat_B[772] +
//             mat_A[985] * mat_B[804] +
//             mat_A[986] * mat_B[836] +
//             mat_A[987] * mat_B[868] +
//             mat_A[988] * mat_B[900] +
//             mat_A[989] * mat_B[932] +
//             mat_A[990] * mat_B[964] +
//             mat_A[991] * mat_B[996];
//  mat_C[965] <= 
//             mat_A[960] * mat_B[5] +
//             mat_A[961] * mat_B[37] +
//             mat_A[962] * mat_B[69] +
//             mat_A[963] * mat_B[101] +
//             mat_A[964] * mat_B[133] +
//             mat_A[965] * mat_B[165] +
//             mat_A[966] * mat_B[197] +
//             mat_A[967] * mat_B[229] +
//             mat_A[968] * mat_B[261] +
//             mat_A[969] * mat_B[293] +
//             mat_A[970] * mat_B[325] +
//             mat_A[971] * mat_B[357] +
//             mat_A[972] * mat_B[389] +
//             mat_A[973] * mat_B[421] +
//             mat_A[974] * mat_B[453] +
//             mat_A[975] * mat_B[485] +
//             mat_A[976] * mat_B[517] +
//             mat_A[977] * mat_B[549] +
//             mat_A[978] * mat_B[581] +
//             mat_A[979] * mat_B[613] +
//             mat_A[980] * mat_B[645] +
//             mat_A[981] * mat_B[677] +
//             mat_A[982] * mat_B[709] +
//             mat_A[983] * mat_B[741] +
//             mat_A[984] * mat_B[773] +
//             mat_A[985] * mat_B[805] +
//             mat_A[986] * mat_B[837] +
//             mat_A[987] * mat_B[869] +
//             mat_A[988] * mat_B[901] +
//             mat_A[989] * mat_B[933] +
//             mat_A[990] * mat_B[965] +
//             mat_A[991] * mat_B[997];
//  mat_C[966] <= 
//             mat_A[960] * mat_B[6] +
//             mat_A[961] * mat_B[38] +
//             mat_A[962] * mat_B[70] +
//             mat_A[963] * mat_B[102] +
//             mat_A[964] * mat_B[134] +
//             mat_A[965] * mat_B[166] +
//             mat_A[966] * mat_B[198] +
//             mat_A[967] * mat_B[230] +
//             mat_A[968] * mat_B[262] +
//             mat_A[969] * mat_B[294] +
//             mat_A[970] * mat_B[326] +
//             mat_A[971] * mat_B[358] +
//             mat_A[972] * mat_B[390] +
//             mat_A[973] * mat_B[422] +
//             mat_A[974] * mat_B[454] +
//             mat_A[975] * mat_B[486] +
//             mat_A[976] * mat_B[518] +
//             mat_A[977] * mat_B[550] +
//             mat_A[978] * mat_B[582] +
//             mat_A[979] * mat_B[614] +
//             mat_A[980] * mat_B[646] +
//             mat_A[981] * mat_B[678] +
//             mat_A[982] * mat_B[710] +
//             mat_A[983] * mat_B[742] +
//             mat_A[984] * mat_B[774] +
//             mat_A[985] * mat_B[806] +
//             mat_A[986] * mat_B[838] +
//             mat_A[987] * mat_B[870] +
//             mat_A[988] * mat_B[902] +
//             mat_A[989] * mat_B[934] +
//             mat_A[990] * mat_B[966] +
//             mat_A[991] * mat_B[998];
//  mat_C[967] <= 
//             mat_A[960] * mat_B[7] +
//             mat_A[961] * mat_B[39] +
//             mat_A[962] * mat_B[71] +
//             mat_A[963] * mat_B[103] +
//             mat_A[964] * mat_B[135] +
//             mat_A[965] * mat_B[167] +
//             mat_A[966] * mat_B[199] +
//             mat_A[967] * mat_B[231] +
//             mat_A[968] * mat_B[263] +
//             mat_A[969] * mat_B[295] +
//             mat_A[970] * mat_B[327] +
//             mat_A[971] * mat_B[359] +
//             mat_A[972] * mat_B[391] +
//             mat_A[973] * mat_B[423] +
//             mat_A[974] * mat_B[455] +
//             mat_A[975] * mat_B[487] +
//             mat_A[976] * mat_B[519] +
//             mat_A[977] * mat_B[551] +
//             mat_A[978] * mat_B[583] +
//             mat_A[979] * mat_B[615] +
//             mat_A[980] * mat_B[647] +
//             mat_A[981] * mat_B[679] +
//             mat_A[982] * mat_B[711] +
//             mat_A[983] * mat_B[743] +
//             mat_A[984] * mat_B[775] +
//             mat_A[985] * mat_B[807] +
//             mat_A[986] * mat_B[839] +
//             mat_A[987] * mat_B[871] +
//             mat_A[988] * mat_B[903] +
//             mat_A[989] * mat_B[935] +
//             mat_A[990] * mat_B[967] +
//             mat_A[991] * mat_B[999];
//  mat_C[968] <= 
//             mat_A[960] * mat_B[8] +
//             mat_A[961] * mat_B[40] +
//             mat_A[962] * mat_B[72] +
//             mat_A[963] * mat_B[104] +
//             mat_A[964] * mat_B[136] +
//             mat_A[965] * mat_B[168] +
//             mat_A[966] * mat_B[200] +
//             mat_A[967] * mat_B[232] +
//             mat_A[968] * mat_B[264] +
//             mat_A[969] * mat_B[296] +
//             mat_A[970] * mat_B[328] +
//             mat_A[971] * mat_B[360] +
//             mat_A[972] * mat_B[392] +
//             mat_A[973] * mat_B[424] +
//             mat_A[974] * mat_B[456] +
//             mat_A[975] * mat_B[488] +
//             mat_A[976] * mat_B[520] +
//             mat_A[977] * mat_B[552] +
//             mat_A[978] * mat_B[584] +
//             mat_A[979] * mat_B[616] +
//             mat_A[980] * mat_B[648] +
//             mat_A[981] * mat_B[680] +
//             mat_A[982] * mat_B[712] +
//             mat_A[983] * mat_B[744] +
//             mat_A[984] * mat_B[776] +
//             mat_A[985] * mat_B[808] +
//             mat_A[986] * mat_B[840] +
//             mat_A[987] * mat_B[872] +
//             mat_A[988] * mat_B[904] +
//             mat_A[989] * mat_B[936] +
//             mat_A[990] * mat_B[968] +
//             mat_A[991] * mat_B[1000];
//  mat_C[969] <= 
//             mat_A[960] * mat_B[9] +
//             mat_A[961] * mat_B[41] +
//             mat_A[962] * mat_B[73] +
//             mat_A[963] * mat_B[105] +
//             mat_A[964] * mat_B[137] +
//             mat_A[965] * mat_B[169] +
//             mat_A[966] * mat_B[201] +
//             mat_A[967] * mat_B[233] +
//             mat_A[968] * mat_B[265] +
//             mat_A[969] * mat_B[297] +
//             mat_A[970] * mat_B[329] +
//             mat_A[971] * mat_B[361] +
//             mat_A[972] * mat_B[393] +
//             mat_A[973] * mat_B[425] +
//             mat_A[974] * mat_B[457] +
//             mat_A[975] * mat_B[489] +
//             mat_A[976] * mat_B[521] +
//             mat_A[977] * mat_B[553] +
//             mat_A[978] * mat_B[585] +
//             mat_A[979] * mat_B[617] +
//             mat_A[980] * mat_B[649] +
//             mat_A[981] * mat_B[681] +
//             mat_A[982] * mat_B[713] +
//             mat_A[983] * mat_B[745] +
//             mat_A[984] * mat_B[777] +
//             mat_A[985] * mat_B[809] +
//             mat_A[986] * mat_B[841] +
//             mat_A[987] * mat_B[873] +
//             mat_A[988] * mat_B[905] +
//             mat_A[989] * mat_B[937] +
//             mat_A[990] * mat_B[969] +
//             mat_A[991] * mat_B[1001];
//  mat_C[970] <= 
//             mat_A[960] * mat_B[10] +
//             mat_A[961] * mat_B[42] +
//             mat_A[962] * mat_B[74] +
//             mat_A[963] * mat_B[106] +
//             mat_A[964] * mat_B[138] +
//             mat_A[965] * mat_B[170] +
//             mat_A[966] * mat_B[202] +
//             mat_A[967] * mat_B[234] +
//             mat_A[968] * mat_B[266] +
//             mat_A[969] * mat_B[298] +
//             mat_A[970] * mat_B[330] +
//             mat_A[971] * mat_B[362] +
//             mat_A[972] * mat_B[394] +
//             mat_A[973] * mat_B[426] +
//             mat_A[974] * mat_B[458] +
//             mat_A[975] * mat_B[490] +
//             mat_A[976] * mat_B[522] +
//             mat_A[977] * mat_B[554] +
//             mat_A[978] * mat_B[586] +
//             mat_A[979] * mat_B[618] +
//             mat_A[980] * mat_B[650] +
//             mat_A[981] * mat_B[682] +
//             mat_A[982] * mat_B[714] +
//             mat_A[983] * mat_B[746] +
//             mat_A[984] * mat_B[778] +
//             mat_A[985] * mat_B[810] +
//             mat_A[986] * mat_B[842] +
//             mat_A[987] * mat_B[874] +
//             mat_A[988] * mat_B[906] +
//             mat_A[989] * mat_B[938] +
//             mat_A[990] * mat_B[970] +
//             mat_A[991] * mat_B[1002];
//  mat_C[971] <= 
//             mat_A[960] * mat_B[11] +
//             mat_A[961] * mat_B[43] +
//             mat_A[962] * mat_B[75] +
//             mat_A[963] * mat_B[107] +
//             mat_A[964] * mat_B[139] +
//             mat_A[965] * mat_B[171] +
//             mat_A[966] * mat_B[203] +
//             mat_A[967] * mat_B[235] +
//             mat_A[968] * mat_B[267] +
//             mat_A[969] * mat_B[299] +
//             mat_A[970] * mat_B[331] +
//             mat_A[971] * mat_B[363] +
//             mat_A[972] * mat_B[395] +
//             mat_A[973] * mat_B[427] +
//             mat_A[974] * mat_B[459] +
//             mat_A[975] * mat_B[491] +
//             mat_A[976] * mat_B[523] +
//             mat_A[977] * mat_B[555] +
//             mat_A[978] * mat_B[587] +
//             mat_A[979] * mat_B[619] +
//             mat_A[980] * mat_B[651] +
//             mat_A[981] * mat_B[683] +
//             mat_A[982] * mat_B[715] +
//             mat_A[983] * mat_B[747] +
//             mat_A[984] * mat_B[779] +
//             mat_A[985] * mat_B[811] +
//             mat_A[986] * mat_B[843] +
//             mat_A[987] * mat_B[875] +
//             mat_A[988] * mat_B[907] +
//             mat_A[989] * mat_B[939] +
//             mat_A[990] * mat_B[971] +
//             mat_A[991] * mat_B[1003];
//  mat_C[972] <= 
//             mat_A[960] * mat_B[12] +
//             mat_A[961] * mat_B[44] +
//             mat_A[962] * mat_B[76] +
//             mat_A[963] * mat_B[108] +
//             mat_A[964] * mat_B[140] +
//             mat_A[965] * mat_B[172] +
//             mat_A[966] * mat_B[204] +
//             mat_A[967] * mat_B[236] +
//             mat_A[968] * mat_B[268] +
//             mat_A[969] * mat_B[300] +
//             mat_A[970] * mat_B[332] +
//             mat_A[971] * mat_B[364] +
//             mat_A[972] * mat_B[396] +
//             mat_A[973] * mat_B[428] +
//             mat_A[974] * mat_B[460] +
//             mat_A[975] * mat_B[492] +
//             mat_A[976] * mat_B[524] +
//             mat_A[977] * mat_B[556] +
//             mat_A[978] * mat_B[588] +
//             mat_A[979] * mat_B[620] +
//             mat_A[980] * mat_B[652] +
//             mat_A[981] * mat_B[684] +
//             mat_A[982] * mat_B[716] +
//             mat_A[983] * mat_B[748] +
//             mat_A[984] * mat_B[780] +
//             mat_A[985] * mat_B[812] +
//             mat_A[986] * mat_B[844] +
//             mat_A[987] * mat_B[876] +
//             mat_A[988] * mat_B[908] +
//             mat_A[989] * mat_B[940] +
//             mat_A[990] * mat_B[972] +
//             mat_A[991] * mat_B[1004];
//  mat_C[973] <= 
//             mat_A[960] * mat_B[13] +
//             mat_A[961] * mat_B[45] +
//             mat_A[962] * mat_B[77] +
//             mat_A[963] * mat_B[109] +
//             mat_A[964] * mat_B[141] +
//             mat_A[965] * mat_B[173] +
//             mat_A[966] * mat_B[205] +
//             mat_A[967] * mat_B[237] +
//             mat_A[968] * mat_B[269] +
//             mat_A[969] * mat_B[301] +
//             mat_A[970] * mat_B[333] +
//             mat_A[971] * mat_B[365] +
//             mat_A[972] * mat_B[397] +
//             mat_A[973] * mat_B[429] +
//             mat_A[974] * mat_B[461] +
//             mat_A[975] * mat_B[493] +
//             mat_A[976] * mat_B[525] +
//             mat_A[977] * mat_B[557] +
//             mat_A[978] * mat_B[589] +
//             mat_A[979] * mat_B[621] +
//             mat_A[980] * mat_B[653] +
//             mat_A[981] * mat_B[685] +
//             mat_A[982] * mat_B[717] +
//             mat_A[983] * mat_B[749] +
//             mat_A[984] * mat_B[781] +
//             mat_A[985] * mat_B[813] +
//             mat_A[986] * mat_B[845] +
//             mat_A[987] * mat_B[877] +
//             mat_A[988] * mat_B[909] +
//             mat_A[989] * mat_B[941] +
//             mat_A[990] * mat_B[973] +
//             mat_A[991] * mat_B[1005];
//  mat_C[974] <= 
//             mat_A[960] * mat_B[14] +
//             mat_A[961] * mat_B[46] +
//             mat_A[962] * mat_B[78] +
//             mat_A[963] * mat_B[110] +
//             mat_A[964] * mat_B[142] +
//             mat_A[965] * mat_B[174] +
//             mat_A[966] * mat_B[206] +
//             mat_A[967] * mat_B[238] +
//             mat_A[968] * mat_B[270] +
//             mat_A[969] * mat_B[302] +
//             mat_A[970] * mat_B[334] +
//             mat_A[971] * mat_B[366] +
//             mat_A[972] * mat_B[398] +
//             mat_A[973] * mat_B[430] +
//             mat_A[974] * mat_B[462] +
//             mat_A[975] * mat_B[494] +
//             mat_A[976] * mat_B[526] +
//             mat_A[977] * mat_B[558] +
//             mat_A[978] * mat_B[590] +
//             mat_A[979] * mat_B[622] +
//             mat_A[980] * mat_B[654] +
//             mat_A[981] * mat_B[686] +
//             mat_A[982] * mat_B[718] +
//             mat_A[983] * mat_B[750] +
//             mat_A[984] * mat_B[782] +
//             mat_A[985] * mat_B[814] +
//             mat_A[986] * mat_B[846] +
//             mat_A[987] * mat_B[878] +
//             mat_A[988] * mat_B[910] +
//             mat_A[989] * mat_B[942] +
//             mat_A[990] * mat_B[974] +
//             mat_A[991] * mat_B[1006];
//  mat_C[975] <= 
//             mat_A[960] * mat_B[15] +
//             mat_A[961] * mat_B[47] +
//             mat_A[962] * mat_B[79] +
//             mat_A[963] * mat_B[111] +
//             mat_A[964] * mat_B[143] +
//             mat_A[965] * mat_B[175] +
//             mat_A[966] * mat_B[207] +
//             mat_A[967] * mat_B[239] +
//             mat_A[968] * mat_B[271] +
//             mat_A[969] * mat_B[303] +
//             mat_A[970] * mat_B[335] +
//             mat_A[971] * mat_B[367] +
//             mat_A[972] * mat_B[399] +
//             mat_A[973] * mat_B[431] +
//             mat_A[974] * mat_B[463] +
//             mat_A[975] * mat_B[495] +
//             mat_A[976] * mat_B[527] +
//             mat_A[977] * mat_B[559] +
//             mat_A[978] * mat_B[591] +
//             mat_A[979] * mat_B[623] +
//             mat_A[980] * mat_B[655] +
//             mat_A[981] * mat_B[687] +
//             mat_A[982] * mat_B[719] +
//             mat_A[983] * mat_B[751] +
//             mat_A[984] * mat_B[783] +
//             mat_A[985] * mat_B[815] +
//             mat_A[986] * mat_B[847] +
//             mat_A[987] * mat_B[879] +
//             mat_A[988] * mat_B[911] +
//             mat_A[989] * mat_B[943] +
//             mat_A[990] * mat_B[975] +
//             mat_A[991] * mat_B[1007];
//  mat_C[976] <= 
//             mat_A[960] * mat_B[16] +
//             mat_A[961] * mat_B[48] +
//             mat_A[962] * mat_B[80] +
//             mat_A[963] * mat_B[112] +
//             mat_A[964] * mat_B[144] +
//             mat_A[965] * mat_B[176] +
//             mat_A[966] * mat_B[208] +
//             mat_A[967] * mat_B[240] +
//             mat_A[968] * mat_B[272] +
//             mat_A[969] * mat_B[304] +
//             mat_A[970] * mat_B[336] +
//             mat_A[971] * mat_B[368] +
//             mat_A[972] * mat_B[400] +
//             mat_A[973] * mat_B[432] +
//             mat_A[974] * mat_B[464] +
//             mat_A[975] * mat_B[496] +
//             mat_A[976] * mat_B[528] +
//             mat_A[977] * mat_B[560] +
//             mat_A[978] * mat_B[592] +
//             mat_A[979] * mat_B[624] +
//             mat_A[980] * mat_B[656] +
//             mat_A[981] * mat_B[688] +
//             mat_A[982] * mat_B[720] +
//             mat_A[983] * mat_B[752] +
//             mat_A[984] * mat_B[784] +
//             mat_A[985] * mat_B[816] +
//             mat_A[986] * mat_B[848] +
//             mat_A[987] * mat_B[880] +
//             mat_A[988] * mat_B[912] +
//             mat_A[989] * mat_B[944] +
//             mat_A[990] * mat_B[976] +
//             mat_A[991] * mat_B[1008];
//  mat_C[977] <= 
//             mat_A[960] * mat_B[17] +
//             mat_A[961] * mat_B[49] +
//             mat_A[962] * mat_B[81] +
//             mat_A[963] * mat_B[113] +
//             mat_A[964] * mat_B[145] +
//             mat_A[965] * mat_B[177] +
//             mat_A[966] * mat_B[209] +
//             mat_A[967] * mat_B[241] +
//             mat_A[968] * mat_B[273] +
//             mat_A[969] * mat_B[305] +
//             mat_A[970] * mat_B[337] +
//             mat_A[971] * mat_B[369] +
//             mat_A[972] * mat_B[401] +
//             mat_A[973] * mat_B[433] +
//             mat_A[974] * mat_B[465] +
//             mat_A[975] * mat_B[497] +
//             mat_A[976] * mat_B[529] +
//             mat_A[977] * mat_B[561] +
//             mat_A[978] * mat_B[593] +
//             mat_A[979] * mat_B[625] +
//             mat_A[980] * mat_B[657] +
//             mat_A[981] * mat_B[689] +
//             mat_A[982] * mat_B[721] +
//             mat_A[983] * mat_B[753] +
//             mat_A[984] * mat_B[785] +
//             mat_A[985] * mat_B[817] +
//             mat_A[986] * mat_B[849] +
//             mat_A[987] * mat_B[881] +
//             mat_A[988] * mat_B[913] +
//             mat_A[989] * mat_B[945] +
//             mat_A[990] * mat_B[977] +
//             mat_A[991] * mat_B[1009];
//  mat_C[978] <= 
//             mat_A[960] * mat_B[18] +
//             mat_A[961] * mat_B[50] +
//             mat_A[962] * mat_B[82] +
//             mat_A[963] * mat_B[114] +
//             mat_A[964] * mat_B[146] +
//             mat_A[965] * mat_B[178] +
//             mat_A[966] * mat_B[210] +
//             mat_A[967] * mat_B[242] +
//             mat_A[968] * mat_B[274] +
//             mat_A[969] * mat_B[306] +
//             mat_A[970] * mat_B[338] +
//             mat_A[971] * mat_B[370] +
//             mat_A[972] * mat_B[402] +
//             mat_A[973] * mat_B[434] +
//             mat_A[974] * mat_B[466] +
//             mat_A[975] * mat_B[498] +
//             mat_A[976] * mat_B[530] +
//             mat_A[977] * mat_B[562] +
//             mat_A[978] * mat_B[594] +
//             mat_A[979] * mat_B[626] +
//             mat_A[980] * mat_B[658] +
//             mat_A[981] * mat_B[690] +
//             mat_A[982] * mat_B[722] +
//             mat_A[983] * mat_B[754] +
//             mat_A[984] * mat_B[786] +
//             mat_A[985] * mat_B[818] +
//             mat_A[986] * mat_B[850] +
//             mat_A[987] * mat_B[882] +
//             mat_A[988] * mat_B[914] +
//             mat_A[989] * mat_B[946] +
//             mat_A[990] * mat_B[978] +
//             mat_A[991] * mat_B[1010];
//  mat_C[979] <= 
//             mat_A[960] * mat_B[19] +
//             mat_A[961] * mat_B[51] +
//             mat_A[962] * mat_B[83] +
//             mat_A[963] * mat_B[115] +
//             mat_A[964] * mat_B[147] +
//             mat_A[965] * mat_B[179] +
//             mat_A[966] * mat_B[211] +
//             mat_A[967] * mat_B[243] +
//             mat_A[968] * mat_B[275] +
//             mat_A[969] * mat_B[307] +
//             mat_A[970] * mat_B[339] +
//             mat_A[971] * mat_B[371] +
//             mat_A[972] * mat_B[403] +
//             mat_A[973] * mat_B[435] +
//             mat_A[974] * mat_B[467] +
//             mat_A[975] * mat_B[499] +
//             mat_A[976] * mat_B[531] +
//             mat_A[977] * mat_B[563] +
//             mat_A[978] * mat_B[595] +
//             mat_A[979] * mat_B[627] +
//             mat_A[980] * mat_B[659] +
//             mat_A[981] * mat_B[691] +
//             mat_A[982] * mat_B[723] +
//             mat_A[983] * mat_B[755] +
//             mat_A[984] * mat_B[787] +
//             mat_A[985] * mat_B[819] +
//             mat_A[986] * mat_B[851] +
//             mat_A[987] * mat_B[883] +
//             mat_A[988] * mat_B[915] +
//             mat_A[989] * mat_B[947] +
//             mat_A[990] * mat_B[979] +
//             mat_A[991] * mat_B[1011];
//  mat_C[980] <= 
//             mat_A[960] * mat_B[20] +
//             mat_A[961] * mat_B[52] +
//             mat_A[962] * mat_B[84] +
//             mat_A[963] * mat_B[116] +
//             mat_A[964] * mat_B[148] +
//             mat_A[965] * mat_B[180] +
//             mat_A[966] * mat_B[212] +
//             mat_A[967] * mat_B[244] +
//             mat_A[968] * mat_B[276] +
//             mat_A[969] * mat_B[308] +
//             mat_A[970] * mat_B[340] +
//             mat_A[971] * mat_B[372] +
//             mat_A[972] * mat_B[404] +
//             mat_A[973] * mat_B[436] +
//             mat_A[974] * mat_B[468] +
//             mat_A[975] * mat_B[500] +
//             mat_A[976] * mat_B[532] +
//             mat_A[977] * mat_B[564] +
//             mat_A[978] * mat_B[596] +
//             mat_A[979] * mat_B[628] +
//             mat_A[980] * mat_B[660] +
//             mat_A[981] * mat_B[692] +
//             mat_A[982] * mat_B[724] +
//             mat_A[983] * mat_B[756] +
//             mat_A[984] * mat_B[788] +
//             mat_A[985] * mat_B[820] +
//             mat_A[986] * mat_B[852] +
//             mat_A[987] * mat_B[884] +
//             mat_A[988] * mat_B[916] +
//             mat_A[989] * mat_B[948] +
//             mat_A[990] * mat_B[980] +
//             mat_A[991] * mat_B[1012];
//  mat_C[981] <= 
//             mat_A[960] * mat_B[21] +
//             mat_A[961] * mat_B[53] +
//             mat_A[962] * mat_B[85] +
//             mat_A[963] * mat_B[117] +
//             mat_A[964] * mat_B[149] +
//             mat_A[965] * mat_B[181] +
//             mat_A[966] * mat_B[213] +
//             mat_A[967] * mat_B[245] +
//             mat_A[968] * mat_B[277] +
//             mat_A[969] * mat_B[309] +
//             mat_A[970] * mat_B[341] +
//             mat_A[971] * mat_B[373] +
//             mat_A[972] * mat_B[405] +
//             mat_A[973] * mat_B[437] +
//             mat_A[974] * mat_B[469] +
//             mat_A[975] * mat_B[501] +
//             mat_A[976] * mat_B[533] +
//             mat_A[977] * mat_B[565] +
//             mat_A[978] * mat_B[597] +
//             mat_A[979] * mat_B[629] +
//             mat_A[980] * mat_B[661] +
//             mat_A[981] * mat_B[693] +
//             mat_A[982] * mat_B[725] +
//             mat_A[983] * mat_B[757] +
//             mat_A[984] * mat_B[789] +
//             mat_A[985] * mat_B[821] +
//             mat_A[986] * mat_B[853] +
//             mat_A[987] * mat_B[885] +
//             mat_A[988] * mat_B[917] +
//             mat_A[989] * mat_B[949] +
//             mat_A[990] * mat_B[981] +
//             mat_A[991] * mat_B[1013];
//  mat_C[982] <= 
//             mat_A[960] * mat_B[22] +
//             mat_A[961] * mat_B[54] +
//             mat_A[962] * mat_B[86] +
//             mat_A[963] * mat_B[118] +
//             mat_A[964] * mat_B[150] +
//             mat_A[965] * mat_B[182] +
//             mat_A[966] * mat_B[214] +
//             mat_A[967] * mat_B[246] +
//             mat_A[968] * mat_B[278] +
//             mat_A[969] * mat_B[310] +
//             mat_A[970] * mat_B[342] +
//             mat_A[971] * mat_B[374] +
//             mat_A[972] * mat_B[406] +
//             mat_A[973] * mat_B[438] +
//             mat_A[974] * mat_B[470] +
//             mat_A[975] * mat_B[502] +
//             mat_A[976] * mat_B[534] +
//             mat_A[977] * mat_B[566] +
//             mat_A[978] * mat_B[598] +
//             mat_A[979] * mat_B[630] +
//             mat_A[980] * mat_B[662] +
//             mat_A[981] * mat_B[694] +
//             mat_A[982] * mat_B[726] +
//             mat_A[983] * mat_B[758] +
//             mat_A[984] * mat_B[790] +
//             mat_A[985] * mat_B[822] +
//             mat_A[986] * mat_B[854] +
//             mat_A[987] * mat_B[886] +
//             mat_A[988] * mat_B[918] +
//             mat_A[989] * mat_B[950] +
//             mat_A[990] * mat_B[982] +
//             mat_A[991] * mat_B[1014];
//  mat_C[983] <= 
//             mat_A[960] * mat_B[23] +
//             mat_A[961] * mat_B[55] +
//             mat_A[962] * mat_B[87] +
//             mat_A[963] * mat_B[119] +
//             mat_A[964] * mat_B[151] +
//             mat_A[965] * mat_B[183] +
//             mat_A[966] * mat_B[215] +
//             mat_A[967] * mat_B[247] +
//             mat_A[968] * mat_B[279] +
//             mat_A[969] * mat_B[311] +
//             mat_A[970] * mat_B[343] +
//             mat_A[971] * mat_B[375] +
//             mat_A[972] * mat_B[407] +
//             mat_A[973] * mat_B[439] +
//             mat_A[974] * mat_B[471] +
//             mat_A[975] * mat_B[503] +
//             mat_A[976] * mat_B[535] +
//             mat_A[977] * mat_B[567] +
//             mat_A[978] * mat_B[599] +
//             mat_A[979] * mat_B[631] +
//             mat_A[980] * mat_B[663] +
//             mat_A[981] * mat_B[695] +
//             mat_A[982] * mat_B[727] +
//             mat_A[983] * mat_B[759] +
//             mat_A[984] * mat_B[791] +
//             mat_A[985] * mat_B[823] +
//             mat_A[986] * mat_B[855] +
//             mat_A[987] * mat_B[887] +
//             mat_A[988] * mat_B[919] +
//             mat_A[989] * mat_B[951] +
//             mat_A[990] * mat_B[983] +
//             mat_A[991] * mat_B[1015];
//  mat_C[984] <= 
//             mat_A[960] * mat_B[24] +
//             mat_A[961] * mat_B[56] +
//             mat_A[962] * mat_B[88] +
//             mat_A[963] * mat_B[120] +
//             mat_A[964] * mat_B[152] +
//             mat_A[965] * mat_B[184] +
//             mat_A[966] * mat_B[216] +
//             mat_A[967] * mat_B[248] +
//             mat_A[968] * mat_B[280] +
//             mat_A[969] * mat_B[312] +
//             mat_A[970] * mat_B[344] +
//             mat_A[971] * mat_B[376] +
//             mat_A[972] * mat_B[408] +
//             mat_A[973] * mat_B[440] +
//             mat_A[974] * mat_B[472] +
//             mat_A[975] * mat_B[504] +
//             mat_A[976] * mat_B[536] +
//             mat_A[977] * mat_B[568] +
//             mat_A[978] * mat_B[600] +
//             mat_A[979] * mat_B[632] +
//             mat_A[980] * mat_B[664] +
//             mat_A[981] * mat_B[696] +
//             mat_A[982] * mat_B[728] +
//             mat_A[983] * mat_B[760] +
//             mat_A[984] * mat_B[792] +
//             mat_A[985] * mat_B[824] +
//             mat_A[986] * mat_B[856] +
//             mat_A[987] * mat_B[888] +
//             mat_A[988] * mat_B[920] +
//             mat_A[989] * mat_B[952] +
//             mat_A[990] * mat_B[984] +
//             mat_A[991] * mat_B[1016];
//  mat_C[985] <= 
//             mat_A[960] * mat_B[25] +
//             mat_A[961] * mat_B[57] +
//             mat_A[962] * mat_B[89] +
//             mat_A[963] * mat_B[121] +
//             mat_A[964] * mat_B[153] +
//             mat_A[965] * mat_B[185] +
//             mat_A[966] * mat_B[217] +
//             mat_A[967] * mat_B[249] +
//             mat_A[968] * mat_B[281] +
//             mat_A[969] * mat_B[313] +
//             mat_A[970] * mat_B[345] +
//             mat_A[971] * mat_B[377] +
//             mat_A[972] * mat_B[409] +
//             mat_A[973] * mat_B[441] +
//             mat_A[974] * mat_B[473] +
//             mat_A[975] * mat_B[505] +
//             mat_A[976] * mat_B[537] +
//             mat_A[977] * mat_B[569] +
//             mat_A[978] * mat_B[601] +
//             mat_A[979] * mat_B[633] +
//             mat_A[980] * mat_B[665] +
//             mat_A[981] * mat_B[697] +
//             mat_A[982] * mat_B[729] +
//             mat_A[983] * mat_B[761] +
//             mat_A[984] * mat_B[793] +
//             mat_A[985] * mat_B[825] +
//             mat_A[986] * mat_B[857] +
//             mat_A[987] * mat_B[889] +
//             mat_A[988] * mat_B[921] +
//             mat_A[989] * mat_B[953] +
//             mat_A[990] * mat_B[985] +
//             mat_A[991] * mat_B[1017];
//  mat_C[986] <= 
//             mat_A[960] * mat_B[26] +
//             mat_A[961] * mat_B[58] +
//             mat_A[962] * mat_B[90] +
//             mat_A[963] * mat_B[122] +
//             mat_A[964] * mat_B[154] +
//             mat_A[965] * mat_B[186] +
//             mat_A[966] * mat_B[218] +
//             mat_A[967] * mat_B[250] +
//             mat_A[968] * mat_B[282] +
//             mat_A[969] * mat_B[314] +
//             mat_A[970] * mat_B[346] +
//             mat_A[971] * mat_B[378] +
//             mat_A[972] * mat_B[410] +
//             mat_A[973] * mat_B[442] +
//             mat_A[974] * mat_B[474] +
//             mat_A[975] * mat_B[506] +
//             mat_A[976] * mat_B[538] +
//             mat_A[977] * mat_B[570] +
//             mat_A[978] * mat_B[602] +
//             mat_A[979] * mat_B[634] +
//             mat_A[980] * mat_B[666] +
//             mat_A[981] * mat_B[698] +
//             mat_A[982] * mat_B[730] +
//             mat_A[983] * mat_B[762] +
//             mat_A[984] * mat_B[794] +
//             mat_A[985] * mat_B[826] +
//             mat_A[986] * mat_B[858] +
//             mat_A[987] * mat_B[890] +
//             mat_A[988] * mat_B[922] +
//             mat_A[989] * mat_B[954] +
//             mat_A[990] * mat_B[986] +
//             mat_A[991] * mat_B[1018];
//  mat_C[987] <= 
//             mat_A[960] * mat_B[27] +
//             mat_A[961] * mat_B[59] +
//             mat_A[962] * mat_B[91] +
//             mat_A[963] * mat_B[123] +
//             mat_A[964] * mat_B[155] +
//             mat_A[965] * mat_B[187] +
//             mat_A[966] * mat_B[219] +
//             mat_A[967] * mat_B[251] +
//             mat_A[968] * mat_B[283] +
//             mat_A[969] * mat_B[315] +
//             mat_A[970] * mat_B[347] +
//             mat_A[971] * mat_B[379] +
//             mat_A[972] * mat_B[411] +
//             mat_A[973] * mat_B[443] +
//             mat_A[974] * mat_B[475] +
//             mat_A[975] * mat_B[507] +
//             mat_A[976] * mat_B[539] +
//             mat_A[977] * mat_B[571] +
//             mat_A[978] * mat_B[603] +
//             mat_A[979] * mat_B[635] +
//             mat_A[980] * mat_B[667] +
//             mat_A[981] * mat_B[699] +
//             mat_A[982] * mat_B[731] +
//             mat_A[983] * mat_B[763] +
//             mat_A[984] * mat_B[795] +
//             mat_A[985] * mat_B[827] +
//             mat_A[986] * mat_B[859] +
//             mat_A[987] * mat_B[891] +
//             mat_A[988] * mat_B[923] +
//             mat_A[989] * mat_B[955] +
//             mat_A[990] * mat_B[987] +
//             mat_A[991] * mat_B[1019];
//  mat_C[988] <= 
//             mat_A[960] * mat_B[28] +
//             mat_A[961] * mat_B[60] +
//             mat_A[962] * mat_B[92] +
//             mat_A[963] * mat_B[124] +
//             mat_A[964] * mat_B[156] +
//             mat_A[965] * mat_B[188] +
//             mat_A[966] * mat_B[220] +
//             mat_A[967] * mat_B[252] +
//             mat_A[968] * mat_B[284] +
//             mat_A[969] * mat_B[316] +
//             mat_A[970] * mat_B[348] +
//             mat_A[971] * mat_B[380] +
//             mat_A[972] * mat_B[412] +
//             mat_A[973] * mat_B[444] +
//             mat_A[974] * mat_B[476] +
//             mat_A[975] * mat_B[508] +
//             mat_A[976] * mat_B[540] +
//             mat_A[977] * mat_B[572] +
//             mat_A[978] * mat_B[604] +
//             mat_A[979] * mat_B[636] +
//             mat_A[980] * mat_B[668] +
//             mat_A[981] * mat_B[700] +
//             mat_A[982] * mat_B[732] +
//             mat_A[983] * mat_B[764] +
//             mat_A[984] * mat_B[796] +
//             mat_A[985] * mat_B[828] +
//             mat_A[986] * mat_B[860] +
//             mat_A[987] * mat_B[892] +
//             mat_A[988] * mat_B[924] +
//             mat_A[989] * mat_B[956] +
//             mat_A[990] * mat_B[988] +
//             mat_A[991] * mat_B[1020];
//  mat_C[989] <= 
//             mat_A[960] * mat_B[29] +
//             mat_A[961] * mat_B[61] +
//             mat_A[962] * mat_B[93] +
//             mat_A[963] * mat_B[125] +
//             mat_A[964] * mat_B[157] +
//             mat_A[965] * mat_B[189] +
//             mat_A[966] * mat_B[221] +
//             mat_A[967] * mat_B[253] +
//             mat_A[968] * mat_B[285] +
//             mat_A[969] * mat_B[317] +
//             mat_A[970] * mat_B[349] +
//             mat_A[971] * mat_B[381] +
//             mat_A[972] * mat_B[413] +
//             mat_A[973] * mat_B[445] +
//             mat_A[974] * mat_B[477] +
//             mat_A[975] * mat_B[509] +
//             mat_A[976] * mat_B[541] +
//             mat_A[977] * mat_B[573] +
//             mat_A[978] * mat_B[605] +
//             mat_A[979] * mat_B[637] +
//             mat_A[980] * mat_B[669] +
//             mat_A[981] * mat_B[701] +
//             mat_A[982] * mat_B[733] +
//             mat_A[983] * mat_B[765] +
//             mat_A[984] * mat_B[797] +
//             mat_A[985] * mat_B[829] +
//             mat_A[986] * mat_B[861] +
//             mat_A[987] * mat_B[893] +
//             mat_A[988] * mat_B[925] +
//             mat_A[989] * mat_B[957] +
//             mat_A[990] * mat_B[989] +
//             mat_A[991] * mat_B[1021];
//  mat_C[990] <= 
//             mat_A[960] * mat_B[30] +
//             mat_A[961] * mat_B[62] +
//             mat_A[962] * mat_B[94] +
//             mat_A[963] * mat_B[126] +
//             mat_A[964] * mat_B[158] +
//             mat_A[965] * mat_B[190] +
//             mat_A[966] * mat_B[222] +
//             mat_A[967] * mat_B[254] +
//             mat_A[968] * mat_B[286] +
//             mat_A[969] * mat_B[318] +
//             mat_A[970] * mat_B[350] +
//             mat_A[971] * mat_B[382] +
//             mat_A[972] * mat_B[414] +
//             mat_A[973] * mat_B[446] +
//             mat_A[974] * mat_B[478] +
//             mat_A[975] * mat_B[510] +
//             mat_A[976] * mat_B[542] +
//             mat_A[977] * mat_B[574] +
//             mat_A[978] * mat_B[606] +
//             mat_A[979] * mat_B[638] +
//             mat_A[980] * mat_B[670] +
//             mat_A[981] * mat_B[702] +
//             mat_A[982] * mat_B[734] +
//             mat_A[983] * mat_B[766] +
//             mat_A[984] * mat_B[798] +
//             mat_A[985] * mat_B[830] +
//             mat_A[986] * mat_B[862] +
//             mat_A[987] * mat_B[894] +
//             mat_A[988] * mat_B[926] +
//             mat_A[989] * mat_B[958] +
//             mat_A[990] * mat_B[990] +
//             mat_A[991] * mat_B[1022];
//  mat_C[991] <= 
//             mat_A[960] * mat_B[31] +
//             mat_A[961] * mat_B[63] +
//             mat_A[962] * mat_B[95] +
//             mat_A[963] * mat_B[127] +
//             mat_A[964] * mat_B[159] +
//             mat_A[965] * mat_B[191] +
//             mat_A[966] * mat_B[223] +
//             mat_A[967] * mat_B[255] +
//             mat_A[968] * mat_B[287] +
//             mat_A[969] * mat_B[319] +
//             mat_A[970] * mat_B[351] +
//             mat_A[971] * mat_B[383] +
//             mat_A[972] * mat_B[415] +
//             mat_A[973] * mat_B[447] +
//             mat_A[974] * mat_B[479] +
//             mat_A[975] * mat_B[511] +
//             mat_A[976] * mat_B[543] +
//             mat_A[977] * mat_B[575] +
//             mat_A[978] * mat_B[607] +
//             mat_A[979] * mat_B[639] +
//             mat_A[980] * mat_B[671] +
//             mat_A[981] * mat_B[703] +
//             mat_A[982] * mat_B[735] +
//             mat_A[983] * mat_B[767] +
//             mat_A[984] * mat_B[799] +
//             mat_A[985] * mat_B[831] +
//             mat_A[986] * mat_B[863] +
//             mat_A[987] * mat_B[895] +
//             mat_A[988] * mat_B[927] +
//             mat_A[989] * mat_B[959] +
//             mat_A[990] * mat_B[991] +
//             mat_A[991] * mat_B[1023];
//  mat_C[992] <= 
//             mat_A[992] * mat_B[0] +
//             mat_A[993] * mat_B[32] +
//             mat_A[994] * mat_B[64] +
//             mat_A[995] * mat_B[96] +
//             mat_A[996] * mat_B[128] +
//             mat_A[997] * mat_B[160] +
//             mat_A[998] * mat_B[192] +
//             mat_A[999] * mat_B[224] +
//             mat_A[1000] * mat_B[256] +
//             mat_A[1001] * mat_B[288] +
//             mat_A[1002] * mat_B[320] +
//             mat_A[1003] * mat_B[352] +
//             mat_A[1004] * mat_B[384] +
//             mat_A[1005] * mat_B[416] +
//             mat_A[1006] * mat_B[448] +
//             mat_A[1007] * mat_B[480] +
//             mat_A[1008] * mat_B[512] +
//             mat_A[1009] * mat_B[544] +
//             mat_A[1010] * mat_B[576] +
//             mat_A[1011] * mat_B[608] +
//             mat_A[1012] * mat_B[640] +
//             mat_A[1013] * mat_B[672] +
//             mat_A[1014] * mat_B[704] +
//             mat_A[1015] * mat_B[736] +
//             mat_A[1016] * mat_B[768] +
//             mat_A[1017] * mat_B[800] +
//             mat_A[1018] * mat_B[832] +
//             mat_A[1019] * mat_B[864] +
//             mat_A[1020] * mat_B[896] +
//             mat_A[1021] * mat_B[928] +
//             mat_A[1022] * mat_B[960] +
//             mat_A[1023] * mat_B[992];
//  mat_C[993] <= 
//             mat_A[992] * mat_B[1] +
//             mat_A[993] * mat_B[33] +
//             mat_A[994] * mat_B[65] +
//             mat_A[995] * mat_B[97] +
//             mat_A[996] * mat_B[129] +
//             mat_A[997] * mat_B[161] +
//             mat_A[998] * mat_B[193] +
//             mat_A[999] * mat_B[225] +
//             mat_A[1000] * mat_B[257] +
//             mat_A[1001] * mat_B[289] +
//             mat_A[1002] * mat_B[321] +
//             mat_A[1003] * mat_B[353] +
//             mat_A[1004] * mat_B[385] +
//             mat_A[1005] * mat_B[417] +
//             mat_A[1006] * mat_B[449] +
//             mat_A[1007] * mat_B[481] +
//             mat_A[1008] * mat_B[513] +
//             mat_A[1009] * mat_B[545] +
//             mat_A[1010] * mat_B[577] +
//             mat_A[1011] * mat_B[609] +
//             mat_A[1012] * mat_B[641] +
//             mat_A[1013] * mat_B[673] +
//             mat_A[1014] * mat_B[705] +
//             mat_A[1015] * mat_B[737] +
//             mat_A[1016] * mat_B[769] +
//             mat_A[1017] * mat_B[801] +
//             mat_A[1018] * mat_B[833] +
//             mat_A[1019] * mat_B[865] +
//             mat_A[1020] * mat_B[897] +
//             mat_A[1021] * mat_B[929] +
//             mat_A[1022] * mat_B[961] +
//             mat_A[1023] * mat_B[993];
//  mat_C[994] <= 
//             mat_A[992] * mat_B[2] +
//             mat_A[993] * mat_B[34] +
//             mat_A[994] * mat_B[66] +
//             mat_A[995] * mat_B[98] +
//             mat_A[996] * mat_B[130] +
//             mat_A[997] * mat_B[162] +
//             mat_A[998] * mat_B[194] +
//             mat_A[999] * mat_B[226] +
//             mat_A[1000] * mat_B[258] +
//             mat_A[1001] * mat_B[290] +
//             mat_A[1002] * mat_B[322] +
//             mat_A[1003] * mat_B[354] +
//             mat_A[1004] * mat_B[386] +
//             mat_A[1005] * mat_B[418] +
//             mat_A[1006] * mat_B[450] +
//             mat_A[1007] * mat_B[482] +
//             mat_A[1008] * mat_B[514] +
//             mat_A[1009] * mat_B[546] +
//             mat_A[1010] * mat_B[578] +
//             mat_A[1011] * mat_B[610] +
//             mat_A[1012] * mat_B[642] +
//             mat_A[1013] * mat_B[674] +
//             mat_A[1014] * mat_B[706] +
//             mat_A[1015] * mat_B[738] +
//             mat_A[1016] * mat_B[770] +
//             mat_A[1017] * mat_B[802] +
//             mat_A[1018] * mat_B[834] +
//             mat_A[1019] * mat_B[866] +
//             mat_A[1020] * mat_B[898] +
//             mat_A[1021] * mat_B[930] +
//             mat_A[1022] * mat_B[962] +
//             mat_A[1023] * mat_B[994];
//  mat_C[995] <= 
//             mat_A[992] * mat_B[3] +
//             mat_A[993] * mat_B[35] +
//             mat_A[994] * mat_B[67] +
//             mat_A[995] * mat_B[99] +
//             mat_A[996] * mat_B[131] +
//             mat_A[997] * mat_B[163] +
//             mat_A[998] * mat_B[195] +
//             mat_A[999] * mat_B[227] +
//             mat_A[1000] * mat_B[259] +
//             mat_A[1001] * mat_B[291] +
//             mat_A[1002] * mat_B[323] +
//             mat_A[1003] * mat_B[355] +
//             mat_A[1004] * mat_B[387] +
//             mat_A[1005] * mat_B[419] +
//             mat_A[1006] * mat_B[451] +
//             mat_A[1007] * mat_B[483] +
//             mat_A[1008] * mat_B[515] +
//             mat_A[1009] * mat_B[547] +
//             mat_A[1010] * mat_B[579] +
//             mat_A[1011] * mat_B[611] +
//             mat_A[1012] * mat_B[643] +
//             mat_A[1013] * mat_B[675] +
//             mat_A[1014] * mat_B[707] +
//             mat_A[1015] * mat_B[739] +
//             mat_A[1016] * mat_B[771] +
//             mat_A[1017] * mat_B[803] +
//             mat_A[1018] * mat_B[835] +
//             mat_A[1019] * mat_B[867] +
//             mat_A[1020] * mat_B[899] +
//             mat_A[1021] * mat_B[931] +
//             mat_A[1022] * mat_B[963] +
//             mat_A[1023] * mat_B[995];
//  mat_C[996] <= 
//             mat_A[992] * mat_B[4] +
//             mat_A[993] * mat_B[36] +
//             mat_A[994] * mat_B[68] +
//             mat_A[995] * mat_B[100] +
//             mat_A[996] * mat_B[132] +
//             mat_A[997] * mat_B[164] +
//             mat_A[998] * mat_B[196] +
//             mat_A[999] * mat_B[228] +
//             mat_A[1000] * mat_B[260] +
//             mat_A[1001] * mat_B[292] +
//             mat_A[1002] * mat_B[324] +
//             mat_A[1003] * mat_B[356] +
//             mat_A[1004] * mat_B[388] +
//             mat_A[1005] * mat_B[420] +
//             mat_A[1006] * mat_B[452] +
//             mat_A[1007] * mat_B[484] +
//             mat_A[1008] * mat_B[516] +
//             mat_A[1009] * mat_B[548] +
//             mat_A[1010] * mat_B[580] +
//             mat_A[1011] * mat_B[612] +
//             mat_A[1012] * mat_B[644] +
//             mat_A[1013] * mat_B[676] +
//             mat_A[1014] * mat_B[708] +
//             mat_A[1015] * mat_B[740] +
//             mat_A[1016] * mat_B[772] +
//             mat_A[1017] * mat_B[804] +
//             mat_A[1018] * mat_B[836] +
//             mat_A[1019] * mat_B[868] +
//             mat_A[1020] * mat_B[900] +
//             mat_A[1021] * mat_B[932] +
//             mat_A[1022] * mat_B[964] +
//             mat_A[1023] * mat_B[996];
//  mat_C[997] <= 
//             mat_A[992] * mat_B[5] +
//             mat_A[993] * mat_B[37] +
//             mat_A[994] * mat_B[69] +
//             mat_A[995] * mat_B[101] +
//             mat_A[996] * mat_B[133] +
//             mat_A[997] * mat_B[165] +
//             mat_A[998] * mat_B[197] +
//             mat_A[999] * mat_B[229] +
//             mat_A[1000] * mat_B[261] +
//             mat_A[1001] * mat_B[293] +
//             mat_A[1002] * mat_B[325] +
//             mat_A[1003] * mat_B[357] +
//             mat_A[1004] * mat_B[389] +
//             mat_A[1005] * mat_B[421] +
//             mat_A[1006] * mat_B[453] +
//             mat_A[1007] * mat_B[485] +
//             mat_A[1008] * mat_B[517] +
//             mat_A[1009] * mat_B[549] +
//             mat_A[1010] * mat_B[581] +
//             mat_A[1011] * mat_B[613] +
//             mat_A[1012] * mat_B[645] +
//             mat_A[1013] * mat_B[677] +
//             mat_A[1014] * mat_B[709] +
//             mat_A[1015] * mat_B[741] +
//             mat_A[1016] * mat_B[773] +
//             mat_A[1017] * mat_B[805] +
//             mat_A[1018] * mat_B[837] +
//             mat_A[1019] * mat_B[869] +
//             mat_A[1020] * mat_B[901] +
//             mat_A[1021] * mat_B[933] +
//             mat_A[1022] * mat_B[965] +
//             mat_A[1023] * mat_B[997];
//  mat_C[998] <= 
//             mat_A[992] * mat_B[6] +
//             mat_A[993] * mat_B[38] +
//             mat_A[994] * mat_B[70] +
//             mat_A[995] * mat_B[102] +
//             mat_A[996] * mat_B[134] +
//             mat_A[997] * mat_B[166] +
//             mat_A[998] * mat_B[198] +
//             mat_A[999] * mat_B[230] +
//             mat_A[1000] * mat_B[262] +
//             mat_A[1001] * mat_B[294] +
//             mat_A[1002] * mat_B[326] +
//             mat_A[1003] * mat_B[358] +
//             mat_A[1004] * mat_B[390] +
//             mat_A[1005] * mat_B[422] +
//             mat_A[1006] * mat_B[454] +
//             mat_A[1007] * mat_B[486] +
//             mat_A[1008] * mat_B[518] +
//             mat_A[1009] * mat_B[550] +
//             mat_A[1010] * mat_B[582] +
//             mat_A[1011] * mat_B[614] +
//             mat_A[1012] * mat_B[646] +
//             mat_A[1013] * mat_B[678] +
//             mat_A[1014] * mat_B[710] +
//             mat_A[1015] * mat_B[742] +
//             mat_A[1016] * mat_B[774] +
//             mat_A[1017] * mat_B[806] +
//             mat_A[1018] * mat_B[838] +
//             mat_A[1019] * mat_B[870] +
//             mat_A[1020] * mat_B[902] +
//             mat_A[1021] * mat_B[934] +
//             mat_A[1022] * mat_B[966] +
//             mat_A[1023] * mat_B[998];
//  mat_C[999] <= 
//             mat_A[992] * mat_B[7] +
//             mat_A[993] * mat_B[39] +
//             mat_A[994] * mat_B[71] +
//             mat_A[995] * mat_B[103] +
//             mat_A[996] * mat_B[135] +
//             mat_A[997] * mat_B[167] +
//             mat_A[998] * mat_B[199] +
//             mat_A[999] * mat_B[231] +
//             mat_A[1000] * mat_B[263] +
//             mat_A[1001] * mat_B[295] +
//             mat_A[1002] * mat_B[327] +
//             mat_A[1003] * mat_B[359] +
//             mat_A[1004] * mat_B[391] +
//             mat_A[1005] * mat_B[423] +
//             mat_A[1006] * mat_B[455] +
//             mat_A[1007] * mat_B[487] +
//             mat_A[1008] * mat_B[519] +
//             mat_A[1009] * mat_B[551] +
//             mat_A[1010] * mat_B[583] +
//             mat_A[1011] * mat_B[615] +
//             mat_A[1012] * mat_B[647] +
//             mat_A[1013] * mat_B[679] +
//             mat_A[1014] * mat_B[711] +
//             mat_A[1015] * mat_B[743] +
//             mat_A[1016] * mat_B[775] +
//             mat_A[1017] * mat_B[807] +
//             mat_A[1018] * mat_B[839] +
//             mat_A[1019] * mat_B[871] +
//             mat_A[1020] * mat_B[903] +
//             mat_A[1021] * mat_B[935] +
//             mat_A[1022] * mat_B[967] +
//             mat_A[1023] * mat_B[999];
//  mat_C[1000] <= 
//             mat_A[992] * mat_B[8] +
//             mat_A[993] * mat_B[40] +
//             mat_A[994] * mat_B[72] +
//             mat_A[995] * mat_B[104] +
//             mat_A[996] * mat_B[136] +
//             mat_A[997] * mat_B[168] +
//             mat_A[998] * mat_B[200] +
//             mat_A[999] * mat_B[232] +
//             mat_A[1000] * mat_B[264] +
//             mat_A[1001] * mat_B[296] +
//             mat_A[1002] * mat_B[328] +
//             mat_A[1003] * mat_B[360] +
//             mat_A[1004] * mat_B[392] +
//             mat_A[1005] * mat_B[424] +
//             mat_A[1006] * mat_B[456] +
//             mat_A[1007] * mat_B[488] +
//             mat_A[1008] * mat_B[520] +
//             mat_A[1009] * mat_B[552] +
//             mat_A[1010] * mat_B[584] +
//             mat_A[1011] * mat_B[616] +
//             mat_A[1012] * mat_B[648] +
//             mat_A[1013] * mat_B[680] +
//             mat_A[1014] * mat_B[712] +
//             mat_A[1015] * mat_B[744] +
//             mat_A[1016] * mat_B[776] +
//             mat_A[1017] * mat_B[808] +
//             mat_A[1018] * mat_B[840] +
//             mat_A[1019] * mat_B[872] +
//             mat_A[1020] * mat_B[904] +
//             mat_A[1021] * mat_B[936] +
//             mat_A[1022] * mat_B[968] +
//             mat_A[1023] * mat_B[1000];
//  mat_C[1001] <= 
//             mat_A[992] * mat_B[9] +
//             mat_A[993] * mat_B[41] +
//             mat_A[994] * mat_B[73] +
//             mat_A[995] * mat_B[105] +
//             mat_A[996] * mat_B[137] +
//             mat_A[997] * mat_B[169] +
//             mat_A[998] * mat_B[201] +
//             mat_A[999] * mat_B[233] +
//             mat_A[1000] * mat_B[265] +
//             mat_A[1001] * mat_B[297] +
//             mat_A[1002] * mat_B[329] +
//             mat_A[1003] * mat_B[361] +
//             mat_A[1004] * mat_B[393] +
//             mat_A[1005] * mat_B[425] +
//             mat_A[1006] * mat_B[457] +
//             mat_A[1007] * mat_B[489] +
//             mat_A[1008] * mat_B[521] +
//             mat_A[1009] * mat_B[553] +
//             mat_A[1010] * mat_B[585] +
//             mat_A[1011] * mat_B[617] +
//             mat_A[1012] * mat_B[649] +
//             mat_A[1013] * mat_B[681] +
//             mat_A[1014] * mat_B[713] +
//             mat_A[1015] * mat_B[745] +
//             mat_A[1016] * mat_B[777] +
//             mat_A[1017] * mat_B[809] +
//             mat_A[1018] * mat_B[841] +
//             mat_A[1019] * mat_B[873] +
//             mat_A[1020] * mat_B[905] +
//             mat_A[1021] * mat_B[937] +
//             mat_A[1022] * mat_B[969] +
//             mat_A[1023] * mat_B[1001];
//  mat_C[1002] <= 
//             mat_A[992] * mat_B[10] +
//             mat_A[993] * mat_B[42] +
//             mat_A[994] * mat_B[74] +
//             mat_A[995] * mat_B[106] +
//             mat_A[996] * mat_B[138] +
//             mat_A[997] * mat_B[170] +
//             mat_A[998] * mat_B[202] +
//             mat_A[999] * mat_B[234] +
//             mat_A[1000] * mat_B[266] +
//             mat_A[1001] * mat_B[298] +
//             mat_A[1002] * mat_B[330] +
//             mat_A[1003] * mat_B[362] +
//             mat_A[1004] * mat_B[394] +
//             mat_A[1005] * mat_B[426] +
//             mat_A[1006] * mat_B[458] +
//             mat_A[1007] * mat_B[490] +
//             mat_A[1008] * mat_B[522] +
//             mat_A[1009] * mat_B[554] +
//             mat_A[1010] * mat_B[586] +
//             mat_A[1011] * mat_B[618] +
//             mat_A[1012] * mat_B[650] +
//             mat_A[1013] * mat_B[682] +
//             mat_A[1014] * mat_B[714] +
//             mat_A[1015] * mat_B[746] +
//             mat_A[1016] * mat_B[778] +
//             mat_A[1017] * mat_B[810] +
//             mat_A[1018] * mat_B[842] +
//             mat_A[1019] * mat_B[874] +
//             mat_A[1020] * mat_B[906] +
//             mat_A[1021] * mat_B[938] +
//             mat_A[1022] * mat_B[970] +
//             mat_A[1023] * mat_B[1002];
//  mat_C[1003] <= 
//             mat_A[992] * mat_B[11] +
//             mat_A[993] * mat_B[43] +
//             mat_A[994] * mat_B[75] +
//             mat_A[995] * mat_B[107] +
//             mat_A[996] * mat_B[139] +
//             mat_A[997] * mat_B[171] +
//             mat_A[998] * mat_B[203] +
//             mat_A[999] * mat_B[235] +
//             mat_A[1000] * mat_B[267] +
//             mat_A[1001] * mat_B[299] +
//             mat_A[1002] * mat_B[331] +
//             mat_A[1003] * mat_B[363] +
//             mat_A[1004] * mat_B[395] +
//             mat_A[1005] * mat_B[427] +
//             mat_A[1006] * mat_B[459] +
//             mat_A[1007] * mat_B[491] +
//             mat_A[1008] * mat_B[523] +
//             mat_A[1009] * mat_B[555] +
//             mat_A[1010] * mat_B[587] +
//             mat_A[1011] * mat_B[619] +
//             mat_A[1012] * mat_B[651] +
//             mat_A[1013] * mat_B[683] +
//             mat_A[1014] * mat_B[715] +
//             mat_A[1015] * mat_B[747] +
//             mat_A[1016] * mat_B[779] +
//             mat_A[1017] * mat_B[811] +
//             mat_A[1018] * mat_B[843] +
//             mat_A[1019] * mat_B[875] +
//             mat_A[1020] * mat_B[907] +
//             mat_A[1021] * mat_B[939] +
//             mat_A[1022] * mat_B[971] +
//             mat_A[1023] * mat_B[1003];
//  mat_C[1004] <= 
//             mat_A[992] * mat_B[12] +
//             mat_A[993] * mat_B[44] +
//             mat_A[994] * mat_B[76] +
//             mat_A[995] * mat_B[108] +
//             mat_A[996] * mat_B[140] +
//             mat_A[997] * mat_B[172] +
//             mat_A[998] * mat_B[204] +
//             mat_A[999] * mat_B[236] +
//             mat_A[1000] * mat_B[268] +
//             mat_A[1001] * mat_B[300] +
//             mat_A[1002] * mat_B[332] +
//             mat_A[1003] * mat_B[364] +
//             mat_A[1004] * mat_B[396] +
//             mat_A[1005] * mat_B[428] +
//             mat_A[1006] * mat_B[460] +
//             mat_A[1007] * mat_B[492] +
//             mat_A[1008] * mat_B[524] +
//             mat_A[1009] * mat_B[556] +
//             mat_A[1010] * mat_B[588] +
//             mat_A[1011] * mat_B[620] +
//             mat_A[1012] * mat_B[652] +
//             mat_A[1013] * mat_B[684] +
//             mat_A[1014] * mat_B[716] +
//             mat_A[1015] * mat_B[748] +
//             mat_A[1016] * mat_B[780] +
//             mat_A[1017] * mat_B[812] +
//             mat_A[1018] * mat_B[844] +
//             mat_A[1019] * mat_B[876] +
//             mat_A[1020] * mat_B[908] +
//             mat_A[1021] * mat_B[940] +
//             mat_A[1022] * mat_B[972] +
//             mat_A[1023] * mat_B[1004];
//  mat_C[1005] <= 
//             mat_A[992] * mat_B[13] +
//             mat_A[993] * mat_B[45] +
//             mat_A[994] * mat_B[77] +
//             mat_A[995] * mat_B[109] +
//             mat_A[996] * mat_B[141] +
//             mat_A[997] * mat_B[173] +
//             mat_A[998] * mat_B[205] +
//             mat_A[999] * mat_B[237] +
//             mat_A[1000] * mat_B[269] +
//             mat_A[1001] * mat_B[301] +
//             mat_A[1002] * mat_B[333] +
//             mat_A[1003] * mat_B[365] +
//             mat_A[1004] * mat_B[397] +
//             mat_A[1005] * mat_B[429] +
//             mat_A[1006] * mat_B[461] +
//             mat_A[1007] * mat_B[493] +
//             mat_A[1008] * mat_B[525] +
//             mat_A[1009] * mat_B[557] +
//             mat_A[1010] * mat_B[589] +
//             mat_A[1011] * mat_B[621] +
//             mat_A[1012] * mat_B[653] +
//             mat_A[1013] * mat_B[685] +
//             mat_A[1014] * mat_B[717] +
//             mat_A[1015] * mat_B[749] +
//             mat_A[1016] * mat_B[781] +
//             mat_A[1017] * mat_B[813] +
//             mat_A[1018] * mat_B[845] +
//             mat_A[1019] * mat_B[877] +
//             mat_A[1020] * mat_B[909] +
//             mat_A[1021] * mat_B[941] +
//             mat_A[1022] * mat_B[973] +
//             mat_A[1023] * mat_B[1005];
//  mat_C[1006] <= 
//             mat_A[992] * mat_B[14] +
//             mat_A[993] * mat_B[46] +
//             mat_A[994] * mat_B[78] +
//             mat_A[995] * mat_B[110] +
//             mat_A[996] * mat_B[142] +
//             mat_A[997] * mat_B[174] +
//             mat_A[998] * mat_B[206] +
//             mat_A[999] * mat_B[238] +
//             mat_A[1000] * mat_B[270] +
//             mat_A[1001] * mat_B[302] +
//             mat_A[1002] * mat_B[334] +
//             mat_A[1003] * mat_B[366] +
//             mat_A[1004] * mat_B[398] +
//             mat_A[1005] * mat_B[430] +
//             mat_A[1006] * mat_B[462] +
//             mat_A[1007] * mat_B[494] +
//             mat_A[1008] * mat_B[526] +
//             mat_A[1009] * mat_B[558] +
//             mat_A[1010] * mat_B[590] +
//             mat_A[1011] * mat_B[622] +
//             mat_A[1012] * mat_B[654] +
//             mat_A[1013] * mat_B[686] +
//             mat_A[1014] * mat_B[718] +
//             mat_A[1015] * mat_B[750] +
//             mat_A[1016] * mat_B[782] +
//             mat_A[1017] * mat_B[814] +
//             mat_A[1018] * mat_B[846] +
//             mat_A[1019] * mat_B[878] +
//             mat_A[1020] * mat_B[910] +
//             mat_A[1021] * mat_B[942] +
//             mat_A[1022] * mat_B[974] +
//             mat_A[1023] * mat_B[1006];
//  mat_C[1007] <= 
//             mat_A[992] * mat_B[15] +
//             mat_A[993] * mat_B[47] +
//             mat_A[994] * mat_B[79] +
//             mat_A[995] * mat_B[111] +
//             mat_A[996] * mat_B[143] +
//             mat_A[997] * mat_B[175] +
//             mat_A[998] * mat_B[207] +
//             mat_A[999] * mat_B[239] +
//             mat_A[1000] * mat_B[271] +
//             mat_A[1001] * mat_B[303] +
//             mat_A[1002] * mat_B[335] +
//             mat_A[1003] * mat_B[367] +
//             mat_A[1004] * mat_B[399] +
//             mat_A[1005] * mat_B[431] +
//             mat_A[1006] * mat_B[463] +
//             mat_A[1007] * mat_B[495] +
//             mat_A[1008] * mat_B[527] +
//             mat_A[1009] * mat_B[559] +
//             mat_A[1010] * mat_B[591] +
//             mat_A[1011] * mat_B[623] +
//             mat_A[1012] * mat_B[655] +
//             mat_A[1013] * mat_B[687] +
//             mat_A[1014] * mat_B[719] +
//             mat_A[1015] * mat_B[751] +
//             mat_A[1016] * mat_B[783] +
//             mat_A[1017] * mat_B[815] +
//             mat_A[1018] * mat_B[847] +
//             mat_A[1019] * mat_B[879] +
//             mat_A[1020] * mat_B[911] +
//             mat_A[1021] * mat_B[943] +
//             mat_A[1022] * mat_B[975] +
//             mat_A[1023] * mat_B[1007];
//  mat_C[1008] <= 
//             mat_A[992] * mat_B[16] +
//             mat_A[993] * mat_B[48] +
//             mat_A[994] * mat_B[80] +
//             mat_A[995] * mat_B[112] +
//             mat_A[996] * mat_B[144] +
//             mat_A[997] * mat_B[176] +
//             mat_A[998] * mat_B[208] +
//             mat_A[999] * mat_B[240] +
//             mat_A[1000] * mat_B[272] +
//             mat_A[1001] * mat_B[304] +
//             mat_A[1002] * mat_B[336] +
//             mat_A[1003] * mat_B[368] +
//             mat_A[1004] * mat_B[400] +
//             mat_A[1005] * mat_B[432] +
//             mat_A[1006] * mat_B[464] +
//             mat_A[1007] * mat_B[496] +
//             mat_A[1008] * mat_B[528] +
//             mat_A[1009] * mat_B[560] +
//             mat_A[1010] * mat_B[592] +
//             mat_A[1011] * mat_B[624] +
//             mat_A[1012] * mat_B[656] +
//             mat_A[1013] * mat_B[688] +
//             mat_A[1014] * mat_B[720] +
//             mat_A[1015] * mat_B[752] +
//             mat_A[1016] * mat_B[784] +
//             mat_A[1017] * mat_B[816] +
//             mat_A[1018] * mat_B[848] +
//             mat_A[1019] * mat_B[880] +
//             mat_A[1020] * mat_B[912] +
//             mat_A[1021] * mat_B[944] +
//             mat_A[1022] * mat_B[976] +
//             mat_A[1023] * mat_B[1008];
//  mat_C[1009] <= 
//             mat_A[992] * mat_B[17] +
//             mat_A[993] * mat_B[49] +
//             mat_A[994] * mat_B[81] +
//             mat_A[995] * mat_B[113] +
//             mat_A[996] * mat_B[145] +
//             mat_A[997] * mat_B[177] +
//             mat_A[998] * mat_B[209] +
//             mat_A[999] * mat_B[241] +
//             mat_A[1000] * mat_B[273] +
//             mat_A[1001] * mat_B[305] +
//             mat_A[1002] * mat_B[337] +
//             mat_A[1003] * mat_B[369] +
//             mat_A[1004] * mat_B[401] +
//             mat_A[1005] * mat_B[433] +
//             mat_A[1006] * mat_B[465] +
//             mat_A[1007] * mat_B[497] +
//             mat_A[1008] * mat_B[529] +
//             mat_A[1009] * mat_B[561] +
//             mat_A[1010] * mat_B[593] +
//             mat_A[1011] * mat_B[625] +
//             mat_A[1012] * mat_B[657] +
//             mat_A[1013] * mat_B[689] +
//             mat_A[1014] * mat_B[721] +
//             mat_A[1015] * mat_B[753] +
//             mat_A[1016] * mat_B[785] +
//             mat_A[1017] * mat_B[817] +
//             mat_A[1018] * mat_B[849] +
//             mat_A[1019] * mat_B[881] +
//             mat_A[1020] * mat_B[913] +
//             mat_A[1021] * mat_B[945] +
//             mat_A[1022] * mat_B[977] +
//             mat_A[1023] * mat_B[1009];
//  mat_C[1010] <= 
//             mat_A[992] * mat_B[18] +
//             mat_A[993] * mat_B[50] +
//             mat_A[994] * mat_B[82] +
//             mat_A[995] * mat_B[114] +
//             mat_A[996] * mat_B[146] +
//             mat_A[997] * mat_B[178] +
//             mat_A[998] * mat_B[210] +
//             mat_A[999] * mat_B[242] +
//             mat_A[1000] * mat_B[274] +
//             mat_A[1001] * mat_B[306] +
//             mat_A[1002] * mat_B[338] +
//             mat_A[1003] * mat_B[370] +
//             mat_A[1004] * mat_B[402] +
//             mat_A[1005] * mat_B[434] +
//             mat_A[1006] * mat_B[466] +
//             mat_A[1007] * mat_B[498] +
//             mat_A[1008] * mat_B[530] +
//             mat_A[1009] * mat_B[562] +
//             mat_A[1010] * mat_B[594] +
//             mat_A[1011] * mat_B[626] +
//             mat_A[1012] * mat_B[658] +
//             mat_A[1013] * mat_B[690] +
//             mat_A[1014] * mat_B[722] +
//             mat_A[1015] * mat_B[754] +
//             mat_A[1016] * mat_B[786] +
//             mat_A[1017] * mat_B[818] +
//             mat_A[1018] * mat_B[850] +
//             mat_A[1019] * mat_B[882] +
//             mat_A[1020] * mat_B[914] +
//             mat_A[1021] * mat_B[946] +
//             mat_A[1022] * mat_B[978] +
//             mat_A[1023] * mat_B[1010];
//  mat_C[1011] <= 
//             mat_A[992] * mat_B[19] +
//             mat_A[993] * mat_B[51] +
//             mat_A[994] * mat_B[83] +
//             mat_A[995] * mat_B[115] +
//             mat_A[996] * mat_B[147] +
//             mat_A[997] * mat_B[179] +
//             mat_A[998] * mat_B[211] +
//             mat_A[999] * mat_B[243] +
//             mat_A[1000] * mat_B[275] +
//             mat_A[1001] * mat_B[307] +
//             mat_A[1002] * mat_B[339] +
//             mat_A[1003] * mat_B[371] +
//             mat_A[1004] * mat_B[403] +
//             mat_A[1005] * mat_B[435] +
//             mat_A[1006] * mat_B[467] +
//             mat_A[1007] * mat_B[499] +
//             mat_A[1008] * mat_B[531] +
//             mat_A[1009] * mat_B[563] +
//             mat_A[1010] * mat_B[595] +
//             mat_A[1011] * mat_B[627] +
//             mat_A[1012] * mat_B[659] +
//             mat_A[1013] * mat_B[691] +
//             mat_A[1014] * mat_B[723] +
//             mat_A[1015] * mat_B[755] +
//             mat_A[1016] * mat_B[787] +
//             mat_A[1017] * mat_B[819] +
//             mat_A[1018] * mat_B[851] +
//             mat_A[1019] * mat_B[883] +
//             mat_A[1020] * mat_B[915] +
//             mat_A[1021] * mat_B[947] +
//             mat_A[1022] * mat_B[979] +
//             mat_A[1023] * mat_B[1011];
//  mat_C[1012] <= 
//             mat_A[992] * mat_B[20] +
//             mat_A[993] * mat_B[52] +
//             mat_A[994] * mat_B[84] +
//             mat_A[995] * mat_B[116] +
//             mat_A[996] * mat_B[148] +
//             mat_A[997] * mat_B[180] +
//             mat_A[998] * mat_B[212] +
//             mat_A[999] * mat_B[244] +
//             mat_A[1000] * mat_B[276] +
//             mat_A[1001] * mat_B[308] +
//             mat_A[1002] * mat_B[340] +
//             mat_A[1003] * mat_B[372] +
//             mat_A[1004] * mat_B[404] +
//             mat_A[1005] * mat_B[436] +
//             mat_A[1006] * mat_B[468] +
//             mat_A[1007] * mat_B[500] +
//             mat_A[1008] * mat_B[532] +
//             mat_A[1009] * mat_B[564] +
//             mat_A[1010] * mat_B[596] +
//             mat_A[1011] * mat_B[628] +
//             mat_A[1012] * mat_B[660] +
//             mat_A[1013] * mat_B[692] +
//             mat_A[1014] * mat_B[724] +
//             mat_A[1015] * mat_B[756] +
//             mat_A[1016] * mat_B[788] +
//             mat_A[1017] * mat_B[820] +
//             mat_A[1018] * mat_B[852] +
//             mat_A[1019] * mat_B[884] +
//             mat_A[1020] * mat_B[916] +
//             mat_A[1021] * mat_B[948] +
//             mat_A[1022] * mat_B[980] +
//             mat_A[1023] * mat_B[1012];
//  mat_C[1013] <= 
//             mat_A[992] * mat_B[21] +
//             mat_A[993] * mat_B[53] +
//             mat_A[994] * mat_B[85] +
//             mat_A[995] * mat_B[117] +
//             mat_A[996] * mat_B[149] +
//             mat_A[997] * mat_B[181] +
//             mat_A[998] * mat_B[213] +
//             mat_A[999] * mat_B[245] +
//             mat_A[1000] * mat_B[277] +
//             mat_A[1001] * mat_B[309] +
//             mat_A[1002] * mat_B[341] +
//             mat_A[1003] * mat_B[373] +
//             mat_A[1004] * mat_B[405] +
//             mat_A[1005] * mat_B[437] +
//             mat_A[1006] * mat_B[469] +
//             mat_A[1007] * mat_B[501] +
//             mat_A[1008] * mat_B[533] +
//             mat_A[1009] * mat_B[565] +
//             mat_A[1010] * mat_B[597] +
//             mat_A[1011] * mat_B[629] +
//             mat_A[1012] * mat_B[661] +
//             mat_A[1013] * mat_B[693] +
//             mat_A[1014] * mat_B[725] +
//             mat_A[1015] * mat_B[757] +
//             mat_A[1016] * mat_B[789] +
//             mat_A[1017] * mat_B[821] +
//             mat_A[1018] * mat_B[853] +
//             mat_A[1019] * mat_B[885] +
//             mat_A[1020] * mat_B[917] +
//             mat_A[1021] * mat_B[949] +
//             mat_A[1022] * mat_B[981] +
//             mat_A[1023] * mat_B[1013];
//  mat_C[1014] <= 
//             mat_A[992] * mat_B[22] +
//             mat_A[993] * mat_B[54] +
//             mat_A[994] * mat_B[86] +
//             mat_A[995] * mat_B[118] +
//             mat_A[996] * mat_B[150] +
//             mat_A[997] * mat_B[182] +
//             mat_A[998] * mat_B[214] +
//             mat_A[999] * mat_B[246] +
//             mat_A[1000] * mat_B[278] +
//             mat_A[1001] * mat_B[310] +
//             mat_A[1002] * mat_B[342] +
//             mat_A[1003] * mat_B[374] +
//             mat_A[1004] * mat_B[406] +
//             mat_A[1005] * mat_B[438] +
//             mat_A[1006] * mat_B[470] +
//             mat_A[1007] * mat_B[502] +
//             mat_A[1008] * mat_B[534] +
//             mat_A[1009] * mat_B[566] +
//             mat_A[1010] * mat_B[598] +
//             mat_A[1011] * mat_B[630] +
//             mat_A[1012] * mat_B[662] +
//             mat_A[1013] * mat_B[694] +
//             mat_A[1014] * mat_B[726] +
//             mat_A[1015] * mat_B[758] +
//             mat_A[1016] * mat_B[790] +
//             mat_A[1017] * mat_B[822] +
//             mat_A[1018] * mat_B[854] +
//             mat_A[1019] * mat_B[886] +
//             mat_A[1020] * mat_B[918] +
//             mat_A[1021] * mat_B[950] +
//             mat_A[1022] * mat_B[982] +
//             mat_A[1023] * mat_B[1014];
//  mat_C[1015] <= 
//             mat_A[992] * mat_B[23] +
//             mat_A[993] * mat_B[55] +
//             mat_A[994] * mat_B[87] +
//             mat_A[995] * mat_B[119] +
//             mat_A[996] * mat_B[151] +
//             mat_A[997] * mat_B[183] +
//             mat_A[998] * mat_B[215] +
//             mat_A[999] * mat_B[247] +
//             mat_A[1000] * mat_B[279] +
//             mat_A[1001] * mat_B[311] +
//             mat_A[1002] * mat_B[343] +
//             mat_A[1003] * mat_B[375] +
//             mat_A[1004] * mat_B[407] +
//             mat_A[1005] * mat_B[439] +
//             mat_A[1006] * mat_B[471] +
//             mat_A[1007] * mat_B[503] +
//             mat_A[1008] * mat_B[535] +
//             mat_A[1009] * mat_B[567] +
//             mat_A[1010] * mat_B[599] +
//             mat_A[1011] * mat_B[631] +
//             mat_A[1012] * mat_B[663] +
//             mat_A[1013] * mat_B[695] +
//             mat_A[1014] * mat_B[727] +
//             mat_A[1015] * mat_B[759] +
//             mat_A[1016] * mat_B[791] +
//             mat_A[1017] * mat_B[823] +
//             mat_A[1018] * mat_B[855] +
//             mat_A[1019] * mat_B[887] +
//             mat_A[1020] * mat_B[919] +
//             mat_A[1021] * mat_B[951] +
//             mat_A[1022] * mat_B[983] +
//             mat_A[1023] * mat_B[1015];
//  mat_C[1016] <= 
//             mat_A[992] * mat_B[24] +
//             mat_A[993] * mat_B[56] +
//             mat_A[994] * mat_B[88] +
//             mat_A[995] * mat_B[120] +
//             mat_A[996] * mat_B[152] +
//             mat_A[997] * mat_B[184] +
//             mat_A[998] * mat_B[216] +
//             mat_A[999] * mat_B[248] +
//             mat_A[1000] * mat_B[280] +
//             mat_A[1001] * mat_B[312] +
//             mat_A[1002] * mat_B[344] +
//             mat_A[1003] * mat_B[376] +
//             mat_A[1004] * mat_B[408] +
//             mat_A[1005] * mat_B[440] +
//             mat_A[1006] * mat_B[472] +
//             mat_A[1007] * mat_B[504] +
//             mat_A[1008] * mat_B[536] +
//             mat_A[1009] * mat_B[568] +
//             mat_A[1010] * mat_B[600] +
//             mat_A[1011] * mat_B[632] +
//             mat_A[1012] * mat_B[664] +
//             mat_A[1013] * mat_B[696] +
//             mat_A[1014] * mat_B[728] +
//             mat_A[1015] * mat_B[760] +
//             mat_A[1016] * mat_B[792] +
//             mat_A[1017] * mat_B[824] +
//             mat_A[1018] * mat_B[856] +
//             mat_A[1019] * mat_B[888] +
//             mat_A[1020] * mat_B[920] +
//             mat_A[1021] * mat_B[952] +
//             mat_A[1022] * mat_B[984] +
//             mat_A[1023] * mat_B[1016];
//  mat_C[1017] <= 
//             mat_A[992] * mat_B[25] +
//             mat_A[993] * mat_B[57] +
//             mat_A[994] * mat_B[89] +
//             mat_A[995] * mat_B[121] +
//             mat_A[996] * mat_B[153] +
//             mat_A[997] * mat_B[185] +
//             mat_A[998] * mat_B[217] +
//             mat_A[999] * mat_B[249] +
//             mat_A[1000] * mat_B[281] +
//             mat_A[1001] * mat_B[313] +
//             mat_A[1002] * mat_B[345] +
//             mat_A[1003] * mat_B[377] +
//             mat_A[1004] * mat_B[409] +
//             mat_A[1005] * mat_B[441] +
//             mat_A[1006] * mat_B[473] +
//             mat_A[1007] * mat_B[505] +
//             mat_A[1008] * mat_B[537] +
//             mat_A[1009] * mat_B[569] +
//             mat_A[1010] * mat_B[601] +
//             mat_A[1011] * mat_B[633] +
//             mat_A[1012] * mat_B[665] +
//             mat_A[1013] * mat_B[697] +
//             mat_A[1014] * mat_B[729] +
//             mat_A[1015] * mat_B[761] +
//             mat_A[1016] * mat_B[793] +
//             mat_A[1017] * mat_B[825] +
//             mat_A[1018] * mat_B[857] +
//             mat_A[1019] * mat_B[889] +
//             mat_A[1020] * mat_B[921] +
//             mat_A[1021] * mat_B[953] +
//             mat_A[1022] * mat_B[985] +
//             mat_A[1023] * mat_B[1017];
//  mat_C[1018] <= 
//             mat_A[992] * mat_B[26] +
//             mat_A[993] * mat_B[58] +
//             mat_A[994] * mat_B[90] +
//             mat_A[995] * mat_B[122] +
//             mat_A[996] * mat_B[154] +
//             mat_A[997] * mat_B[186] +
//             mat_A[998] * mat_B[218] +
//             mat_A[999] * mat_B[250] +
//             mat_A[1000] * mat_B[282] +
//             mat_A[1001] * mat_B[314] +
//             mat_A[1002] * mat_B[346] +
//             mat_A[1003] * mat_B[378] +
//             mat_A[1004] * mat_B[410] +
//             mat_A[1005] * mat_B[442] +
//             mat_A[1006] * mat_B[474] +
//             mat_A[1007] * mat_B[506] +
//             mat_A[1008] * mat_B[538] +
//             mat_A[1009] * mat_B[570] +
//             mat_A[1010] * mat_B[602] +
//             mat_A[1011] * mat_B[634] +
//             mat_A[1012] * mat_B[666] +
//             mat_A[1013] * mat_B[698] +
//             mat_A[1014] * mat_B[730] +
//             mat_A[1015] * mat_B[762] +
//             mat_A[1016] * mat_B[794] +
//             mat_A[1017] * mat_B[826] +
//             mat_A[1018] * mat_B[858] +
//             mat_A[1019] * mat_B[890] +
//             mat_A[1020] * mat_B[922] +
//             mat_A[1021] * mat_B[954] +
//             mat_A[1022] * mat_B[986] +
//             mat_A[1023] * mat_B[1018];
//  mat_C[1019] <= 
//             mat_A[992] * mat_B[27] +
//             mat_A[993] * mat_B[59] +
//             mat_A[994] * mat_B[91] +
//             mat_A[995] * mat_B[123] +
//             mat_A[996] * mat_B[155] +
//             mat_A[997] * mat_B[187] +
//             mat_A[998] * mat_B[219] +
//             mat_A[999] * mat_B[251] +
//             mat_A[1000] * mat_B[283] +
//             mat_A[1001] * mat_B[315] +
//             mat_A[1002] * mat_B[347] +
//             mat_A[1003] * mat_B[379] +
//             mat_A[1004] * mat_B[411] +
//             mat_A[1005] * mat_B[443] +
//             mat_A[1006] * mat_B[475] +
//             mat_A[1007] * mat_B[507] +
//             mat_A[1008] * mat_B[539] +
//             mat_A[1009] * mat_B[571] +
//             mat_A[1010] * mat_B[603] +
//             mat_A[1011] * mat_B[635] +
//             mat_A[1012] * mat_B[667] +
//             mat_A[1013] * mat_B[699] +
//             mat_A[1014] * mat_B[731] +
//             mat_A[1015] * mat_B[763] +
//             mat_A[1016] * mat_B[795] +
//             mat_A[1017] * mat_B[827] +
//             mat_A[1018] * mat_B[859] +
//             mat_A[1019] * mat_B[891] +
//             mat_A[1020] * mat_B[923] +
//             mat_A[1021] * mat_B[955] +
//             mat_A[1022] * mat_B[987] +
//             mat_A[1023] * mat_B[1019];
//  mat_C[1020] <= 
//             mat_A[992] * mat_B[28] +
//             mat_A[993] * mat_B[60] +
//             mat_A[994] * mat_B[92] +
//             mat_A[995] * mat_B[124] +
//             mat_A[996] * mat_B[156] +
//             mat_A[997] * mat_B[188] +
//             mat_A[998] * mat_B[220] +
//             mat_A[999] * mat_B[252] +
//             mat_A[1000] * mat_B[284] +
//             mat_A[1001] * mat_B[316] +
//             mat_A[1002] * mat_B[348] +
//             mat_A[1003] * mat_B[380] +
//             mat_A[1004] * mat_B[412] +
//             mat_A[1005] * mat_B[444] +
//             mat_A[1006] * mat_B[476] +
//             mat_A[1007] * mat_B[508] +
//             mat_A[1008] * mat_B[540] +
//             mat_A[1009] * mat_B[572] +
//             mat_A[1010] * mat_B[604] +
//             mat_A[1011] * mat_B[636] +
//             mat_A[1012] * mat_B[668] +
//             mat_A[1013] * mat_B[700] +
//             mat_A[1014] * mat_B[732] +
//             mat_A[1015] * mat_B[764] +
//             mat_A[1016] * mat_B[796] +
//             mat_A[1017] * mat_B[828] +
//             mat_A[1018] * mat_B[860] +
//             mat_A[1019] * mat_B[892] +
//             mat_A[1020] * mat_B[924] +
//             mat_A[1021] * mat_B[956] +
//             mat_A[1022] * mat_B[988] +
//             mat_A[1023] * mat_B[1020];
//  mat_C[1021] <= 
//             mat_A[992] * mat_B[29] +
//             mat_A[993] * mat_B[61] +
//             mat_A[994] * mat_B[93] +
//             mat_A[995] * mat_B[125] +
//             mat_A[996] * mat_B[157] +
//             mat_A[997] * mat_B[189] +
//             mat_A[998] * mat_B[221] +
//             mat_A[999] * mat_B[253] +
//             mat_A[1000] * mat_B[285] +
//             mat_A[1001] * mat_B[317] +
//             mat_A[1002] * mat_B[349] +
//             mat_A[1003] * mat_B[381] +
//             mat_A[1004] * mat_B[413] +
//             mat_A[1005] * mat_B[445] +
//             mat_A[1006] * mat_B[477] +
//             mat_A[1007] * mat_B[509] +
//             mat_A[1008] * mat_B[541] +
//             mat_A[1009] * mat_B[573] +
//             mat_A[1010] * mat_B[605] +
//             mat_A[1011] * mat_B[637] +
//             mat_A[1012] * mat_B[669] +
//             mat_A[1013] * mat_B[701] +
//             mat_A[1014] * mat_B[733] +
//             mat_A[1015] * mat_B[765] +
//             mat_A[1016] * mat_B[797] +
//             mat_A[1017] * mat_B[829] +
//             mat_A[1018] * mat_B[861] +
//             mat_A[1019] * mat_B[893] +
//             mat_A[1020] * mat_B[925] +
//             mat_A[1021] * mat_B[957] +
//             mat_A[1022] * mat_B[989] +
//             mat_A[1023] * mat_B[1021];
//  mat_C[1022] <= 
//             mat_A[992] * mat_B[30] +
//             mat_A[993] * mat_B[62] +
//             mat_A[994] * mat_B[94] +
//             mat_A[995] * mat_B[126] +
//             mat_A[996] * mat_B[158] +
//             mat_A[997] * mat_B[190] +
//             mat_A[998] * mat_B[222] +
//             mat_A[999] * mat_B[254] +
//             mat_A[1000] * mat_B[286] +
//             mat_A[1001] * mat_B[318] +
//             mat_A[1002] * mat_B[350] +
//             mat_A[1003] * mat_B[382] +
//             mat_A[1004] * mat_B[414] +
//             mat_A[1005] * mat_B[446] +
//             mat_A[1006] * mat_B[478] +
//             mat_A[1007] * mat_B[510] +
//             mat_A[1008] * mat_B[542] +
//             mat_A[1009] * mat_B[574] +
//             mat_A[1010] * mat_B[606] +
//             mat_A[1011] * mat_B[638] +
//             mat_A[1012] * mat_B[670] +
//             mat_A[1013] * mat_B[702] +
//             mat_A[1014] * mat_B[734] +
//             mat_A[1015] * mat_B[766] +
//             mat_A[1016] * mat_B[798] +
//             mat_A[1017] * mat_B[830] +
//             mat_A[1018] * mat_B[862] +
//             mat_A[1019] * mat_B[894] +
//             mat_A[1020] * mat_B[926] +
//             mat_A[1021] * mat_B[958] +
//             mat_A[1022] * mat_B[990] +
//             mat_A[1023] * mat_B[1022];
//  mat_C[1023] <= 
//             mat_A[992] * mat_B[31] +
//             mat_A[993] * mat_B[63] +
//             mat_A[994] * mat_B[95] +
//             mat_A[995] * mat_B[127] +
//             mat_A[996] * mat_B[159] +
//             mat_A[997] * mat_B[191] +
//             mat_A[998] * mat_B[223] +
//             mat_A[999] * mat_B[255] +
//             mat_A[1000] * mat_B[287] +
//             mat_A[1001] * mat_B[319] +
//             mat_A[1002] * mat_B[351] +
//             mat_A[1003] * mat_B[383] +
//             mat_A[1004] * mat_B[415] +
//             mat_A[1005] * mat_B[447] +
//             mat_A[1006] * mat_B[479] +
//             mat_A[1007] * mat_B[511] +
//             mat_A[1008] * mat_B[543] +
//             mat_A[1009] * mat_B[575] +
//             mat_A[1010] * mat_B[607] +
//             mat_A[1011] * mat_B[639] +
//             mat_A[1012] * mat_B[671] +
//             mat_A[1013] * mat_B[703] +
//             mat_A[1014] * mat_B[735] +
//             mat_A[1015] * mat_B[767] +
//             mat_A[1016] * mat_B[799] +
//             mat_A[1017] * mat_B[831] +
//             mat_A[1018] * mat_B[863] +
//             mat_A[1019] * mat_B[895] +
//             mat_A[1020] * mat_B[927] +
//             mat_A[1021] * mat_B[959] +
//             mat_A[1022] * mat_B[991] +
//             mat_A[1023] * mat_B[1023];
  end
endmodule
