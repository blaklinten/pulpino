module multiply_long #(
  parameter mat_size = 2,
  parameter dat_size = 8
) (
  input  logic            start        ,
  input  logic            clk          , //kanske ej behövs
  input  logic [3:0][7:0] mat_A [255:0],
  input  logic [3:0][7:0] mat_B [255:0],
  output logic [3:0][7:0] mat_C [255:0],
  output logic            done
);

  always @(posedge clk)
  begin
    mat_C[0][0] <= 
                  mat_A[0][0] * mat_B[0][0] +
                  mat_A[0][1] * mat_B[1][0] +
                  mat_A[0][2] * mat_B[2][0] +
                  mat_A[0][3] * mat_B[3][0] +
                  mat_A[0][4] * mat_B[4][0] +
                  mat_A[0][5] * mat_B[5][0] +
                  mat_A[0][6] * mat_B[6][0] +
                  mat_A[0][7] * mat_B[7][0] +
                  mat_A[0][8] * mat_B[8][0] +
                  mat_A[0][9] * mat_B[9][0] +
                  mat_A[0][10] * mat_B[10][0] +
                  mat_A[0][11] * mat_B[11][0] +
                  mat_A[0][12] * mat_B[12][0] +
                  mat_A[0][13] * mat_B[13][0] +
                  mat_A[0][14] * mat_B[14][0] +
                  mat_A[0][15] * mat_B[15][0] +
                  mat_A[0][16] * mat_B[16][0] +
                  mat_A[0][17] * mat_B[17][0] +
                  mat_A[0][18] * mat_B[18][0] +
                  mat_A[0][19] * mat_B[19][0] +
                  mat_A[0][20] * mat_B[20][0] +
                  mat_A[0][21] * mat_B[21][0] +
                  mat_A[0][22] * mat_B[22][0] +
                  mat_A[0][23] * mat_B[23][0] +
                  mat_A[0][24] * mat_B[24][0] +
                  mat_A[0][25] * mat_B[25][0] +
                  mat_A[0][26] * mat_B[26][0] +
                  mat_A[0][27] * mat_B[27][0] +
                  mat_A[0][28] * mat_B[28][0] +
                  mat_A[0][29] * mat_B[29][0] +
                  mat_A[0][30] * mat_B[30][0] +
                  mat_A[0][31] * mat_B[31][0];
    mat_C[0][1] <= 
                  mat_A[0][0] * mat_B[0][1] +
                  mat_A[0][1] * mat_B[1][1] +
                  mat_A[0][2] * mat_B[2][1] +
                  mat_A[0][3] * mat_B[3][1] +
                  mat_A[0][4] * mat_B[4][1] +
                  mat_A[0][5] * mat_B[5][1] +
                  mat_A[0][6] * mat_B[6][1] +
                  mat_A[0][7] * mat_B[7][1] +
                  mat_A[0][8] * mat_B[8][1] +
                  mat_A[0][9] * mat_B[9][1] +
                  mat_A[0][10] * mat_B[10][1] +
                  mat_A[0][11] * mat_B[11][1] +
                  mat_A[0][12] * mat_B[12][1] +
                  mat_A[0][13] * mat_B[13][1] +
                  mat_A[0][14] * mat_B[14][1] +
                  mat_A[0][15] * mat_B[15][1] +
                  mat_A[0][16] * mat_B[16][1] +
                  mat_A[0][17] * mat_B[17][1] +
                  mat_A[0][18] * mat_B[18][1] +
                  mat_A[0][19] * mat_B[19][1] +
                  mat_A[0][20] * mat_B[20][1] +
                  mat_A[0][21] * mat_B[21][1] +
                  mat_A[0][22] * mat_B[22][1] +
                  mat_A[0][23] * mat_B[23][1] +
                  mat_A[0][24] * mat_B[24][1] +
                  mat_A[0][25] * mat_B[25][1] +
                  mat_A[0][26] * mat_B[26][1] +
                  mat_A[0][27] * mat_B[27][1] +
                  mat_A[0][28] * mat_B[28][1] +
                  mat_A[0][29] * mat_B[29][1] +
                  mat_A[0][30] * mat_B[30][1] +
                  mat_A[0][31] * mat_B[31][1];
    mat_C[0][2] <= 
                  mat_A[0][0] * mat_B[0][2] +
                  mat_A[0][1] * mat_B[1][2] +
                  mat_A[0][2] * mat_B[2][2] +
                  mat_A[0][3] * mat_B[3][2] +
                  mat_A[0][4] * mat_B[4][2] +
                  mat_A[0][5] * mat_B[5][2] +
                  mat_A[0][6] * mat_B[6][2] +
                  mat_A[0][7] * mat_B[7][2] +
                  mat_A[0][8] * mat_B[8][2] +
                  mat_A[0][9] * mat_B[9][2] +
                  mat_A[0][10] * mat_B[10][2] +
                  mat_A[0][11] * mat_B[11][2] +
                  mat_A[0][12] * mat_B[12][2] +
                  mat_A[0][13] * mat_B[13][2] +
                  mat_A[0][14] * mat_B[14][2] +
                  mat_A[0][15] * mat_B[15][2] +
                  mat_A[0][16] * mat_B[16][2] +
                  mat_A[0][17] * mat_B[17][2] +
                  mat_A[0][18] * mat_B[18][2] +
                  mat_A[0][19] * mat_B[19][2] +
                  mat_A[0][20] * mat_B[20][2] +
                  mat_A[0][21] * mat_B[21][2] +
                  mat_A[0][22] * mat_B[22][2] +
                  mat_A[0][23] * mat_B[23][2] +
                  mat_A[0][24] * mat_B[24][2] +
                  mat_A[0][25] * mat_B[25][2] +
                  mat_A[0][26] * mat_B[26][2] +
                  mat_A[0][27] * mat_B[27][2] +
                  mat_A[0][28] * mat_B[28][2] +
                  mat_A[0][29] * mat_B[29][2] +
                  mat_A[0][30] * mat_B[30][2] +
                  mat_A[0][31] * mat_B[31][2];
    mat_C[0][3] <= 
                  mat_A[0][0] * mat_B[0][3] +
                  mat_A[0][1] * mat_B[1][3] +
                  mat_A[0][2] * mat_B[2][3] +
                  mat_A[0][3] * mat_B[3][3] +
                  mat_A[0][4] * mat_B[4][3] +
                  mat_A[0][5] * mat_B[5][3] +
                  mat_A[0][6] * mat_B[6][3] +
                  mat_A[0][7] * mat_B[7][3] +
                  mat_A[0][8] * mat_B[8][3] +
                  mat_A[0][9] * mat_B[9][3] +
                  mat_A[0][10] * mat_B[10][3] +
                  mat_A[0][11] * mat_B[11][3] +
                  mat_A[0][12] * mat_B[12][3] +
                  mat_A[0][13] * mat_B[13][3] +
                  mat_A[0][14] * mat_B[14][3] +
                  mat_A[0][15] * mat_B[15][3] +
                  mat_A[0][16] * mat_B[16][3] +
                  mat_A[0][17] * mat_B[17][3] +
                  mat_A[0][18] * mat_B[18][3] +
                  mat_A[0][19] * mat_B[19][3] +
                  mat_A[0][20] * mat_B[20][3] +
                  mat_A[0][21] * mat_B[21][3] +
                  mat_A[0][22] * mat_B[22][3] +
                  mat_A[0][23] * mat_B[23][3] +
                  mat_A[0][24] * mat_B[24][3] +
                  mat_A[0][25] * mat_B[25][3] +
                  mat_A[0][26] * mat_B[26][3] +
                  mat_A[0][27] * mat_B[27][3] +
                  mat_A[0][28] * mat_B[28][3] +
                  mat_A[0][29] * mat_B[29][3] +
                  mat_A[0][30] * mat_B[30][3] +
                  mat_A[0][31] * mat_B[31][3];
    mat_C[0][4] <= 
                  mat_A[0][0] * mat_B[0][4] +
                  mat_A[0][1] * mat_B[1][4] +
                  mat_A[0][2] * mat_B[2][4] +
                  mat_A[0][3] * mat_B[3][4] +
                  mat_A[0][4] * mat_B[4][4] +
                  mat_A[0][5] * mat_B[5][4] +
                  mat_A[0][6] * mat_B[6][4] +
                  mat_A[0][7] * mat_B[7][4] +
                  mat_A[0][8] * mat_B[8][4] +
                  mat_A[0][9] * mat_B[9][4] +
                  mat_A[0][10] * mat_B[10][4] +
                  mat_A[0][11] * mat_B[11][4] +
                  mat_A[0][12] * mat_B[12][4] +
                  mat_A[0][13] * mat_B[13][4] +
                  mat_A[0][14] * mat_B[14][4] +
                  mat_A[0][15] * mat_B[15][4] +
                  mat_A[0][16] * mat_B[16][4] +
                  mat_A[0][17] * mat_B[17][4] +
                  mat_A[0][18] * mat_B[18][4] +
                  mat_A[0][19] * mat_B[19][4] +
                  mat_A[0][20] * mat_B[20][4] +
                  mat_A[0][21] * mat_B[21][4] +
                  mat_A[0][22] * mat_B[22][4] +
                  mat_A[0][23] * mat_B[23][4] +
                  mat_A[0][24] * mat_B[24][4] +
                  mat_A[0][25] * mat_B[25][4] +
                  mat_A[0][26] * mat_B[26][4] +
                  mat_A[0][27] * mat_B[27][4] +
                  mat_A[0][28] * mat_B[28][4] +
                  mat_A[0][29] * mat_B[29][4] +
                  mat_A[0][30] * mat_B[30][4] +
                  mat_A[0][31] * mat_B[31][4];
    mat_C[0][5] <= 
                  mat_A[0][0] * mat_B[0][5] +
                  mat_A[0][1] * mat_B[1][5] +
                  mat_A[0][2] * mat_B[2][5] +
                  mat_A[0][3] * mat_B[3][5] +
                  mat_A[0][4] * mat_B[4][5] +
                  mat_A[0][5] * mat_B[5][5] +
                  mat_A[0][6] * mat_B[6][5] +
                  mat_A[0][7] * mat_B[7][5] +
                  mat_A[0][8] * mat_B[8][5] +
                  mat_A[0][9] * mat_B[9][5] +
                  mat_A[0][10] * mat_B[10][5] +
                  mat_A[0][11] * mat_B[11][5] +
                  mat_A[0][12] * mat_B[12][5] +
                  mat_A[0][13] * mat_B[13][5] +
                  mat_A[0][14] * mat_B[14][5] +
                  mat_A[0][15] * mat_B[15][5] +
                  mat_A[0][16] * mat_B[16][5] +
                  mat_A[0][17] * mat_B[17][5] +
                  mat_A[0][18] * mat_B[18][5] +
                  mat_A[0][19] * mat_B[19][5] +
                  mat_A[0][20] * mat_B[20][5] +
                  mat_A[0][21] * mat_B[21][5] +
                  mat_A[0][22] * mat_B[22][5] +
                  mat_A[0][23] * mat_B[23][5] +
                  mat_A[0][24] * mat_B[24][5] +
                  mat_A[0][25] * mat_B[25][5] +
                  mat_A[0][26] * mat_B[26][5] +
                  mat_A[0][27] * mat_B[27][5] +
                  mat_A[0][28] * mat_B[28][5] +
                  mat_A[0][29] * mat_B[29][5] +
                  mat_A[0][30] * mat_B[30][5] +
                  mat_A[0][31] * mat_B[31][5];
    mat_C[0][6] <= 
                  mat_A[0][0] * mat_B[0][6] +
                  mat_A[0][1] * mat_B[1][6] +
                  mat_A[0][2] * mat_B[2][6] +
                  mat_A[0][3] * mat_B[3][6] +
                  mat_A[0][4] * mat_B[4][6] +
                  mat_A[0][5] * mat_B[5][6] +
                  mat_A[0][6] * mat_B[6][6] +
                  mat_A[0][7] * mat_B[7][6] +
                  mat_A[0][8] * mat_B[8][6] +
                  mat_A[0][9] * mat_B[9][6] +
                  mat_A[0][10] * mat_B[10][6] +
                  mat_A[0][11] * mat_B[11][6] +
                  mat_A[0][12] * mat_B[12][6] +
                  mat_A[0][13] * mat_B[13][6] +
                  mat_A[0][14] * mat_B[14][6] +
                  mat_A[0][15] * mat_B[15][6] +
                  mat_A[0][16] * mat_B[16][6] +
                  mat_A[0][17] * mat_B[17][6] +
                  mat_A[0][18] * mat_B[18][6] +
                  mat_A[0][19] * mat_B[19][6] +
                  mat_A[0][20] * mat_B[20][6] +
                  mat_A[0][21] * mat_B[21][6] +
                  mat_A[0][22] * mat_B[22][6] +
                  mat_A[0][23] * mat_B[23][6] +
                  mat_A[0][24] * mat_B[24][6] +
                  mat_A[0][25] * mat_B[25][6] +
                  mat_A[0][26] * mat_B[26][6] +
                  mat_A[0][27] * mat_B[27][6] +
                  mat_A[0][28] * mat_B[28][6] +
                  mat_A[0][29] * mat_B[29][6] +
                  mat_A[0][30] * mat_B[30][6] +
                  mat_A[0][31] * mat_B[31][6];
    mat_C[0][7] <= 
                  mat_A[0][0] * mat_B[0][7] +
                  mat_A[0][1] * mat_B[1][7] +
                  mat_A[0][2] * mat_B[2][7] +
                  mat_A[0][3] * mat_B[3][7] +
                  mat_A[0][4] * mat_B[4][7] +
                  mat_A[0][5] * mat_B[5][7] +
                  mat_A[0][6] * mat_B[6][7] +
                  mat_A[0][7] * mat_B[7][7] +
                  mat_A[0][8] * mat_B[8][7] +
                  mat_A[0][9] * mat_B[9][7] +
                  mat_A[0][10] * mat_B[10][7] +
                  mat_A[0][11] * mat_B[11][7] +
                  mat_A[0][12] * mat_B[12][7] +
                  mat_A[0][13] * mat_B[13][7] +
                  mat_A[0][14] * mat_B[14][7] +
                  mat_A[0][15] * mat_B[15][7] +
                  mat_A[0][16] * mat_B[16][7] +
                  mat_A[0][17] * mat_B[17][7] +
                  mat_A[0][18] * mat_B[18][7] +
                  mat_A[0][19] * mat_B[19][7] +
                  mat_A[0][20] * mat_B[20][7] +
                  mat_A[0][21] * mat_B[21][7] +
                  mat_A[0][22] * mat_B[22][7] +
                  mat_A[0][23] * mat_B[23][7] +
                  mat_A[0][24] * mat_B[24][7] +
                  mat_A[0][25] * mat_B[25][7] +
                  mat_A[0][26] * mat_B[26][7] +
                  mat_A[0][27] * mat_B[27][7] +
                  mat_A[0][28] * mat_B[28][7] +
                  mat_A[0][29] * mat_B[29][7] +
                  mat_A[0][30] * mat_B[30][7] +
                  mat_A[0][31] * mat_B[31][7];
    mat_C[0][8] <= 
                  mat_A[0][0] * mat_B[0][8] +
                  mat_A[0][1] * mat_B[1][8] +
                  mat_A[0][2] * mat_B[2][8] +
                  mat_A[0][3] * mat_B[3][8] +
                  mat_A[0][4] * mat_B[4][8] +
                  mat_A[0][5] * mat_B[5][8] +
                  mat_A[0][6] * mat_B[6][8] +
                  mat_A[0][7] * mat_B[7][8] +
                  mat_A[0][8] * mat_B[8][8] +
                  mat_A[0][9] * mat_B[9][8] +
                  mat_A[0][10] * mat_B[10][8] +
                  mat_A[0][11] * mat_B[11][8] +
                  mat_A[0][12] * mat_B[12][8] +
                  mat_A[0][13] * mat_B[13][8] +
                  mat_A[0][14] * mat_B[14][8] +
                  mat_A[0][15] * mat_B[15][8] +
                  mat_A[0][16] * mat_B[16][8] +
                  mat_A[0][17] * mat_B[17][8] +
                  mat_A[0][18] * mat_B[18][8] +
                  mat_A[0][19] * mat_B[19][8] +
                  mat_A[0][20] * mat_B[20][8] +
                  mat_A[0][21] * mat_B[21][8] +
                  mat_A[0][22] * mat_B[22][8] +
                  mat_A[0][23] * mat_B[23][8] +
                  mat_A[0][24] * mat_B[24][8] +
                  mat_A[0][25] * mat_B[25][8] +
                  mat_A[0][26] * mat_B[26][8] +
                  mat_A[0][27] * mat_B[27][8] +
                  mat_A[0][28] * mat_B[28][8] +
                  mat_A[0][29] * mat_B[29][8] +
                  mat_A[0][30] * mat_B[30][8] +
                  mat_A[0][31] * mat_B[31][8];
    mat_C[0][9] <= 
                  mat_A[0][0] * mat_B[0][9] +
                  mat_A[0][1] * mat_B[1][9] +
                  mat_A[0][2] * mat_B[2][9] +
                  mat_A[0][3] * mat_B[3][9] +
                  mat_A[0][4] * mat_B[4][9] +
                  mat_A[0][5] * mat_B[5][9] +
                  mat_A[0][6] * mat_B[6][9] +
                  mat_A[0][7] * mat_B[7][9] +
                  mat_A[0][8] * mat_B[8][9] +
                  mat_A[0][9] * mat_B[9][9] +
                  mat_A[0][10] * mat_B[10][9] +
                  mat_A[0][11] * mat_B[11][9] +
                  mat_A[0][12] * mat_B[12][9] +
                  mat_A[0][13] * mat_B[13][9] +
                  mat_A[0][14] * mat_B[14][9] +
                  mat_A[0][15] * mat_B[15][9] +
                  mat_A[0][16] * mat_B[16][9] +
                  mat_A[0][17] * mat_B[17][9] +
                  mat_A[0][18] * mat_B[18][9] +
                  mat_A[0][19] * mat_B[19][9] +
                  mat_A[0][20] * mat_B[20][9] +
                  mat_A[0][21] * mat_B[21][9] +
                  mat_A[0][22] * mat_B[22][9] +
                  mat_A[0][23] * mat_B[23][9] +
                  mat_A[0][24] * mat_B[24][9] +
                  mat_A[0][25] * mat_B[25][9] +
                  mat_A[0][26] * mat_B[26][9] +
                  mat_A[0][27] * mat_B[27][9] +
                  mat_A[0][28] * mat_B[28][9] +
                  mat_A[0][29] * mat_B[29][9] +
                  mat_A[0][30] * mat_B[30][9] +
                  mat_A[0][31] * mat_B[31][9];
    mat_C[0][10] <= 
                  mat_A[0][0] * mat_B[0][10] +
                  mat_A[0][1] * mat_B[1][10] +
                  mat_A[0][2] * mat_B[2][10] +
                  mat_A[0][3] * mat_B[3][10] +
                  mat_A[0][4] * mat_B[4][10] +
                  mat_A[0][5] * mat_B[5][10] +
                  mat_A[0][6] * mat_B[6][10] +
                  mat_A[0][7] * mat_B[7][10] +
                  mat_A[0][8] * mat_B[8][10] +
                  mat_A[0][9] * mat_B[9][10] +
                  mat_A[0][10] * mat_B[10][10] +
                  mat_A[0][11] * mat_B[11][10] +
                  mat_A[0][12] * mat_B[12][10] +
                  mat_A[0][13] * mat_B[13][10] +
                  mat_A[0][14] * mat_B[14][10] +
                  mat_A[0][15] * mat_B[15][10] +
                  mat_A[0][16] * mat_B[16][10] +
                  mat_A[0][17] * mat_B[17][10] +
                  mat_A[0][18] * mat_B[18][10] +
                  mat_A[0][19] * mat_B[19][10] +
                  mat_A[0][20] * mat_B[20][10] +
                  mat_A[0][21] * mat_B[21][10] +
                  mat_A[0][22] * mat_B[22][10] +
                  mat_A[0][23] * mat_B[23][10] +
                  mat_A[0][24] * mat_B[24][10] +
                  mat_A[0][25] * mat_B[25][10] +
                  mat_A[0][26] * mat_B[26][10] +
                  mat_A[0][27] * mat_B[27][10] +
                  mat_A[0][28] * mat_B[28][10] +
                  mat_A[0][29] * mat_B[29][10] +
                  mat_A[0][30] * mat_B[30][10] +
                  mat_A[0][31] * mat_B[31][10];
    mat_C[0][11] <= 
                  mat_A[0][0] * mat_B[0][11] +
                  mat_A[0][1] * mat_B[1][11] +
                  mat_A[0][2] * mat_B[2][11] +
                  mat_A[0][3] * mat_B[3][11] +
                  mat_A[0][4] * mat_B[4][11] +
                  mat_A[0][5] * mat_B[5][11] +
                  mat_A[0][6] * mat_B[6][11] +
                  mat_A[0][7] * mat_B[7][11] +
                  mat_A[0][8] * mat_B[8][11] +
                  mat_A[0][9] * mat_B[9][11] +
                  mat_A[0][10] * mat_B[10][11] +
                  mat_A[0][11] * mat_B[11][11] +
                  mat_A[0][12] * mat_B[12][11] +
                  mat_A[0][13] * mat_B[13][11] +
                  mat_A[0][14] * mat_B[14][11] +
                  mat_A[0][15] * mat_B[15][11] +
                  mat_A[0][16] * mat_B[16][11] +
                  mat_A[0][17] * mat_B[17][11] +
                  mat_A[0][18] * mat_B[18][11] +
                  mat_A[0][19] * mat_B[19][11] +
                  mat_A[0][20] * mat_B[20][11] +
                  mat_A[0][21] * mat_B[21][11] +
                  mat_A[0][22] * mat_B[22][11] +
                  mat_A[0][23] * mat_B[23][11] +
                  mat_A[0][24] * mat_B[24][11] +
                  mat_A[0][25] * mat_B[25][11] +
                  mat_A[0][26] * mat_B[26][11] +
                  mat_A[0][27] * mat_B[27][11] +
                  mat_A[0][28] * mat_B[28][11] +
                  mat_A[0][29] * mat_B[29][11] +
                  mat_A[0][30] * mat_B[30][11] +
                  mat_A[0][31] * mat_B[31][11];
    mat_C[0][12] <= 
                  mat_A[0][0] * mat_B[0][12] +
                  mat_A[0][1] * mat_B[1][12] +
                  mat_A[0][2] * mat_B[2][12] +
                  mat_A[0][3] * mat_B[3][12] +
                  mat_A[0][4] * mat_B[4][12] +
                  mat_A[0][5] * mat_B[5][12] +
                  mat_A[0][6] * mat_B[6][12] +
                  mat_A[0][7] * mat_B[7][12] +
                  mat_A[0][8] * mat_B[8][12] +
                  mat_A[0][9] * mat_B[9][12] +
                  mat_A[0][10] * mat_B[10][12] +
                  mat_A[0][11] * mat_B[11][12] +
                  mat_A[0][12] * mat_B[12][12] +
                  mat_A[0][13] * mat_B[13][12] +
                  mat_A[0][14] * mat_B[14][12] +
                  mat_A[0][15] * mat_B[15][12] +
                  mat_A[0][16] * mat_B[16][12] +
                  mat_A[0][17] * mat_B[17][12] +
                  mat_A[0][18] * mat_B[18][12] +
                  mat_A[0][19] * mat_B[19][12] +
                  mat_A[0][20] * mat_B[20][12] +
                  mat_A[0][21] * mat_B[21][12] +
                  mat_A[0][22] * mat_B[22][12] +
                  mat_A[0][23] * mat_B[23][12] +
                  mat_A[0][24] * mat_B[24][12] +
                  mat_A[0][25] * mat_B[25][12] +
                  mat_A[0][26] * mat_B[26][12] +
                  mat_A[0][27] * mat_B[27][12] +
                  mat_A[0][28] * mat_B[28][12] +
                  mat_A[0][29] * mat_B[29][12] +
                  mat_A[0][30] * mat_B[30][12] +
                  mat_A[0][31] * mat_B[31][12];
    mat_C[0][13] <= 
                  mat_A[0][0] * mat_B[0][13] +
                  mat_A[0][1] * mat_B[1][13] +
                  mat_A[0][2] * mat_B[2][13] +
                  mat_A[0][3] * mat_B[3][13] +
                  mat_A[0][4] * mat_B[4][13] +
                  mat_A[0][5] * mat_B[5][13] +
                  mat_A[0][6] * mat_B[6][13] +
                  mat_A[0][7] * mat_B[7][13] +
                  mat_A[0][8] * mat_B[8][13] +
                  mat_A[0][9] * mat_B[9][13] +
                  mat_A[0][10] * mat_B[10][13] +
                  mat_A[0][11] * mat_B[11][13] +
                  mat_A[0][12] * mat_B[12][13] +
                  mat_A[0][13] * mat_B[13][13] +
                  mat_A[0][14] * mat_B[14][13] +
                  mat_A[0][15] * mat_B[15][13] +
                  mat_A[0][16] * mat_B[16][13] +
                  mat_A[0][17] * mat_B[17][13] +
                  mat_A[0][18] * mat_B[18][13] +
                  mat_A[0][19] * mat_B[19][13] +
                  mat_A[0][20] * mat_B[20][13] +
                  mat_A[0][21] * mat_B[21][13] +
                  mat_A[0][22] * mat_B[22][13] +
                  mat_A[0][23] * mat_B[23][13] +
                  mat_A[0][24] * mat_B[24][13] +
                  mat_A[0][25] * mat_B[25][13] +
                  mat_A[0][26] * mat_B[26][13] +
                  mat_A[0][27] * mat_B[27][13] +
                  mat_A[0][28] * mat_B[28][13] +
                  mat_A[0][29] * mat_B[29][13] +
                  mat_A[0][30] * mat_B[30][13] +
                  mat_A[0][31] * mat_B[31][13];
    mat_C[0][14] <= 
                  mat_A[0][0] * mat_B[0][14] +
                  mat_A[0][1] * mat_B[1][14] +
                  mat_A[0][2] * mat_B[2][14] +
                  mat_A[0][3] * mat_B[3][14] +
                  mat_A[0][4] * mat_B[4][14] +
                  mat_A[0][5] * mat_B[5][14] +
                  mat_A[0][6] * mat_B[6][14] +
                  mat_A[0][7] * mat_B[7][14] +
                  mat_A[0][8] * mat_B[8][14] +
                  mat_A[0][9] * mat_B[9][14] +
                  mat_A[0][10] * mat_B[10][14] +
                  mat_A[0][11] * mat_B[11][14] +
                  mat_A[0][12] * mat_B[12][14] +
                  mat_A[0][13] * mat_B[13][14] +
                  mat_A[0][14] * mat_B[14][14] +
                  mat_A[0][15] * mat_B[15][14] +
                  mat_A[0][16] * mat_B[16][14] +
                  mat_A[0][17] * mat_B[17][14] +
                  mat_A[0][18] * mat_B[18][14] +
                  mat_A[0][19] * mat_B[19][14] +
                  mat_A[0][20] * mat_B[20][14] +
                  mat_A[0][21] * mat_B[21][14] +
                  mat_A[0][22] * mat_B[22][14] +
                  mat_A[0][23] * mat_B[23][14] +
                  mat_A[0][24] * mat_B[24][14] +
                  mat_A[0][25] * mat_B[25][14] +
                  mat_A[0][26] * mat_B[26][14] +
                  mat_A[0][27] * mat_B[27][14] +
                  mat_A[0][28] * mat_B[28][14] +
                  mat_A[0][29] * mat_B[29][14] +
                  mat_A[0][30] * mat_B[30][14] +
                  mat_A[0][31] * mat_B[31][14];
    mat_C[0][15] <= 
                  mat_A[0][0] * mat_B[0][15] +
                  mat_A[0][1] * mat_B[1][15] +
                  mat_A[0][2] * mat_B[2][15] +
                  mat_A[0][3] * mat_B[3][15] +
                  mat_A[0][4] * mat_B[4][15] +
                  mat_A[0][5] * mat_B[5][15] +
                  mat_A[0][6] * mat_B[6][15] +
                  mat_A[0][7] * mat_B[7][15] +
                  mat_A[0][8] * mat_B[8][15] +
                  mat_A[0][9] * mat_B[9][15] +
                  mat_A[0][10] * mat_B[10][15] +
                  mat_A[0][11] * mat_B[11][15] +
                  mat_A[0][12] * mat_B[12][15] +
                  mat_A[0][13] * mat_B[13][15] +
                  mat_A[0][14] * mat_B[14][15] +
                  mat_A[0][15] * mat_B[15][15] +
                  mat_A[0][16] * mat_B[16][15] +
                  mat_A[0][17] * mat_B[17][15] +
                  mat_A[0][18] * mat_B[18][15] +
                  mat_A[0][19] * mat_B[19][15] +
                  mat_A[0][20] * mat_B[20][15] +
                  mat_A[0][21] * mat_B[21][15] +
                  mat_A[0][22] * mat_B[22][15] +
                  mat_A[0][23] * mat_B[23][15] +
                  mat_A[0][24] * mat_B[24][15] +
                  mat_A[0][25] * mat_B[25][15] +
                  mat_A[0][26] * mat_B[26][15] +
                  mat_A[0][27] * mat_B[27][15] +
                  mat_A[0][28] * mat_B[28][15] +
                  mat_A[0][29] * mat_B[29][15] +
                  mat_A[0][30] * mat_B[30][15] +
                  mat_A[0][31] * mat_B[31][15];
    mat_C[0][16] <= 
                  mat_A[0][0] * mat_B[0][16] +
                  mat_A[0][1] * mat_B[1][16] +
                  mat_A[0][2] * mat_B[2][16] +
                  mat_A[0][3] * mat_B[3][16] +
                  mat_A[0][4] * mat_B[4][16] +
                  mat_A[0][5] * mat_B[5][16] +
                  mat_A[0][6] * mat_B[6][16] +
                  mat_A[0][7] * mat_B[7][16] +
                  mat_A[0][8] * mat_B[8][16] +
                  mat_A[0][9] * mat_B[9][16] +
                  mat_A[0][10] * mat_B[10][16] +
                  mat_A[0][11] * mat_B[11][16] +
                  mat_A[0][12] * mat_B[12][16] +
                  mat_A[0][13] * mat_B[13][16] +
                  mat_A[0][14] * mat_B[14][16] +
                  mat_A[0][15] * mat_B[15][16] +
                  mat_A[0][16] * mat_B[16][16] +
                  mat_A[0][17] * mat_B[17][16] +
                  mat_A[0][18] * mat_B[18][16] +
                  mat_A[0][19] * mat_B[19][16] +
                  mat_A[0][20] * mat_B[20][16] +
                  mat_A[0][21] * mat_B[21][16] +
                  mat_A[0][22] * mat_B[22][16] +
                  mat_A[0][23] * mat_B[23][16] +
                  mat_A[0][24] * mat_B[24][16] +
                  mat_A[0][25] * mat_B[25][16] +
                  mat_A[0][26] * mat_B[26][16] +
                  mat_A[0][27] * mat_B[27][16] +
                  mat_A[0][28] * mat_B[28][16] +
                  mat_A[0][29] * mat_B[29][16] +
                  mat_A[0][30] * mat_B[30][16] +
                  mat_A[0][31] * mat_B[31][16];
    mat_C[0][17] <= 
                  mat_A[0][0] * mat_B[0][17] +
                  mat_A[0][1] * mat_B[1][17] +
                  mat_A[0][2] * mat_B[2][17] +
                  mat_A[0][3] * mat_B[3][17] +
                  mat_A[0][4] * mat_B[4][17] +
                  mat_A[0][5] * mat_B[5][17] +
                  mat_A[0][6] * mat_B[6][17] +
                  mat_A[0][7] * mat_B[7][17] +
                  mat_A[0][8] * mat_B[8][17] +
                  mat_A[0][9] * mat_B[9][17] +
                  mat_A[0][10] * mat_B[10][17] +
                  mat_A[0][11] * mat_B[11][17] +
                  mat_A[0][12] * mat_B[12][17] +
                  mat_A[0][13] * mat_B[13][17] +
                  mat_A[0][14] * mat_B[14][17] +
                  mat_A[0][15] * mat_B[15][17] +
                  mat_A[0][16] * mat_B[16][17] +
                  mat_A[0][17] * mat_B[17][17] +
                  mat_A[0][18] * mat_B[18][17] +
                  mat_A[0][19] * mat_B[19][17] +
                  mat_A[0][20] * mat_B[20][17] +
                  mat_A[0][21] * mat_B[21][17] +
                  mat_A[0][22] * mat_B[22][17] +
                  mat_A[0][23] * mat_B[23][17] +
                  mat_A[0][24] * mat_B[24][17] +
                  mat_A[0][25] * mat_B[25][17] +
                  mat_A[0][26] * mat_B[26][17] +
                  mat_A[0][27] * mat_B[27][17] +
                  mat_A[0][28] * mat_B[28][17] +
                  mat_A[0][29] * mat_B[29][17] +
                  mat_A[0][30] * mat_B[30][17] +
                  mat_A[0][31] * mat_B[31][17];
    mat_C[0][18] <= 
                  mat_A[0][0] * mat_B[0][18] +
                  mat_A[0][1] * mat_B[1][18] +
                  mat_A[0][2] * mat_B[2][18] +
                  mat_A[0][3] * mat_B[3][18] +
                  mat_A[0][4] * mat_B[4][18] +
                  mat_A[0][5] * mat_B[5][18] +
                  mat_A[0][6] * mat_B[6][18] +
                  mat_A[0][7] * mat_B[7][18] +
                  mat_A[0][8] * mat_B[8][18] +
                  mat_A[0][9] * mat_B[9][18] +
                  mat_A[0][10] * mat_B[10][18] +
                  mat_A[0][11] * mat_B[11][18] +
                  mat_A[0][12] * mat_B[12][18] +
                  mat_A[0][13] * mat_B[13][18] +
                  mat_A[0][14] * mat_B[14][18] +
                  mat_A[0][15] * mat_B[15][18] +
                  mat_A[0][16] * mat_B[16][18] +
                  mat_A[0][17] * mat_B[17][18] +
                  mat_A[0][18] * mat_B[18][18] +
                  mat_A[0][19] * mat_B[19][18] +
                  mat_A[0][20] * mat_B[20][18] +
                  mat_A[0][21] * mat_B[21][18] +
                  mat_A[0][22] * mat_B[22][18] +
                  mat_A[0][23] * mat_B[23][18] +
                  mat_A[0][24] * mat_B[24][18] +
                  mat_A[0][25] * mat_B[25][18] +
                  mat_A[0][26] * mat_B[26][18] +
                  mat_A[0][27] * mat_B[27][18] +
                  mat_A[0][28] * mat_B[28][18] +
                  mat_A[0][29] * mat_B[29][18] +
                  mat_A[0][30] * mat_B[30][18] +
                  mat_A[0][31] * mat_B[31][18];
    mat_C[0][19] <= 
                  mat_A[0][0] * mat_B[0][19] +
                  mat_A[0][1] * mat_B[1][19] +
                  mat_A[0][2] * mat_B[2][19] +
                  mat_A[0][3] * mat_B[3][19] +
                  mat_A[0][4] * mat_B[4][19] +
                  mat_A[0][5] * mat_B[5][19] +
                  mat_A[0][6] * mat_B[6][19] +
                  mat_A[0][7] * mat_B[7][19] +
                  mat_A[0][8] * mat_B[8][19] +
                  mat_A[0][9] * mat_B[9][19] +
                  mat_A[0][10] * mat_B[10][19] +
                  mat_A[0][11] * mat_B[11][19] +
                  mat_A[0][12] * mat_B[12][19] +
                  mat_A[0][13] * mat_B[13][19] +
                  mat_A[0][14] * mat_B[14][19] +
                  mat_A[0][15] * mat_B[15][19] +
                  mat_A[0][16] * mat_B[16][19] +
                  mat_A[0][17] * mat_B[17][19] +
                  mat_A[0][18] * mat_B[18][19] +
                  mat_A[0][19] * mat_B[19][19] +
                  mat_A[0][20] * mat_B[20][19] +
                  mat_A[0][21] * mat_B[21][19] +
                  mat_A[0][22] * mat_B[22][19] +
                  mat_A[0][23] * mat_B[23][19] +
                  mat_A[0][24] * mat_B[24][19] +
                  mat_A[0][25] * mat_B[25][19] +
                  mat_A[0][26] * mat_B[26][19] +
                  mat_A[0][27] * mat_B[27][19] +
                  mat_A[0][28] * mat_B[28][19] +
                  mat_A[0][29] * mat_B[29][19] +
                  mat_A[0][30] * mat_B[30][19] +
                  mat_A[0][31] * mat_B[31][19];
    mat_C[0][20] <= 
                  mat_A[0][0] * mat_B[0][20] +
                  mat_A[0][1] * mat_B[1][20] +
                  mat_A[0][2] * mat_B[2][20] +
                  mat_A[0][3] * mat_B[3][20] +
                  mat_A[0][4] * mat_B[4][20] +
                  mat_A[0][5] * mat_B[5][20] +
                  mat_A[0][6] * mat_B[6][20] +
                  mat_A[0][7] * mat_B[7][20] +
                  mat_A[0][8] * mat_B[8][20] +
                  mat_A[0][9] * mat_B[9][20] +
                  mat_A[0][10] * mat_B[10][20] +
                  mat_A[0][11] * mat_B[11][20] +
                  mat_A[0][12] * mat_B[12][20] +
                  mat_A[0][13] * mat_B[13][20] +
                  mat_A[0][14] * mat_B[14][20] +
                  mat_A[0][15] * mat_B[15][20] +
                  mat_A[0][16] * mat_B[16][20] +
                  mat_A[0][17] * mat_B[17][20] +
                  mat_A[0][18] * mat_B[18][20] +
                  mat_A[0][19] * mat_B[19][20] +
                  mat_A[0][20] * mat_B[20][20] +
                  mat_A[0][21] * mat_B[21][20] +
                  mat_A[0][22] * mat_B[22][20] +
                  mat_A[0][23] * mat_B[23][20] +
                  mat_A[0][24] * mat_B[24][20] +
                  mat_A[0][25] * mat_B[25][20] +
                  mat_A[0][26] * mat_B[26][20] +
                  mat_A[0][27] * mat_B[27][20] +
                  mat_A[0][28] * mat_B[28][20] +
                  mat_A[0][29] * mat_B[29][20] +
                  mat_A[0][30] * mat_B[30][20] +
                  mat_A[0][31] * mat_B[31][20];
    mat_C[0][21] <= 
                  mat_A[0][0] * mat_B[0][21] +
                  mat_A[0][1] * mat_B[1][21] +
                  mat_A[0][2] * mat_B[2][21] +
                  mat_A[0][3] * mat_B[3][21] +
                  mat_A[0][4] * mat_B[4][21] +
                  mat_A[0][5] * mat_B[5][21] +
                  mat_A[0][6] * mat_B[6][21] +
                  mat_A[0][7] * mat_B[7][21] +
                  mat_A[0][8] * mat_B[8][21] +
                  mat_A[0][9] * mat_B[9][21] +
                  mat_A[0][10] * mat_B[10][21] +
                  mat_A[0][11] * mat_B[11][21] +
                  mat_A[0][12] * mat_B[12][21] +
                  mat_A[0][13] * mat_B[13][21] +
                  mat_A[0][14] * mat_B[14][21] +
                  mat_A[0][15] * mat_B[15][21] +
                  mat_A[0][16] * mat_B[16][21] +
                  mat_A[0][17] * mat_B[17][21] +
                  mat_A[0][18] * mat_B[18][21] +
                  mat_A[0][19] * mat_B[19][21] +
                  mat_A[0][20] * mat_B[20][21] +
                  mat_A[0][21] * mat_B[21][21] +
                  mat_A[0][22] * mat_B[22][21] +
                  mat_A[0][23] * mat_B[23][21] +
                  mat_A[0][24] * mat_B[24][21] +
                  mat_A[0][25] * mat_B[25][21] +
                  mat_A[0][26] * mat_B[26][21] +
                  mat_A[0][27] * mat_B[27][21] +
                  mat_A[0][28] * mat_B[28][21] +
                  mat_A[0][29] * mat_B[29][21] +
                  mat_A[0][30] * mat_B[30][21] +
                  mat_A[0][31] * mat_B[31][21];
    mat_C[0][22] <= 
                  mat_A[0][0] * mat_B[0][22] +
                  mat_A[0][1] * mat_B[1][22] +
                  mat_A[0][2] * mat_B[2][22] +
                  mat_A[0][3] * mat_B[3][22] +
                  mat_A[0][4] * mat_B[4][22] +
                  mat_A[0][5] * mat_B[5][22] +
                  mat_A[0][6] * mat_B[6][22] +
                  mat_A[0][7] * mat_B[7][22] +
                  mat_A[0][8] * mat_B[8][22] +
                  mat_A[0][9] * mat_B[9][22] +
                  mat_A[0][10] * mat_B[10][22] +
                  mat_A[0][11] * mat_B[11][22] +
                  mat_A[0][12] * mat_B[12][22] +
                  mat_A[0][13] * mat_B[13][22] +
                  mat_A[0][14] * mat_B[14][22] +
                  mat_A[0][15] * mat_B[15][22] +
                  mat_A[0][16] * mat_B[16][22] +
                  mat_A[0][17] * mat_B[17][22] +
                  mat_A[0][18] * mat_B[18][22] +
                  mat_A[0][19] * mat_B[19][22] +
                  mat_A[0][20] * mat_B[20][22] +
                  mat_A[0][21] * mat_B[21][22] +
                  mat_A[0][22] * mat_B[22][22] +
                  mat_A[0][23] * mat_B[23][22] +
                  mat_A[0][24] * mat_B[24][22] +
                  mat_A[0][25] * mat_B[25][22] +
                  mat_A[0][26] * mat_B[26][22] +
                  mat_A[0][27] * mat_B[27][22] +
                  mat_A[0][28] * mat_B[28][22] +
                  mat_A[0][29] * mat_B[29][22] +
                  mat_A[0][30] * mat_B[30][22] +
                  mat_A[0][31] * mat_B[31][22];
    mat_C[0][23] <= 
                  mat_A[0][0] * mat_B[0][23] +
                  mat_A[0][1] * mat_B[1][23] +
                  mat_A[0][2] * mat_B[2][23] +
                  mat_A[0][3] * mat_B[3][23] +
                  mat_A[0][4] * mat_B[4][23] +
                  mat_A[0][5] * mat_B[5][23] +
                  mat_A[0][6] * mat_B[6][23] +
                  mat_A[0][7] * mat_B[7][23] +
                  mat_A[0][8] * mat_B[8][23] +
                  mat_A[0][9] * mat_B[9][23] +
                  mat_A[0][10] * mat_B[10][23] +
                  mat_A[0][11] * mat_B[11][23] +
                  mat_A[0][12] * mat_B[12][23] +
                  mat_A[0][13] * mat_B[13][23] +
                  mat_A[0][14] * mat_B[14][23] +
                  mat_A[0][15] * mat_B[15][23] +
                  mat_A[0][16] * mat_B[16][23] +
                  mat_A[0][17] * mat_B[17][23] +
                  mat_A[0][18] * mat_B[18][23] +
                  mat_A[0][19] * mat_B[19][23] +
                  mat_A[0][20] * mat_B[20][23] +
                  mat_A[0][21] * mat_B[21][23] +
                  mat_A[0][22] * mat_B[22][23] +
                  mat_A[0][23] * mat_B[23][23] +
                  mat_A[0][24] * mat_B[24][23] +
                  mat_A[0][25] * mat_B[25][23] +
                  mat_A[0][26] * mat_B[26][23] +
                  mat_A[0][27] * mat_B[27][23] +
                  mat_A[0][28] * mat_B[28][23] +
                  mat_A[0][29] * mat_B[29][23] +
                  mat_A[0][30] * mat_B[30][23] +
                  mat_A[0][31] * mat_B[31][23];
    mat_C[0][24] <= 
                  mat_A[0][0] * mat_B[0][24] +
                  mat_A[0][1] * mat_B[1][24] +
                  mat_A[0][2] * mat_B[2][24] +
                  mat_A[0][3] * mat_B[3][24] +
                  mat_A[0][4] * mat_B[4][24] +
                  mat_A[0][5] * mat_B[5][24] +
                  mat_A[0][6] * mat_B[6][24] +
                  mat_A[0][7] * mat_B[7][24] +
                  mat_A[0][8] * mat_B[8][24] +
                  mat_A[0][9] * mat_B[9][24] +
                  mat_A[0][10] * mat_B[10][24] +
                  mat_A[0][11] * mat_B[11][24] +
                  mat_A[0][12] * mat_B[12][24] +
                  mat_A[0][13] * mat_B[13][24] +
                  mat_A[0][14] * mat_B[14][24] +
                  mat_A[0][15] * mat_B[15][24] +
                  mat_A[0][16] * mat_B[16][24] +
                  mat_A[0][17] * mat_B[17][24] +
                  mat_A[0][18] * mat_B[18][24] +
                  mat_A[0][19] * mat_B[19][24] +
                  mat_A[0][20] * mat_B[20][24] +
                  mat_A[0][21] * mat_B[21][24] +
                  mat_A[0][22] * mat_B[22][24] +
                  mat_A[0][23] * mat_B[23][24] +
                  mat_A[0][24] * mat_B[24][24] +
                  mat_A[0][25] * mat_B[25][24] +
                  mat_A[0][26] * mat_B[26][24] +
                  mat_A[0][27] * mat_B[27][24] +
                  mat_A[0][28] * mat_B[28][24] +
                  mat_A[0][29] * mat_B[29][24] +
                  mat_A[0][30] * mat_B[30][24] +
                  mat_A[0][31] * mat_B[31][24];
    mat_C[0][25] <= 
                  mat_A[0][0] * mat_B[0][25] +
                  mat_A[0][1] * mat_B[1][25] +
                  mat_A[0][2] * mat_B[2][25] +
                  mat_A[0][3] * mat_B[3][25] +
                  mat_A[0][4] * mat_B[4][25] +
                  mat_A[0][5] * mat_B[5][25] +
                  mat_A[0][6] * mat_B[6][25] +
                  mat_A[0][7] * mat_B[7][25] +
                  mat_A[0][8] * mat_B[8][25] +
                  mat_A[0][9] * mat_B[9][25] +
                  mat_A[0][10] * mat_B[10][25] +
                  mat_A[0][11] * mat_B[11][25] +
                  mat_A[0][12] * mat_B[12][25] +
                  mat_A[0][13] * mat_B[13][25] +
                  mat_A[0][14] * mat_B[14][25] +
                  mat_A[0][15] * mat_B[15][25] +
                  mat_A[0][16] * mat_B[16][25] +
                  mat_A[0][17] * mat_B[17][25] +
                  mat_A[0][18] * mat_B[18][25] +
                  mat_A[0][19] * mat_B[19][25] +
                  mat_A[0][20] * mat_B[20][25] +
                  mat_A[0][21] * mat_B[21][25] +
                  mat_A[0][22] * mat_B[22][25] +
                  mat_A[0][23] * mat_B[23][25] +
                  mat_A[0][24] * mat_B[24][25] +
                  mat_A[0][25] * mat_B[25][25] +
                  mat_A[0][26] * mat_B[26][25] +
                  mat_A[0][27] * mat_B[27][25] +
                  mat_A[0][28] * mat_B[28][25] +
                  mat_A[0][29] * mat_B[29][25] +
                  mat_A[0][30] * mat_B[30][25] +
                  mat_A[0][31] * mat_B[31][25];
    mat_C[0][26] <= 
                  mat_A[0][0] * mat_B[0][26] +
                  mat_A[0][1] * mat_B[1][26] +
                  mat_A[0][2] * mat_B[2][26] +
                  mat_A[0][3] * mat_B[3][26] +
                  mat_A[0][4] * mat_B[4][26] +
                  mat_A[0][5] * mat_B[5][26] +
                  mat_A[0][6] * mat_B[6][26] +
                  mat_A[0][7] * mat_B[7][26] +
                  mat_A[0][8] * mat_B[8][26] +
                  mat_A[0][9] * mat_B[9][26] +
                  mat_A[0][10] * mat_B[10][26] +
                  mat_A[0][11] * mat_B[11][26] +
                  mat_A[0][12] * mat_B[12][26] +
                  mat_A[0][13] * mat_B[13][26] +
                  mat_A[0][14] * mat_B[14][26] +
                  mat_A[0][15] * mat_B[15][26] +
                  mat_A[0][16] * mat_B[16][26] +
                  mat_A[0][17] * mat_B[17][26] +
                  mat_A[0][18] * mat_B[18][26] +
                  mat_A[0][19] * mat_B[19][26] +
                  mat_A[0][20] * mat_B[20][26] +
                  mat_A[0][21] * mat_B[21][26] +
                  mat_A[0][22] * mat_B[22][26] +
                  mat_A[0][23] * mat_B[23][26] +
                  mat_A[0][24] * mat_B[24][26] +
                  mat_A[0][25] * mat_B[25][26] +
                  mat_A[0][26] * mat_B[26][26] +
                  mat_A[0][27] * mat_B[27][26] +
                  mat_A[0][28] * mat_B[28][26] +
                  mat_A[0][29] * mat_B[29][26] +
                  mat_A[0][30] * mat_B[30][26] +
                  mat_A[0][31] * mat_B[31][26];
    mat_C[0][27] <= 
                  mat_A[0][0] * mat_B[0][27] +
                  mat_A[0][1] * mat_B[1][27] +
                  mat_A[0][2] * mat_B[2][27] +
                  mat_A[0][3] * mat_B[3][27] +
                  mat_A[0][4] * mat_B[4][27] +
                  mat_A[0][5] * mat_B[5][27] +
                  mat_A[0][6] * mat_B[6][27] +
                  mat_A[0][7] * mat_B[7][27] +
                  mat_A[0][8] * mat_B[8][27] +
                  mat_A[0][9] * mat_B[9][27] +
                  mat_A[0][10] * mat_B[10][27] +
                  mat_A[0][11] * mat_B[11][27] +
                  mat_A[0][12] * mat_B[12][27] +
                  mat_A[0][13] * mat_B[13][27] +
                  mat_A[0][14] * mat_B[14][27] +
                  mat_A[0][15] * mat_B[15][27] +
                  mat_A[0][16] * mat_B[16][27] +
                  mat_A[0][17] * mat_B[17][27] +
                  mat_A[0][18] * mat_B[18][27] +
                  mat_A[0][19] * mat_B[19][27] +
                  mat_A[0][20] * mat_B[20][27] +
                  mat_A[0][21] * mat_B[21][27] +
                  mat_A[0][22] * mat_B[22][27] +
                  mat_A[0][23] * mat_B[23][27] +
                  mat_A[0][24] * mat_B[24][27] +
                  mat_A[0][25] * mat_B[25][27] +
                  mat_A[0][26] * mat_B[26][27] +
                  mat_A[0][27] * mat_B[27][27] +
                  mat_A[0][28] * mat_B[28][27] +
                  mat_A[0][29] * mat_B[29][27] +
                  mat_A[0][30] * mat_B[30][27] +
                  mat_A[0][31] * mat_B[31][27];
    mat_C[0][28] <= 
                  mat_A[0][0] * mat_B[0][28] +
                  mat_A[0][1] * mat_B[1][28] +
                  mat_A[0][2] * mat_B[2][28] +
                  mat_A[0][3] * mat_B[3][28] +
                  mat_A[0][4] * mat_B[4][28] +
                  mat_A[0][5] * mat_B[5][28] +
                  mat_A[0][6] * mat_B[6][28] +
                  mat_A[0][7] * mat_B[7][28] +
                  mat_A[0][8] * mat_B[8][28] +
                  mat_A[0][9] * mat_B[9][28] +
                  mat_A[0][10] * mat_B[10][28] +
                  mat_A[0][11] * mat_B[11][28] +
                  mat_A[0][12] * mat_B[12][28] +
                  mat_A[0][13] * mat_B[13][28] +
                  mat_A[0][14] * mat_B[14][28] +
                  mat_A[0][15] * mat_B[15][28] +
                  mat_A[0][16] * mat_B[16][28] +
                  mat_A[0][17] * mat_B[17][28] +
                  mat_A[0][18] * mat_B[18][28] +
                  mat_A[0][19] * mat_B[19][28] +
                  mat_A[0][20] * mat_B[20][28] +
                  mat_A[0][21] * mat_B[21][28] +
                  mat_A[0][22] * mat_B[22][28] +
                  mat_A[0][23] * mat_B[23][28] +
                  mat_A[0][24] * mat_B[24][28] +
                  mat_A[0][25] * mat_B[25][28] +
                  mat_A[0][26] * mat_B[26][28] +
                  mat_A[0][27] * mat_B[27][28] +
                  mat_A[0][28] * mat_B[28][28] +
                  mat_A[0][29] * mat_B[29][28] +
                  mat_A[0][30] * mat_B[30][28] +
                  mat_A[0][31] * mat_B[31][28];
    mat_C[0][29] <= 
                  mat_A[0][0] * mat_B[0][29] +
                  mat_A[0][1] * mat_B[1][29] +
                  mat_A[0][2] * mat_B[2][29] +
                  mat_A[0][3] * mat_B[3][29] +
                  mat_A[0][4] * mat_B[4][29] +
                  mat_A[0][5] * mat_B[5][29] +
                  mat_A[0][6] * mat_B[6][29] +
                  mat_A[0][7] * mat_B[7][29] +
                  mat_A[0][8] * mat_B[8][29] +
                  mat_A[0][9] * mat_B[9][29] +
                  mat_A[0][10] * mat_B[10][29] +
                  mat_A[0][11] * mat_B[11][29] +
                  mat_A[0][12] * mat_B[12][29] +
                  mat_A[0][13] * mat_B[13][29] +
                  mat_A[0][14] * mat_B[14][29] +
                  mat_A[0][15] * mat_B[15][29] +
                  mat_A[0][16] * mat_B[16][29] +
                  mat_A[0][17] * mat_B[17][29] +
                  mat_A[0][18] * mat_B[18][29] +
                  mat_A[0][19] * mat_B[19][29] +
                  mat_A[0][20] * mat_B[20][29] +
                  mat_A[0][21] * mat_B[21][29] +
                  mat_A[0][22] * mat_B[22][29] +
                  mat_A[0][23] * mat_B[23][29] +
                  mat_A[0][24] * mat_B[24][29] +
                  mat_A[0][25] * mat_B[25][29] +
                  mat_A[0][26] * mat_B[26][29] +
                  mat_A[0][27] * mat_B[27][29] +
                  mat_A[0][28] * mat_B[28][29] +
                  mat_A[0][29] * mat_B[29][29] +
                  mat_A[0][30] * mat_B[30][29] +
                  mat_A[0][31] * mat_B[31][29];
    mat_C[0][30] <= 
                  mat_A[0][0] * mat_B[0][30] +
                  mat_A[0][1] * mat_B[1][30] +
                  mat_A[0][2] * mat_B[2][30] +
                  mat_A[0][3] * mat_B[3][30] +
                  mat_A[0][4] * mat_B[4][30] +
                  mat_A[0][5] * mat_B[5][30] +
                  mat_A[0][6] * mat_B[6][30] +
                  mat_A[0][7] * mat_B[7][30] +
                  mat_A[0][8] * mat_B[8][30] +
                  mat_A[0][9] * mat_B[9][30] +
                  mat_A[0][10] * mat_B[10][30] +
                  mat_A[0][11] * mat_B[11][30] +
                  mat_A[0][12] * mat_B[12][30] +
                  mat_A[0][13] * mat_B[13][30] +
                  mat_A[0][14] * mat_B[14][30] +
                  mat_A[0][15] * mat_B[15][30] +
                  mat_A[0][16] * mat_B[16][30] +
                  mat_A[0][17] * mat_B[17][30] +
                  mat_A[0][18] * mat_B[18][30] +
                  mat_A[0][19] * mat_B[19][30] +
                  mat_A[0][20] * mat_B[20][30] +
                  mat_A[0][21] * mat_B[21][30] +
                  mat_A[0][22] * mat_B[22][30] +
                  mat_A[0][23] * mat_B[23][30] +
                  mat_A[0][24] * mat_B[24][30] +
                  mat_A[0][25] * mat_B[25][30] +
                  mat_A[0][26] * mat_B[26][30] +
                  mat_A[0][27] * mat_B[27][30] +
                  mat_A[0][28] * mat_B[28][30] +
                  mat_A[0][29] * mat_B[29][30] +
                  mat_A[0][30] * mat_B[30][30] +
                  mat_A[0][31] * mat_B[31][30];
    mat_C[0][31] <= 
                  mat_A[0][0] * mat_B[0][31] +
                  mat_A[0][1] * mat_B[1][31] +
                  mat_A[0][2] * mat_B[2][31] +
                  mat_A[0][3] * mat_B[3][31] +
                  mat_A[0][4] * mat_B[4][31] +
                  mat_A[0][5] * mat_B[5][31] +
                  mat_A[0][6] * mat_B[6][31] +
                  mat_A[0][7] * mat_B[7][31] +
                  mat_A[0][8] * mat_B[8][31] +
                  mat_A[0][9] * mat_B[9][31] +
                  mat_A[0][10] * mat_B[10][31] +
                  mat_A[0][11] * mat_B[11][31] +
                  mat_A[0][12] * mat_B[12][31] +
                  mat_A[0][13] * mat_B[13][31] +
                  mat_A[0][14] * mat_B[14][31] +
                  mat_A[0][15] * mat_B[15][31] +
                  mat_A[0][16] * mat_B[16][31] +
                  mat_A[0][17] * mat_B[17][31] +
                  mat_A[0][18] * mat_B[18][31] +
                  mat_A[0][19] * mat_B[19][31] +
                  mat_A[0][20] * mat_B[20][31] +
                  mat_A[0][21] * mat_B[21][31] +
                  mat_A[0][22] * mat_B[22][31] +
                  mat_A[0][23] * mat_B[23][31] +
                  mat_A[0][24] * mat_B[24][31] +
                  mat_A[0][25] * mat_B[25][31] +
                  mat_A[0][26] * mat_B[26][31] +
                  mat_A[0][27] * mat_B[27][31] +
                  mat_A[0][28] * mat_B[28][31] +
                  mat_A[0][29] * mat_B[29][31] +
                  mat_A[0][30] * mat_B[30][31] +
                  mat_A[0][31] * mat_B[31][31];
    mat_C[1][0] <= 
                  mat_A[1][0] * mat_B[0][0] +
                  mat_A[1][1] * mat_B[1][0] +
                  mat_A[1][2] * mat_B[2][0] +
                  mat_A[1][3] * mat_B[3][0] +
                  mat_A[1][4] * mat_B[4][0] +
                  mat_A[1][5] * mat_B[5][0] +
                  mat_A[1][6] * mat_B[6][0] +
                  mat_A[1][7] * mat_B[7][0] +
                  mat_A[1][8] * mat_B[8][0] +
                  mat_A[1][9] * mat_B[9][0] +
                  mat_A[1][10] * mat_B[10][0] +
                  mat_A[1][11] * mat_B[11][0] +
                  mat_A[1][12] * mat_B[12][0] +
                  mat_A[1][13] * mat_B[13][0] +
                  mat_A[1][14] * mat_B[14][0] +
                  mat_A[1][15] * mat_B[15][0] +
                  mat_A[1][16] * mat_B[16][0] +
                  mat_A[1][17] * mat_B[17][0] +
                  mat_A[1][18] * mat_B[18][0] +
                  mat_A[1][19] * mat_B[19][0] +
                  mat_A[1][20] * mat_B[20][0] +
                  mat_A[1][21] * mat_B[21][0] +
                  mat_A[1][22] * mat_B[22][0] +
                  mat_A[1][23] * mat_B[23][0] +
                  mat_A[1][24] * mat_B[24][0] +
                  mat_A[1][25] * mat_B[25][0] +
                  mat_A[1][26] * mat_B[26][0] +
                  mat_A[1][27] * mat_B[27][0] +
                  mat_A[1][28] * mat_B[28][0] +
                  mat_A[1][29] * mat_B[29][0] +
                  mat_A[1][30] * mat_B[30][0] +
                  mat_A[1][31] * mat_B[31][0];
    mat_C[1][1] <= 
                  mat_A[1][0] * mat_B[0][1] +
                  mat_A[1][1] * mat_B[1][1] +
                  mat_A[1][2] * mat_B[2][1] +
                  mat_A[1][3] * mat_B[3][1] +
                  mat_A[1][4] * mat_B[4][1] +
                  mat_A[1][5] * mat_B[5][1] +
                  mat_A[1][6] * mat_B[6][1] +
                  mat_A[1][7] * mat_B[7][1] +
                  mat_A[1][8] * mat_B[8][1] +
                  mat_A[1][9] * mat_B[9][1] +
                  mat_A[1][10] * mat_B[10][1] +
                  mat_A[1][11] * mat_B[11][1] +
                  mat_A[1][12] * mat_B[12][1] +
                  mat_A[1][13] * mat_B[13][1] +
                  mat_A[1][14] * mat_B[14][1] +
                  mat_A[1][15] * mat_B[15][1] +
                  mat_A[1][16] * mat_B[16][1] +
                  mat_A[1][17] * mat_B[17][1] +
                  mat_A[1][18] * mat_B[18][1] +
                  mat_A[1][19] * mat_B[19][1] +
                  mat_A[1][20] * mat_B[20][1] +
                  mat_A[1][21] * mat_B[21][1] +
                  mat_A[1][22] * mat_B[22][1] +
                  mat_A[1][23] * mat_B[23][1] +
                  mat_A[1][24] * mat_B[24][1] +
                  mat_A[1][25] * mat_B[25][1] +
                  mat_A[1][26] * mat_B[26][1] +
                  mat_A[1][27] * mat_B[27][1] +
                  mat_A[1][28] * mat_B[28][1] +
                  mat_A[1][29] * mat_B[29][1] +
                  mat_A[1][30] * mat_B[30][1] +
                  mat_A[1][31] * mat_B[31][1];
    mat_C[1][2] <= 
                  mat_A[1][0] * mat_B[0][2] +
                  mat_A[1][1] * mat_B[1][2] +
                  mat_A[1][2] * mat_B[2][2] +
                  mat_A[1][3] * mat_B[3][2] +
                  mat_A[1][4] * mat_B[4][2] +
                  mat_A[1][5] * mat_B[5][2] +
                  mat_A[1][6] * mat_B[6][2] +
                  mat_A[1][7] * mat_B[7][2] +
                  mat_A[1][8] * mat_B[8][2] +
                  mat_A[1][9] * mat_B[9][2] +
                  mat_A[1][10] * mat_B[10][2] +
                  mat_A[1][11] * mat_B[11][2] +
                  mat_A[1][12] * mat_B[12][2] +
                  mat_A[1][13] * mat_B[13][2] +
                  mat_A[1][14] * mat_B[14][2] +
                  mat_A[1][15] * mat_B[15][2] +
                  mat_A[1][16] * mat_B[16][2] +
                  mat_A[1][17] * mat_B[17][2] +
                  mat_A[1][18] * mat_B[18][2] +
                  mat_A[1][19] * mat_B[19][2] +
                  mat_A[1][20] * mat_B[20][2] +
                  mat_A[1][21] * mat_B[21][2] +
                  mat_A[1][22] * mat_B[22][2] +
                  mat_A[1][23] * mat_B[23][2] +
                  mat_A[1][24] * mat_B[24][2] +
                  mat_A[1][25] * mat_B[25][2] +
                  mat_A[1][26] * mat_B[26][2] +
                  mat_A[1][27] * mat_B[27][2] +
                  mat_A[1][28] * mat_B[28][2] +
                  mat_A[1][29] * mat_B[29][2] +
                  mat_A[1][30] * mat_B[30][2] +
                  mat_A[1][31] * mat_B[31][2];
    mat_C[1][3] <= 
                  mat_A[1][0] * mat_B[0][3] +
                  mat_A[1][1] * mat_B[1][3] +
                  mat_A[1][2] * mat_B[2][3] +
                  mat_A[1][3] * mat_B[3][3] +
                  mat_A[1][4] * mat_B[4][3] +
                  mat_A[1][5] * mat_B[5][3] +
                  mat_A[1][6] * mat_B[6][3] +
                  mat_A[1][7] * mat_B[7][3] +
                  mat_A[1][8] * mat_B[8][3] +
                  mat_A[1][9] * mat_B[9][3] +
                  mat_A[1][10] * mat_B[10][3] +
                  mat_A[1][11] * mat_B[11][3] +
                  mat_A[1][12] * mat_B[12][3] +
                  mat_A[1][13] * mat_B[13][3] +
                  mat_A[1][14] * mat_B[14][3] +
                  mat_A[1][15] * mat_B[15][3] +
                  mat_A[1][16] * mat_B[16][3] +
                  mat_A[1][17] * mat_B[17][3] +
                  mat_A[1][18] * mat_B[18][3] +
                  mat_A[1][19] * mat_B[19][3] +
                  mat_A[1][20] * mat_B[20][3] +
                  mat_A[1][21] * mat_B[21][3] +
                  mat_A[1][22] * mat_B[22][3] +
                  mat_A[1][23] * mat_B[23][3] +
                  mat_A[1][24] * mat_B[24][3] +
                  mat_A[1][25] * mat_B[25][3] +
                  mat_A[1][26] * mat_B[26][3] +
                  mat_A[1][27] * mat_B[27][3] +
                  mat_A[1][28] * mat_B[28][3] +
                  mat_A[1][29] * mat_B[29][3] +
                  mat_A[1][30] * mat_B[30][3] +
                  mat_A[1][31] * mat_B[31][3];
    mat_C[1][4] <= 
                  mat_A[1][0] * mat_B[0][4] +
                  mat_A[1][1] * mat_B[1][4] +
                  mat_A[1][2] * mat_B[2][4] +
                  mat_A[1][3] * mat_B[3][4] +
                  mat_A[1][4] * mat_B[4][4] +
                  mat_A[1][5] * mat_B[5][4] +
                  mat_A[1][6] * mat_B[6][4] +
                  mat_A[1][7] * mat_B[7][4] +
                  mat_A[1][8] * mat_B[8][4] +
                  mat_A[1][9] * mat_B[9][4] +
                  mat_A[1][10] * mat_B[10][4] +
                  mat_A[1][11] * mat_B[11][4] +
                  mat_A[1][12] * mat_B[12][4] +
                  mat_A[1][13] * mat_B[13][4] +
                  mat_A[1][14] * mat_B[14][4] +
                  mat_A[1][15] * mat_B[15][4] +
                  mat_A[1][16] * mat_B[16][4] +
                  mat_A[1][17] * mat_B[17][4] +
                  mat_A[1][18] * mat_B[18][4] +
                  mat_A[1][19] * mat_B[19][4] +
                  mat_A[1][20] * mat_B[20][4] +
                  mat_A[1][21] * mat_B[21][4] +
                  mat_A[1][22] * mat_B[22][4] +
                  mat_A[1][23] * mat_B[23][4] +
                  mat_A[1][24] * mat_B[24][4] +
                  mat_A[1][25] * mat_B[25][4] +
                  mat_A[1][26] * mat_B[26][4] +
                  mat_A[1][27] * mat_B[27][4] +
                  mat_A[1][28] * mat_B[28][4] +
                  mat_A[1][29] * mat_B[29][4] +
                  mat_A[1][30] * mat_B[30][4] +
                  mat_A[1][31] * mat_B[31][4];
    mat_C[1][5] <= 
                  mat_A[1][0] * mat_B[0][5] +
                  mat_A[1][1] * mat_B[1][5] +
                  mat_A[1][2] * mat_B[2][5] +
                  mat_A[1][3] * mat_B[3][5] +
                  mat_A[1][4] * mat_B[4][5] +
                  mat_A[1][5] * mat_B[5][5] +
                  mat_A[1][6] * mat_B[6][5] +
                  mat_A[1][7] * mat_B[7][5] +
                  mat_A[1][8] * mat_B[8][5] +
                  mat_A[1][9] * mat_B[9][5] +
                  mat_A[1][10] * mat_B[10][5] +
                  mat_A[1][11] * mat_B[11][5] +
                  mat_A[1][12] * mat_B[12][5] +
                  mat_A[1][13] * mat_B[13][5] +
                  mat_A[1][14] * mat_B[14][5] +
                  mat_A[1][15] * mat_B[15][5] +
                  mat_A[1][16] * mat_B[16][5] +
                  mat_A[1][17] * mat_B[17][5] +
                  mat_A[1][18] * mat_B[18][5] +
                  mat_A[1][19] * mat_B[19][5] +
                  mat_A[1][20] * mat_B[20][5] +
                  mat_A[1][21] * mat_B[21][5] +
                  mat_A[1][22] * mat_B[22][5] +
                  mat_A[1][23] * mat_B[23][5] +
                  mat_A[1][24] * mat_B[24][5] +
                  mat_A[1][25] * mat_B[25][5] +
                  mat_A[1][26] * mat_B[26][5] +
                  mat_A[1][27] * mat_B[27][5] +
                  mat_A[1][28] * mat_B[28][5] +
                  mat_A[1][29] * mat_B[29][5] +
                  mat_A[1][30] * mat_B[30][5] +
                  mat_A[1][31] * mat_B[31][5];
    mat_C[1][6] <= 
                  mat_A[1][0] * mat_B[0][6] +
                  mat_A[1][1] * mat_B[1][6] +
                  mat_A[1][2] * mat_B[2][6] +
                  mat_A[1][3] * mat_B[3][6] +
                  mat_A[1][4] * mat_B[4][6] +
                  mat_A[1][5] * mat_B[5][6] +
                  mat_A[1][6] * mat_B[6][6] +
                  mat_A[1][7] * mat_B[7][6] +
                  mat_A[1][8] * mat_B[8][6] +
                  mat_A[1][9] * mat_B[9][6] +
                  mat_A[1][10] * mat_B[10][6] +
                  mat_A[1][11] * mat_B[11][6] +
                  mat_A[1][12] * mat_B[12][6] +
                  mat_A[1][13] * mat_B[13][6] +
                  mat_A[1][14] * mat_B[14][6] +
                  mat_A[1][15] * mat_B[15][6] +
                  mat_A[1][16] * mat_B[16][6] +
                  mat_A[1][17] * mat_B[17][6] +
                  mat_A[1][18] * mat_B[18][6] +
                  mat_A[1][19] * mat_B[19][6] +
                  mat_A[1][20] * mat_B[20][6] +
                  mat_A[1][21] * mat_B[21][6] +
                  mat_A[1][22] * mat_B[22][6] +
                  mat_A[1][23] * mat_B[23][6] +
                  mat_A[1][24] * mat_B[24][6] +
                  mat_A[1][25] * mat_B[25][6] +
                  mat_A[1][26] * mat_B[26][6] +
                  mat_A[1][27] * mat_B[27][6] +
                  mat_A[1][28] * mat_B[28][6] +
                  mat_A[1][29] * mat_B[29][6] +
                  mat_A[1][30] * mat_B[30][6] +
                  mat_A[1][31] * mat_B[31][6];
    mat_C[1][7] <= 
                  mat_A[1][0] * mat_B[0][7] +
                  mat_A[1][1] * mat_B[1][7] +
                  mat_A[1][2] * mat_B[2][7] +
                  mat_A[1][3] * mat_B[3][7] +
                  mat_A[1][4] * mat_B[4][7] +
                  mat_A[1][5] * mat_B[5][7] +
                  mat_A[1][6] * mat_B[6][7] +
                  mat_A[1][7] * mat_B[7][7] +
                  mat_A[1][8] * mat_B[8][7] +
                  mat_A[1][9] * mat_B[9][7] +
                  mat_A[1][10] * mat_B[10][7] +
                  mat_A[1][11] * mat_B[11][7] +
                  mat_A[1][12] * mat_B[12][7] +
                  mat_A[1][13] * mat_B[13][7] +
                  mat_A[1][14] * mat_B[14][7] +
                  mat_A[1][15] * mat_B[15][7] +
                  mat_A[1][16] * mat_B[16][7] +
                  mat_A[1][17] * mat_B[17][7] +
                  mat_A[1][18] * mat_B[18][7] +
                  mat_A[1][19] * mat_B[19][7] +
                  mat_A[1][20] * mat_B[20][7] +
                  mat_A[1][21] * mat_B[21][7] +
                  mat_A[1][22] * mat_B[22][7] +
                  mat_A[1][23] * mat_B[23][7] +
                  mat_A[1][24] * mat_B[24][7] +
                  mat_A[1][25] * mat_B[25][7] +
                  mat_A[1][26] * mat_B[26][7] +
                  mat_A[1][27] * mat_B[27][7] +
                  mat_A[1][28] * mat_B[28][7] +
                  mat_A[1][29] * mat_B[29][7] +
                  mat_A[1][30] * mat_B[30][7] +
                  mat_A[1][31] * mat_B[31][7];
    mat_C[1][8] <= 
                  mat_A[1][0] * mat_B[0][8] +
                  mat_A[1][1] * mat_B[1][8] +
                  mat_A[1][2] * mat_B[2][8] +
                  mat_A[1][3] * mat_B[3][8] +
                  mat_A[1][4] * mat_B[4][8] +
                  mat_A[1][5] * mat_B[5][8] +
                  mat_A[1][6] * mat_B[6][8] +
                  mat_A[1][7] * mat_B[7][8] +
                  mat_A[1][8] * mat_B[8][8] +
                  mat_A[1][9] * mat_B[9][8] +
                  mat_A[1][10] * mat_B[10][8] +
                  mat_A[1][11] * mat_B[11][8] +
                  mat_A[1][12] * mat_B[12][8] +
                  mat_A[1][13] * mat_B[13][8] +
                  mat_A[1][14] * mat_B[14][8] +
                  mat_A[1][15] * mat_B[15][8] +
                  mat_A[1][16] * mat_B[16][8] +
                  mat_A[1][17] * mat_B[17][8] +
                  mat_A[1][18] * mat_B[18][8] +
                  mat_A[1][19] * mat_B[19][8] +
                  mat_A[1][20] * mat_B[20][8] +
                  mat_A[1][21] * mat_B[21][8] +
                  mat_A[1][22] * mat_B[22][8] +
                  mat_A[1][23] * mat_B[23][8] +
                  mat_A[1][24] * mat_B[24][8] +
                  mat_A[1][25] * mat_B[25][8] +
                  mat_A[1][26] * mat_B[26][8] +
                  mat_A[1][27] * mat_B[27][8] +
                  mat_A[1][28] * mat_B[28][8] +
                  mat_A[1][29] * mat_B[29][8] +
                  mat_A[1][30] * mat_B[30][8] +
                  mat_A[1][31] * mat_B[31][8];
    mat_C[1][9] <= 
                  mat_A[1][0] * mat_B[0][9] +
                  mat_A[1][1] * mat_B[1][9] +
                  mat_A[1][2] * mat_B[2][9] +
                  mat_A[1][3] * mat_B[3][9] +
                  mat_A[1][4] * mat_B[4][9] +
                  mat_A[1][5] * mat_B[5][9] +
                  mat_A[1][6] * mat_B[6][9] +
                  mat_A[1][7] * mat_B[7][9] +
                  mat_A[1][8] * mat_B[8][9] +
                  mat_A[1][9] * mat_B[9][9] +
                  mat_A[1][10] * mat_B[10][9] +
                  mat_A[1][11] * mat_B[11][9] +
                  mat_A[1][12] * mat_B[12][9] +
                  mat_A[1][13] * mat_B[13][9] +
                  mat_A[1][14] * mat_B[14][9] +
                  mat_A[1][15] * mat_B[15][9] +
                  mat_A[1][16] * mat_B[16][9] +
                  mat_A[1][17] * mat_B[17][9] +
                  mat_A[1][18] * mat_B[18][9] +
                  mat_A[1][19] * mat_B[19][9] +
                  mat_A[1][20] * mat_B[20][9] +
                  mat_A[1][21] * mat_B[21][9] +
                  mat_A[1][22] * mat_B[22][9] +
                  mat_A[1][23] * mat_B[23][9] +
                  mat_A[1][24] * mat_B[24][9] +
                  mat_A[1][25] * mat_B[25][9] +
                  mat_A[1][26] * mat_B[26][9] +
                  mat_A[1][27] * mat_B[27][9] +
                  mat_A[1][28] * mat_B[28][9] +
                  mat_A[1][29] * mat_B[29][9] +
                  mat_A[1][30] * mat_B[30][9] +
                  mat_A[1][31] * mat_B[31][9];
    mat_C[1][10] <= 
                  mat_A[1][0] * mat_B[0][10] +
                  mat_A[1][1] * mat_B[1][10] +
                  mat_A[1][2] * mat_B[2][10] +
                  mat_A[1][3] * mat_B[3][10] +
                  mat_A[1][4] * mat_B[4][10] +
                  mat_A[1][5] * mat_B[5][10] +
                  mat_A[1][6] * mat_B[6][10] +
                  mat_A[1][7] * mat_B[7][10] +
                  mat_A[1][8] * mat_B[8][10] +
                  mat_A[1][9] * mat_B[9][10] +
                  mat_A[1][10] * mat_B[10][10] +
                  mat_A[1][11] * mat_B[11][10] +
                  mat_A[1][12] * mat_B[12][10] +
                  mat_A[1][13] * mat_B[13][10] +
                  mat_A[1][14] * mat_B[14][10] +
                  mat_A[1][15] * mat_B[15][10] +
                  mat_A[1][16] * mat_B[16][10] +
                  mat_A[1][17] * mat_B[17][10] +
                  mat_A[1][18] * mat_B[18][10] +
                  mat_A[1][19] * mat_B[19][10] +
                  mat_A[1][20] * mat_B[20][10] +
                  mat_A[1][21] * mat_B[21][10] +
                  mat_A[1][22] * mat_B[22][10] +
                  mat_A[1][23] * mat_B[23][10] +
                  mat_A[1][24] * mat_B[24][10] +
                  mat_A[1][25] * mat_B[25][10] +
                  mat_A[1][26] * mat_B[26][10] +
                  mat_A[1][27] * mat_B[27][10] +
                  mat_A[1][28] * mat_B[28][10] +
                  mat_A[1][29] * mat_B[29][10] +
                  mat_A[1][30] * mat_B[30][10] +
                  mat_A[1][31] * mat_B[31][10];
    mat_C[1][11] <= 
                  mat_A[1][0] * mat_B[0][11] +
                  mat_A[1][1] * mat_B[1][11] +
                  mat_A[1][2] * mat_B[2][11] +
                  mat_A[1][3] * mat_B[3][11] +
                  mat_A[1][4] * mat_B[4][11] +
                  mat_A[1][5] * mat_B[5][11] +
                  mat_A[1][6] * mat_B[6][11] +
                  mat_A[1][7] * mat_B[7][11] +
                  mat_A[1][8] * mat_B[8][11] +
                  mat_A[1][9] * mat_B[9][11] +
                  mat_A[1][10] * mat_B[10][11] +
                  mat_A[1][11] * mat_B[11][11] +
                  mat_A[1][12] * mat_B[12][11] +
                  mat_A[1][13] * mat_B[13][11] +
                  mat_A[1][14] * mat_B[14][11] +
                  mat_A[1][15] * mat_B[15][11] +
                  mat_A[1][16] * mat_B[16][11] +
                  mat_A[1][17] * mat_B[17][11] +
                  mat_A[1][18] * mat_B[18][11] +
                  mat_A[1][19] * mat_B[19][11] +
                  mat_A[1][20] * mat_B[20][11] +
                  mat_A[1][21] * mat_B[21][11] +
                  mat_A[1][22] * mat_B[22][11] +
                  mat_A[1][23] * mat_B[23][11] +
                  mat_A[1][24] * mat_B[24][11] +
                  mat_A[1][25] * mat_B[25][11] +
                  mat_A[1][26] * mat_B[26][11] +
                  mat_A[1][27] * mat_B[27][11] +
                  mat_A[1][28] * mat_B[28][11] +
                  mat_A[1][29] * mat_B[29][11] +
                  mat_A[1][30] * mat_B[30][11] +
                  mat_A[1][31] * mat_B[31][11];
    mat_C[1][12] <= 
                  mat_A[1][0] * mat_B[0][12] +
                  mat_A[1][1] * mat_B[1][12] +
                  mat_A[1][2] * mat_B[2][12] +
                  mat_A[1][3] * mat_B[3][12] +
                  mat_A[1][4] * mat_B[4][12] +
                  mat_A[1][5] * mat_B[5][12] +
                  mat_A[1][6] * mat_B[6][12] +
                  mat_A[1][7] * mat_B[7][12] +
                  mat_A[1][8] * mat_B[8][12] +
                  mat_A[1][9] * mat_B[9][12] +
                  mat_A[1][10] * mat_B[10][12] +
                  mat_A[1][11] * mat_B[11][12] +
                  mat_A[1][12] * mat_B[12][12] +
                  mat_A[1][13] * mat_B[13][12] +
                  mat_A[1][14] * mat_B[14][12] +
                  mat_A[1][15] * mat_B[15][12] +
                  mat_A[1][16] * mat_B[16][12] +
                  mat_A[1][17] * mat_B[17][12] +
                  mat_A[1][18] * mat_B[18][12] +
                  mat_A[1][19] * mat_B[19][12] +
                  mat_A[1][20] * mat_B[20][12] +
                  mat_A[1][21] * mat_B[21][12] +
                  mat_A[1][22] * mat_B[22][12] +
                  mat_A[1][23] * mat_B[23][12] +
                  mat_A[1][24] * mat_B[24][12] +
                  mat_A[1][25] * mat_B[25][12] +
                  mat_A[1][26] * mat_B[26][12] +
                  mat_A[1][27] * mat_B[27][12] +
                  mat_A[1][28] * mat_B[28][12] +
                  mat_A[1][29] * mat_B[29][12] +
                  mat_A[1][30] * mat_B[30][12] +
                  mat_A[1][31] * mat_B[31][12];
    mat_C[1][13] <= 
                  mat_A[1][0] * mat_B[0][13] +
                  mat_A[1][1] * mat_B[1][13] +
                  mat_A[1][2] * mat_B[2][13] +
                  mat_A[1][3] * mat_B[3][13] +
                  mat_A[1][4] * mat_B[4][13] +
                  mat_A[1][5] * mat_B[5][13] +
                  mat_A[1][6] * mat_B[6][13] +
                  mat_A[1][7] * mat_B[7][13] +
                  mat_A[1][8] * mat_B[8][13] +
                  mat_A[1][9] * mat_B[9][13] +
                  mat_A[1][10] * mat_B[10][13] +
                  mat_A[1][11] * mat_B[11][13] +
                  mat_A[1][12] * mat_B[12][13] +
                  mat_A[1][13] * mat_B[13][13] +
                  mat_A[1][14] * mat_B[14][13] +
                  mat_A[1][15] * mat_B[15][13] +
                  mat_A[1][16] * mat_B[16][13] +
                  mat_A[1][17] * mat_B[17][13] +
                  mat_A[1][18] * mat_B[18][13] +
                  mat_A[1][19] * mat_B[19][13] +
                  mat_A[1][20] * mat_B[20][13] +
                  mat_A[1][21] * mat_B[21][13] +
                  mat_A[1][22] * mat_B[22][13] +
                  mat_A[1][23] * mat_B[23][13] +
                  mat_A[1][24] * mat_B[24][13] +
                  mat_A[1][25] * mat_B[25][13] +
                  mat_A[1][26] * mat_B[26][13] +
                  mat_A[1][27] * mat_B[27][13] +
                  mat_A[1][28] * mat_B[28][13] +
                  mat_A[1][29] * mat_B[29][13] +
                  mat_A[1][30] * mat_B[30][13] +
                  mat_A[1][31] * mat_B[31][13];
    mat_C[1][14] <= 
                  mat_A[1][0] * mat_B[0][14] +
                  mat_A[1][1] * mat_B[1][14] +
                  mat_A[1][2] * mat_B[2][14] +
                  mat_A[1][3] * mat_B[3][14] +
                  mat_A[1][4] * mat_B[4][14] +
                  mat_A[1][5] * mat_B[5][14] +
                  mat_A[1][6] * mat_B[6][14] +
                  mat_A[1][7] * mat_B[7][14] +
                  mat_A[1][8] * mat_B[8][14] +
                  mat_A[1][9] * mat_B[9][14] +
                  mat_A[1][10] * mat_B[10][14] +
                  mat_A[1][11] * mat_B[11][14] +
                  mat_A[1][12] * mat_B[12][14] +
                  mat_A[1][13] * mat_B[13][14] +
                  mat_A[1][14] * mat_B[14][14] +
                  mat_A[1][15] * mat_B[15][14] +
                  mat_A[1][16] * mat_B[16][14] +
                  mat_A[1][17] * mat_B[17][14] +
                  mat_A[1][18] * mat_B[18][14] +
                  mat_A[1][19] * mat_B[19][14] +
                  mat_A[1][20] * mat_B[20][14] +
                  mat_A[1][21] * mat_B[21][14] +
                  mat_A[1][22] * mat_B[22][14] +
                  mat_A[1][23] * mat_B[23][14] +
                  mat_A[1][24] * mat_B[24][14] +
                  mat_A[1][25] * mat_B[25][14] +
                  mat_A[1][26] * mat_B[26][14] +
                  mat_A[1][27] * mat_B[27][14] +
                  mat_A[1][28] * mat_B[28][14] +
                  mat_A[1][29] * mat_B[29][14] +
                  mat_A[1][30] * mat_B[30][14] +
                  mat_A[1][31] * mat_B[31][14];
    mat_C[1][15] <= 
                  mat_A[1][0] * mat_B[0][15] +
                  mat_A[1][1] * mat_B[1][15] +
                  mat_A[1][2] * mat_B[2][15] +
                  mat_A[1][3] * mat_B[3][15] +
                  mat_A[1][4] * mat_B[4][15] +
                  mat_A[1][5] * mat_B[5][15] +
                  mat_A[1][6] * mat_B[6][15] +
                  mat_A[1][7] * mat_B[7][15] +
                  mat_A[1][8] * mat_B[8][15] +
                  mat_A[1][9] * mat_B[9][15] +
                  mat_A[1][10] * mat_B[10][15] +
                  mat_A[1][11] * mat_B[11][15] +
                  mat_A[1][12] * mat_B[12][15] +
                  mat_A[1][13] * mat_B[13][15] +
                  mat_A[1][14] * mat_B[14][15] +
                  mat_A[1][15] * mat_B[15][15] +
                  mat_A[1][16] * mat_B[16][15] +
                  mat_A[1][17] * mat_B[17][15] +
                  mat_A[1][18] * mat_B[18][15] +
                  mat_A[1][19] * mat_B[19][15] +
                  mat_A[1][20] * mat_B[20][15] +
                  mat_A[1][21] * mat_B[21][15] +
                  mat_A[1][22] * mat_B[22][15] +
                  mat_A[1][23] * mat_B[23][15] +
                  mat_A[1][24] * mat_B[24][15] +
                  mat_A[1][25] * mat_B[25][15] +
                  mat_A[1][26] * mat_B[26][15] +
                  mat_A[1][27] * mat_B[27][15] +
                  mat_A[1][28] * mat_B[28][15] +
                  mat_A[1][29] * mat_B[29][15] +
                  mat_A[1][30] * mat_B[30][15] +
                  mat_A[1][31] * mat_B[31][15];
    mat_C[1][16] <= 
                  mat_A[1][0] * mat_B[0][16] +
                  mat_A[1][1] * mat_B[1][16] +
                  mat_A[1][2] * mat_B[2][16] +
                  mat_A[1][3] * mat_B[3][16] +
                  mat_A[1][4] * mat_B[4][16] +
                  mat_A[1][5] * mat_B[5][16] +
                  mat_A[1][6] * mat_B[6][16] +
                  mat_A[1][7] * mat_B[7][16] +
                  mat_A[1][8] * mat_B[8][16] +
                  mat_A[1][9] * mat_B[9][16] +
                  mat_A[1][10] * mat_B[10][16] +
                  mat_A[1][11] * mat_B[11][16] +
                  mat_A[1][12] * mat_B[12][16] +
                  mat_A[1][13] * mat_B[13][16] +
                  mat_A[1][14] * mat_B[14][16] +
                  mat_A[1][15] * mat_B[15][16] +
                  mat_A[1][16] * mat_B[16][16] +
                  mat_A[1][17] * mat_B[17][16] +
                  mat_A[1][18] * mat_B[18][16] +
                  mat_A[1][19] * mat_B[19][16] +
                  mat_A[1][20] * mat_B[20][16] +
                  mat_A[1][21] * mat_B[21][16] +
                  mat_A[1][22] * mat_B[22][16] +
                  mat_A[1][23] * mat_B[23][16] +
                  mat_A[1][24] * mat_B[24][16] +
                  mat_A[1][25] * mat_B[25][16] +
                  mat_A[1][26] * mat_B[26][16] +
                  mat_A[1][27] * mat_B[27][16] +
                  mat_A[1][28] * mat_B[28][16] +
                  mat_A[1][29] * mat_B[29][16] +
                  mat_A[1][30] * mat_B[30][16] +
                  mat_A[1][31] * mat_B[31][16];
    mat_C[1][17] <= 
                  mat_A[1][0] * mat_B[0][17] +
                  mat_A[1][1] * mat_B[1][17] +
                  mat_A[1][2] * mat_B[2][17] +
                  mat_A[1][3] * mat_B[3][17] +
                  mat_A[1][4] * mat_B[4][17] +
                  mat_A[1][5] * mat_B[5][17] +
                  mat_A[1][6] * mat_B[6][17] +
                  mat_A[1][7] * mat_B[7][17] +
                  mat_A[1][8] * mat_B[8][17] +
                  mat_A[1][9] * mat_B[9][17] +
                  mat_A[1][10] * mat_B[10][17] +
                  mat_A[1][11] * mat_B[11][17] +
                  mat_A[1][12] * mat_B[12][17] +
                  mat_A[1][13] * mat_B[13][17] +
                  mat_A[1][14] * mat_B[14][17] +
                  mat_A[1][15] * mat_B[15][17] +
                  mat_A[1][16] * mat_B[16][17] +
                  mat_A[1][17] * mat_B[17][17] +
                  mat_A[1][18] * mat_B[18][17] +
                  mat_A[1][19] * mat_B[19][17] +
                  mat_A[1][20] * mat_B[20][17] +
                  mat_A[1][21] * mat_B[21][17] +
                  mat_A[1][22] * mat_B[22][17] +
                  mat_A[1][23] * mat_B[23][17] +
                  mat_A[1][24] * mat_B[24][17] +
                  mat_A[1][25] * mat_B[25][17] +
                  mat_A[1][26] * mat_B[26][17] +
                  mat_A[1][27] * mat_B[27][17] +
                  mat_A[1][28] * mat_B[28][17] +
                  mat_A[1][29] * mat_B[29][17] +
                  mat_A[1][30] * mat_B[30][17] +
                  mat_A[1][31] * mat_B[31][17];
    mat_C[1][18] <= 
                  mat_A[1][0] * mat_B[0][18] +
                  mat_A[1][1] * mat_B[1][18] +
                  mat_A[1][2] * mat_B[2][18] +
                  mat_A[1][3] * mat_B[3][18] +
                  mat_A[1][4] * mat_B[4][18] +
                  mat_A[1][5] * mat_B[5][18] +
                  mat_A[1][6] * mat_B[6][18] +
                  mat_A[1][7] * mat_B[7][18] +
                  mat_A[1][8] * mat_B[8][18] +
                  mat_A[1][9] * mat_B[9][18] +
                  mat_A[1][10] * mat_B[10][18] +
                  mat_A[1][11] * mat_B[11][18] +
                  mat_A[1][12] * mat_B[12][18] +
                  mat_A[1][13] * mat_B[13][18] +
                  mat_A[1][14] * mat_B[14][18] +
                  mat_A[1][15] * mat_B[15][18] +
                  mat_A[1][16] * mat_B[16][18] +
                  mat_A[1][17] * mat_B[17][18] +
                  mat_A[1][18] * mat_B[18][18] +
                  mat_A[1][19] * mat_B[19][18] +
                  mat_A[1][20] * mat_B[20][18] +
                  mat_A[1][21] * mat_B[21][18] +
                  mat_A[1][22] * mat_B[22][18] +
                  mat_A[1][23] * mat_B[23][18] +
                  mat_A[1][24] * mat_B[24][18] +
                  mat_A[1][25] * mat_B[25][18] +
                  mat_A[1][26] * mat_B[26][18] +
                  mat_A[1][27] * mat_B[27][18] +
                  mat_A[1][28] * mat_B[28][18] +
                  mat_A[1][29] * mat_B[29][18] +
                  mat_A[1][30] * mat_B[30][18] +
                  mat_A[1][31] * mat_B[31][18];
    mat_C[1][19] <= 
                  mat_A[1][0] * mat_B[0][19] +
                  mat_A[1][1] * mat_B[1][19] +
                  mat_A[1][2] * mat_B[2][19] +
                  mat_A[1][3] * mat_B[3][19] +
                  mat_A[1][4] * mat_B[4][19] +
                  mat_A[1][5] * mat_B[5][19] +
                  mat_A[1][6] * mat_B[6][19] +
                  mat_A[1][7] * mat_B[7][19] +
                  mat_A[1][8] * mat_B[8][19] +
                  mat_A[1][9] * mat_B[9][19] +
                  mat_A[1][10] * mat_B[10][19] +
                  mat_A[1][11] * mat_B[11][19] +
                  mat_A[1][12] * mat_B[12][19] +
                  mat_A[1][13] * mat_B[13][19] +
                  mat_A[1][14] * mat_B[14][19] +
                  mat_A[1][15] * mat_B[15][19] +
                  mat_A[1][16] * mat_B[16][19] +
                  mat_A[1][17] * mat_B[17][19] +
                  mat_A[1][18] * mat_B[18][19] +
                  mat_A[1][19] * mat_B[19][19] +
                  mat_A[1][20] * mat_B[20][19] +
                  mat_A[1][21] * mat_B[21][19] +
                  mat_A[1][22] * mat_B[22][19] +
                  mat_A[1][23] * mat_B[23][19] +
                  mat_A[1][24] * mat_B[24][19] +
                  mat_A[1][25] * mat_B[25][19] +
                  mat_A[1][26] * mat_B[26][19] +
                  mat_A[1][27] * mat_B[27][19] +
                  mat_A[1][28] * mat_B[28][19] +
                  mat_A[1][29] * mat_B[29][19] +
                  mat_A[1][30] * mat_B[30][19] +
                  mat_A[1][31] * mat_B[31][19];
    mat_C[1][20] <= 
                  mat_A[1][0] * mat_B[0][20] +
                  mat_A[1][1] * mat_B[1][20] +
                  mat_A[1][2] * mat_B[2][20] +
                  mat_A[1][3] * mat_B[3][20] +
                  mat_A[1][4] * mat_B[4][20] +
                  mat_A[1][5] * mat_B[5][20] +
                  mat_A[1][6] * mat_B[6][20] +
                  mat_A[1][7] * mat_B[7][20] +
                  mat_A[1][8] * mat_B[8][20] +
                  mat_A[1][9] * mat_B[9][20] +
                  mat_A[1][10] * mat_B[10][20] +
                  mat_A[1][11] * mat_B[11][20] +
                  mat_A[1][12] * mat_B[12][20] +
                  mat_A[1][13] * mat_B[13][20] +
                  mat_A[1][14] * mat_B[14][20] +
                  mat_A[1][15] * mat_B[15][20] +
                  mat_A[1][16] * mat_B[16][20] +
                  mat_A[1][17] * mat_B[17][20] +
                  mat_A[1][18] * mat_B[18][20] +
                  mat_A[1][19] * mat_B[19][20] +
                  mat_A[1][20] * mat_B[20][20] +
                  mat_A[1][21] * mat_B[21][20] +
                  mat_A[1][22] * mat_B[22][20] +
                  mat_A[1][23] * mat_B[23][20] +
                  mat_A[1][24] * mat_B[24][20] +
                  mat_A[1][25] * mat_B[25][20] +
                  mat_A[1][26] * mat_B[26][20] +
                  mat_A[1][27] * mat_B[27][20] +
                  mat_A[1][28] * mat_B[28][20] +
                  mat_A[1][29] * mat_B[29][20] +
                  mat_A[1][30] * mat_B[30][20] +
                  mat_A[1][31] * mat_B[31][20];
    mat_C[1][21] <= 
                  mat_A[1][0] * mat_B[0][21] +
                  mat_A[1][1] * mat_B[1][21] +
                  mat_A[1][2] * mat_B[2][21] +
                  mat_A[1][3] * mat_B[3][21] +
                  mat_A[1][4] * mat_B[4][21] +
                  mat_A[1][5] * mat_B[5][21] +
                  mat_A[1][6] * mat_B[6][21] +
                  mat_A[1][7] * mat_B[7][21] +
                  mat_A[1][8] * mat_B[8][21] +
                  mat_A[1][9] * mat_B[9][21] +
                  mat_A[1][10] * mat_B[10][21] +
                  mat_A[1][11] * mat_B[11][21] +
                  mat_A[1][12] * mat_B[12][21] +
                  mat_A[1][13] * mat_B[13][21] +
                  mat_A[1][14] * mat_B[14][21] +
                  mat_A[1][15] * mat_B[15][21] +
                  mat_A[1][16] * mat_B[16][21] +
                  mat_A[1][17] * mat_B[17][21] +
                  mat_A[1][18] * mat_B[18][21] +
                  mat_A[1][19] * mat_B[19][21] +
                  mat_A[1][20] * mat_B[20][21] +
                  mat_A[1][21] * mat_B[21][21] +
                  mat_A[1][22] * mat_B[22][21] +
                  mat_A[1][23] * mat_B[23][21] +
                  mat_A[1][24] * mat_B[24][21] +
                  mat_A[1][25] * mat_B[25][21] +
                  mat_A[1][26] * mat_B[26][21] +
                  mat_A[1][27] * mat_B[27][21] +
                  mat_A[1][28] * mat_B[28][21] +
                  mat_A[1][29] * mat_B[29][21] +
                  mat_A[1][30] * mat_B[30][21] +
                  mat_A[1][31] * mat_B[31][21];
    mat_C[1][22] <= 
                  mat_A[1][0] * mat_B[0][22] +
                  mat_A[1][1] * mat_B[1][22] +
                  mat_A[1][2] * mat_B[2][22] +
                  mat_A[1][3] * mat_B[3][22] +
                  mat_A[1][4] * mat_B[4][22] +
                  mat_A[1][5] * mat_B[5][22] +
                  mat_A[1][6] * mat_B[6][22] +
                  mat_A[1][7] * mat_B[7][22] +
                  mat_A[1][8] * mat_B[8][22] +
                  mat_A[1][9] * mat_B[9][22] +
                  mat_A[1][10] * mat_B[10][22] +
                  mat_A[1][11] * mat_B[11][22] +
                  mat_A[1][12] * mat_B[12][22] +
                  mat_A[1][13] * mat_B[13][22] +
                  mat_A[1][14] * mat_B[14][22] +
                  mat_A[1][15] * mat_B[15][22] +
                  mat_A[1][16] * mat_B[16][22] +
                  mat_A[1][17] * mat_B[17][22] +
                  mat_A[1][18] * mat_B[18][22] +
                  mat_A[1][19] * mat_B[19][22] +
                  mat_A[1][20] * mat_B[20][22] +
                  mat_A[1][21] * mat_B[21][22] +
                  mat_A[1][22] * mat_B[22][22] +
                  mat_A[1][23] * mat_B[23][22] +
                  mat_A[1][24] * mat_B[24][22] +
                  mat_A[1][25] * mat_B[25][22] +
                  mat_A[1][26] * mat_B[26][22] +
                  mat_A[1][27] * mat_B[27][22] +
                  mat_A[1][28] * mat_B[28][22] +
                  mat_A[1][29] * mat_B[29][22] +
                  mat_A[1][30] * mat_B[30][22] +
                  mat_A[1][31] * mat_B[31][22];
    mat_C[1][23] <= 
                  mat_A[1][0] * mat_B[0][23] +
                  mat_A[1][1] * mat_B[1][23] +
                  mat_A[1][2] * mat_B[2][23] +
                  mat_A[1][3] * mat_B[3][23] +
                  mat_A[1][4] * mat_B[4][23] +
                  mat_A[1][5] * mat_B[5][23] +
                  mat_A[1][6] * mat_B[6][23] +
                  mat_A[1][7] * mat_B[7][23] +
                  mat_A[1][8] * mat_B[8][23] +
                  mat_A[1][9] * mat_B[9][23] +
                  mat_A[1][10] * mat_B[10][23] +
                  mat_A[1][11] * mat_B[11][23] +
                  mat_A[1][12] * mat_B[12][23] +
                  mat_A[1][13] * mat_B[13][23] +
                  mat_A[1][14] * mat_B[14][23] +
                  mat_A[1][15] * mat_B[15][23] +
                  mat_A[1][16] * mat_B[16][23] +
                  mat_A[1][17] * mat_B[17][23] +
                  mat_A[1][18] * mat_B[18][23] +
                  mat_A[1][19] * mat_B[19][23] +
                  mat_A[1][20] * mat_B[20][23] +
                  mat_A[1][21] * mat_B[21][23] +
                  mat_A[1][22] * mat_B[22][23] +
                  mat_A[1][23] * mat_B[23][23] +
                  mat_A[1][24] * mat_B[24][23] +
                  mat_A[1][25] * mat_B[25][23] +
                  mat_A[1][26] * mat_B[26][23] +
                  mat_A[1][27] * mat_B[27][23] +
                  mat_A[1][28] * mat_B[28][23] +
                  mat_A[1][29] * mat_B[29][23] +
                  mat_A[1][30] * mat_B[30][23] +
                  mat_A[1][31] * mat_B[31][23];
    mat_C[1][24] <= 
                  mat_A[1][0] * mat_B[0][24] +
                  mat_A[1][1] * mat_B[1][24] +
                  mat_A[1][2] * mat_B[2][24] +
                  mat_A[1][3] * mat_B[3][24] +
                  mat_A[1][4] * mat_B[4][24] +
                  mat_A[1][5] * mat_B[5][24] +
                  mat_A[1][6] * mat_B[6][24] +
                  mat_A[1][7] * mat_B[7][24] +
                  mat_A[1][8] * mat_B[8][24] +
                  mat_A[1][9] * mat_B[9][24] +
                  mat_A[1][10] * mat_B[10][24] +
                  mat_A[1][11] * mat_B[11][24] +
                  mat_A[1][12] * mat_B[12][24] +
                  mat_A[1][13] * mat_B[13][24] +
                  mat_A[1][14] * mat_B[14][24] +
                  mat_A[1][15] * mat_B[15][24] +
                  mat_A[1][16] * mat_B[16][24] +
                  mat_A[1][17] * mat_B[17][24] +
                  mat_A[1][18] * mat_B[18][24] +
                  mat_A[1][19] * mat_B[19][24] +
                  mat_A[1][20] * mat_B[20][24] +
                  mat_A[1][21] * mat_B[21][24] +
                  mat_A[1][22] * mat_B[22][24] +
                  mat_A[1][23] * mat_B[23][24] +
                  mat_A[1][24] * mat_B[24][24] +
                  mat_A[1][25] * mat_B[25][24] +
                  mat_A[1][26] * mat_B[26][24] +
                  mat_A[1][27] * mat_B[27][24] +
                  mat_A[1][28] * mat_B[28][24] +
                  mat_A[1][29] * mat_B[29][24] +
                  mat_A[1][30] * mat_B[30][24] +
                  mat_A[1][31] * mat_B[31][24];
    mat_C[1][25] <= 
                  mat_A[1][0] * mat_B[0][25] +
                  mat_A[1][1] * mat_B[1][25] +
                  mat_A[1][2] * mat_B[2][25] +
                  mat_A[1][3] * mat_B[3][25] +
                  mat_A[1][4] * mat_B[4][25] +
                  mat_A[1][5] * mat_B[5][25] +
                  mat_A[1][6] * mat_B[6][25] +
                  mat_A[1][7] * mat_B[7][25] +
                  mat_A[1][8] * mat_B[8][25] +
                  mat_A[1][9] * mat_B[9][25] +
                  mat_A[1][10] * mat_B[10][25] +
                  mat_A[1][11] * mat_B[11][25] +
                  mat_A[1][12] * mat_B[12][25] +
                  mat_A[1][13] * mat_B[13][25] +
                  mat_A[1][14] * mat_B[14][25] +
                  mat_A[1][15] * mat_B[15][25] +
                  mat_A[1][16] * mat_B[16][25] +
                  mat_A[1][17] * mat_B[17][25] +
                  mat_A[1][18] * mat_B[18][25] +
                  mat_A[1][19] * mat_B[19][25] +
                  mat_A[1][20] * mat_B[20][25] +
                  mat_A[1][21] * mat_B[21][25] +
                  mat_A[1][22] * mat_B[22][25] +
                  mat_A[1][23] * mat_B[23][25] +
                  mat_A[1][24] * mat_B[24][25] +
                  mat_A[1][25] * mat_B[25][25] +
                  mat_A[1][26] * mat_B[26][25] +
                  mat_A[1][27] * mat_B[27][25] +
                  mat_A[1][28] * mat_B[28][25] +
                  mat_A[1][29] * mat_B[29][25] +
                  mat_A[1][30] * mat_B[30][25] +
                  mat_A[1][31] * mat_B[31][25];
    mat_C[1][26] <= 
                  mat_A[1][0] * mat_B[0][26] +
                  mat_A[1][1] * mat_B[1][26] +
                  mat_A[1][2] * mat_B[2][26] +
                  mat_A[1][3] * mat_B[3][26] +
                  mat_A[1][4] * mat_B[4][26] +
                  mat_A[1][5] * mat_B[5][26] +
                  mat_A[1][6] * mat_B[6][26] +
                  mat_A[1][7] * mat_B[7][26] +
                  mat_A[1][8] * mat_B[8][26] +
                  mat_A[1][9] * mat_B[9][26] +
                  mat_A[1][10] * mat_B[10][26] +
                  mat_A[1][11] * mat_B[11][26] +
                  mat_A[1][12] * mat_B[12][26] +
                  mat_A[1][13] * mat_B[13][26] +
                  mat_A[1][14] * mat_B[14][26] +
                  mat_A[1][15] * mat_B[15][26] +
                  mat_A[1][16] * mat_B[16][26] +
                  mat_A[1][17] * mat_B[17][26] +
                  mat_A[1][18] * mat_B[18][26] +
                  mat_A[1][19] * mat_B[19][26] +
                  mat_A[1][20] * mat_B[20][26] +
                  mat_A[1][21] * mat_B[21][26] +
                  mat_A[1][22] * mat_B[22][26] +
                  mat_A[1][23] * mat_B[23][26] +
                  mat_A[1][24] * mat_B[24][26] +
                  mat_A[1][25] * mat_B[25][26] +
                  mat_A[1][26] * mat_B[26][26] +
                  mat_A[1][27] * mat_B[27][26] +
                  mat_A[1][28] * mat_B[28][26] +
                  mat_A[1][29] * mat_B[29][26] +
                  mat_A[1][30] * mat_B[30][26] +
                  mat_A[1][31] * mat_B[31][26];
    mat_C[1][27] <= 
                  mat_A[1][0] * mat_B[0][27] +
                  mat_A[1][1] * mat_B[1][27] +
                  mat_A[1][2] * mat_B[2][27] +
                  mat_A[1][3] * mat_B[3][27] +
                  mat_A[1][4] * mat_B[4][27] +
                  mat_A[1][5] * mat_B[5][27] +
                  mat_A[1][6] * mat_B[6][27] +
                  mat_A[1][7] * mat_B[7][27] +
                  mat_A[1][8] * mat_B[8][27] +
                  mat_A[1][9] * mat_B[9][27] +
                  mat_A[1][10] * mat_B[10][27] +
                  mat_A[1][11] * mat_B[11][27] +
                  mat_A[1][12] * mat_B[12][27] +
                  mat_A[1][13] * mat_B[13][27] +
                  mat_A[1][14] * mat_B[14][27] +
                  mat_A[1][15] * mat_B[15][27] +
                  mat_A[1][16] * mat_B[16][27] +
                  mat_A[1][17] * mat_B[17][27] +
                  mat_A[1][18] * mat_B[18][27] +
                  mat_A[1][19] * mat_B[19][27] +
                  mat_A[1][20] * mat_B[20][27] +
                  mat_A[1][21] * mat_B[21][27] +
                  mat_A[1][22] * mat_B[22][27] +
                  mat_A[1][23] * mat_B[23][27] +
                  mat_A[1][24] * mat_B[24][27] +
                  mat_A[1][25] * mat_B[25][27] +
                  mat_A[1][26] * mat_B[26][27] +
                  mat_A[1][27] * mat_B[27][27] +
                  mat_A[1][28] * mat_B[28][27] +
                  mat_A[1][29] * mat_B[29][27] +
                  mat_A[1][30] * mat_B[30][27] +
                  mat_A[1][31] * mat_B[31][27];
    mat_C[1][28] <= 
                  mat_A[1][0] * mat_B[0][28] +
                  mat_A[1][1] * mat_B[1][28] +
                  mat_A[1][2] * mat_B[2][28] +
                  mat_A[1][3] * mat_B[3][28] +
                  mat_A[1][4] * mat_B[4][28] +
                  mat_A[1][5] * mat_B[5][28] +
                  mat_A[1][6] * mat_B[6][28] +
                  mat_A[1][7] * mat_B[7][28] +
                  mat_A[1][8] * mat_B[8][28] +
                  mat_A[1][9] * mat_B[9][28] +
                  mat_A[1][10] * mat_B[10][28] +
                  mat_A[1][11] * mat_B[11][28] +
                  mat_A[1][12] * mat_B[12][28] +
                  mat_A[1][13] * mat_B[13][28] +
                  mat_A[1][14] * mat_B[14][28] +
                  mat_A[1][15] * mat_B[15][28] +
                  mat_A[1][16] * mat_B[16][28] +
                  mat_A[1][17] * mat_B[17][28] +
                  mat_A[1][18] * mat_B[18][28] +
                  mat_A[1][19] * mat_B[19][28] +
                  mat_A[1][20] * mat_B[20][28] +
                  mat_A[1][21] * mat_B[21][28] +
                  mat_A[1][22] * mat_B[22][28] +
                  mat_A[1][23] * mat_B[23][28] +
                  mat_A[1][24] * mat_B[24][28] +
                  mat_A[1][25] * mat_B[25][28] +
                  mat_A[1][26] * mat_B[26][28] +
                  mat_A[1][27] * mat_B[27][28] +
                  mat_A[1][28] * mat_B[28][28] +
                  mat_A[1][29] * mat_B[29][28] +
                  mat_A[1][30] * mat_B[30][28] +
                  mat_A[1][31] * mat_B[31][28];
    mat_C[1][29] <= 
                  mat_A[1][0] * mat_B[0][29] +
                  mat_A[1][1] * mat_B[1][29] +
                  mat_A[1][2] * mat_B[2][29] +
                  mat_A[1][3] * mat_B[3][29] +
                  mat_A[1][4] * mat_B[4][29] +
                  mat_A[1][5] * mat_B[5][29] +
                  mat_A[1][6] * mat_B[6][29] +
                  mat_A[1][7] * mat_B[7][29] +
                  mat_A[1][8] * mat_B[8][29] +
                  mat_A[1][9] * mat_B[9][29] +
                  mat_A[1][10] * mat_B[10][29] +
                  mat_A[1][11] * mat_B[11][29] +
                  mat_A[1][12] * mat_B[12][29] +
                  mat_A[1][13] * mat_B[13][29] +
                  mat_A[1][14] * mat_B[14][29] +
                  mat_A[1][15] * mat_B[15][29] +
                  mat_A[1][16] * mat_B[16][29] +
                  mat_A[1][17] * mat_B[17][29] +
                  mat_A[1][18] * mat_B[18][29] +
                  mat_A[1][19] * mat_B[19][29] +
                  mat_A[1][20] * mat_B[20][29] +
                  mat_A[1][21] * mat_B[21][29] +
                  mat_A[1][22] * mat_B[22][29] +
                  mat_A[1][23] * mat_B[23][29] +
                  mat_A[1][24] * mat_B[24][29] +
                  mat_A[1][25] * mat_B[25][29] +
                  mat_A[1][26] * mat_B[26][29] +
                  mat_A[1][27] * mat_B[27][29] +
                  mat_A[1][28] * mat_B[28][29] +
                  mat_A[1][29] * mat_B[29][29] +
                  mat_A[1][30] * mat_B[30][29] +
                  mat_A[1][31] * mat_B[31][29];
    mat_C[1][30] <= 
                  mat_A[1][0] * mat_B[0][30] +
                  mat_A[1][1] * mat_B[1][30] +
                  mat_A[1][2] * mat_B[2][30] +
                  mat_A[1][3] * mat_B[3][30] +
                  mat_A[1][4] * mat_B[4][30] +
                  mat_A[1][5] * mat_B[5][30] +
                  mat_A[1][6] * mat_B[6][30] +
                  mat_A[1][7] * mat_B[7][30] +
                  mat_A[1][8] * mat_B[8][30] +
                  mat_A[1][9] * mat_B[9][30] +
                  mat_A[1][10] * mat_B[10][30] +
                  mat_A[1][11] * mat_B[11][30] +
                  mat_A[1][12] * mat_B[12][30] +
                  mat_A[1][13] * mat_B[13][30] +
                  mat_A[1][14] * mat_B[14][30] +
                  mat_A[1][15] * mat_B[15][30] +
                  mat_A[1][16] * mat_B[16][30] +
                  mat_A[1][17] * mat_B[17][30] +
                  mat_A[1][18] * mat_B[18][30] +
                  mat_A[1][19] * mat_B[19][30] +
                  mat_A[1][20] * mat_B[20][30] +
                  mat_A[1][21] * mat_B[21][30] +
                  mat_A[1][22] * mat_B[22][30] +
                  mat_A[1][23] * mat_B[23][30] +
                  mat_A[1][24] * mat_B[24][30] +
                  mat_A[1][25] * mat_B[25][30] +
                  mat_A[1][26] * mat_B[26][30] +
                  mat_A[1][27] * mat_B[27][30] +
                  mat_A[1][28] * mat_B[28][30] +
                  mat_A[1][29] * mat_B[29][30] +
                  mat_A[1][30] * mat_B[30][30] +
                  mat_A[1][31] * mat_B[31][30];
    mat_C[1][31] <= 
                  mat_A[1][0] * mat_B[0][31] +
                  mat_A[1][1] * mat_B[1][31] +
                  mat_A[1][2] * mat_B[2][31] +
                  mat_A[1][3] * mat_B[3][31] +
                  mat_A[1][4] * mat_B[4][31] +
                  mat_A[1][5] * mat_B[5][31] +
                  mat_A[1][6] * mat_B[6][31] +
                  mat_A[1][7] * mat_B[7][31] +
                  mat_A[1][8] * mat_B[8][31] +
                  mat_A[1][9] * mat_B[9][31] +
                  mat_A[1][10] * mat_B[10][31] +
                  mat_A[1][11] * mat_B[11][31] +
                  mat_A[1][12] * mat_B[12][31] +
                  mat_A[1][13] * mat_B[13][31] +
                  mat_A[1][14] * mat_B[14][31] +
                  mat_A[1][15] * mat_B[15][31] +
                  mat_A[1][16] * mat_B[16][31] +
                  mat_A[1][17] * mat_B[17][31] +
                  mat_A[1][18] * mat_B[18][31] +
                  mat_A[1][19] * mat_B[19][31] +
                  mat_A[1][20] * mat_B[20][31] +
                  mat_A[1][21] * mat_B[21][31] +
                  mat_A[1][22] * mat_B[22][31] +
                  mat_A[1][23] * mat_B[23][31] +
                  mat_A[1][24] * mat_B[24][31] +
                  mat_A[1][25] * mat_B[25][31] +
                  mat_A[1][26] * mat_B[26][31] +
                  mat_A[1][27] * mat_B[27][31] +
                  mat_A[1][28] * mat_B[28][31] +
                  mat_A[1][29] * mat_B[29][31] +
                  mat_A[1][30] * mat_B[30][31] +
                  mat_A[1][31] * mat_B[31][31];
    mat_C[2][0] <= 
                  mat_A[2][0] * mat_B[0][0] +
                  mat_A[2][1] * mat_B[1][0] +
                  mat_A[2][2] * mat_B[2][0] +
                  mat_A[2][3] * mat_B[3][0] +
                  mat_A[2][4] * mat_B[4][0] +
                  mat_A[2][5] * mat_B[5][0] +
                  mat_A[2][6] * mat_B[6][0] +
                  mat_A[2][7] * mat_B[7][0] +
                  mat_A[2][8] * mat_B[8][0] +
                  mat_A[2][9] * mat_B[9][0] +
                  mat_A[2][10] * mat_B[10][0] +
                  mat_A[2][11] * mat_B[11][0] +
                  mat_A[2][12] * mat_B[12][0] +
                  mat_A[2][13] * mat_B[13][0] +
                  mat_A[2][14] * mat_B[14][0] +
                  mat_A[2][15] * mat_B[15][0] +
                  mat_A[2][16] * mat_B[16][0] +
                  mat_A[2][17] * mat_B[17][0] +
                  mat_A[2][18] * mat_B[18][0] +
                  mat_A[2][19] * mat_B[19][0] +
                  mat_A[2][20] * mat_B[20][0] +
                  mat_A[2][21] * mat_B[21][0] +
                  mat_A[2][22] * mat_B[22][0] +
                  mat_A[2][23] * mat_B[23][0] +
                  mat_A[2][24] * mat_B[24][0] +
                  mat_A[2][25] * mat_B[25][0] +
                  mat_A[2][26] * mat_B[26][0] +
                  mat_A[2][27] * mat_B[27][0] +
                  mat_A[2][28] * mat_B[28][0] +
                  mat_A[2][29] * mat_B[29][0] +
                  mat_A[2][30] * mat_B[30][0] +
                  mat_A[2][31] * mat_B[31][0];
    mat_C[2][1] <= 
                  mat_A[2][0] * mat_B[0][1] +
                  mat_A[2][1] * mat_B[1][1] +
                  mat_A[2][2] * mat_B[2][1] +
                  mat_A[2][3] * mat_B[3][1] +
                  mat_A[2][4] * mat_B[4][1] +
                  mat_A[2][5] * mat_B[5][1] +
                  mat_A[2][6] * mat_B[6][1] +
                  mat_A[2][7] * mat_B[7][1] +
                  mat_A[2][8] * mat_B[8][1] +
                  mat_A[2][9] * mat_B[9][1] +
                  mat_A[2][10] * mat_B[10][1] +
                  mat_A[2][11] * mat_B[11][1] +
                  mat_A[2][12] * mat_B[12][1] +
                  mat_A[2][13] * mat_B[13][1] +
                  mat_A[2][14] * mat_B[14][1] +
                  mat_A[2][15] * mat_B[15][1] +
                  mat_A[2][16] * mat_B[16][1] +
                  mat_A[2][17] * mat_B[17][1] +
                  mat_A[2][18] * mat_B[18][1] +
                  mat_A[2][19] * mat_B[19][1] +
                  mat_A[2][20] * mat_B[20][1] +
                  mat_A[2][21] * mat_B[21][1] +
                  mat_A[2][22] * mat_B[22][1] +
                  mat_A[2][23] * mat_B[23][1] +
                  mat_A[2][24] * mat_B[24][1] +
                  mat_A[2][25] * mat_B[25][1] +
                  mat_A[2][26] * mat_B[26][1] +
                  mat_A[2][27] * mat_B[27][1] +
                  mat_A[2][28] * mat_B[28][1] +
                  mat_A[2][29] * mat_B[29][1] +
                  mat_A[2][30] * mat_B[30][1] +
                  mat_A[2][31] * mat_B[31][1];
    mat_C[2][2] <= 
                  mat_A[2][0] * mat_B[0][2] +
                  mat_A[2][1] * mat_B[1][2] +
                  mat_A[2][2] * mat_B[2][2] +
                  mat_A[2][3] * mat_B[3][2] +
                  mat_A[2][4] * mat_B[4][2] +
                  mat_A[2][5] * mat_B[5][2] +
                  mat_A[2][6] * mat_B[6][2] +
                  mat_A[2][7] * mat_B[7][2] +
                  mat_A[2][8] * mat_B[8][2] +
                  mat_A[2][9] * mat_B[9][2] +
                  mat_A[2][10] * mat_B[10][2] +
                  mat_A[2][11] * mat_B[11][2] +
                  mat_A[2][12] * mat_B[12][2] +
                  mat_A[2][13] * mat_B[13][2] +
                  mat_A[2][14] * mat_B[14][2] +
                  mat_A[2][15] * mat_B[15][2] +
                  mat_A[2][16] * mat_B[16][2] +
                  mat_A[2][17] * mat_B[17][2] +
                  mat_A[2][18] * mat_B[18][2] +
                  mat_A[2][19] * mat_B[19][2] +
                  mat_A[2][20] * mat_B[20][2] +
                  mat_A[2][21] * mat_B[21][2] +
                  mat_A[2][22] * mat_B[22][2] +
                  mat_A[2][23] * mat_B[23][2] +
                  mat_A[2][24] * mat_B[24][2] +
                  mat_A[2][25] * mat_B[25][2] +
                  mat_A[2][26] * mat_B[26][2] +
                  mat_A[2][27] * mat_B[27][2] +
                  mat_A[2][28] * mat_B[28][2] +
                  mat_A[2][29] * mat_B[29][2] +
                  mat_A[2][30] * mat_B[30][2] +
                  mat_A[2][31] * mat_B[31][2];
    mat_C[2][3] <= 
                  mat_A[2][0] * mat_B[0][3] +
                  mat_A[2][1] * mat_B[1][3] +
                  mat_A[2][2] * mat_B[2][3] +
                  mat_A[2][3] * mat_B[3][3] +
                  mat_A[2][4] * mat_B[4][3] +
                  mat_A[2][5] * mat_B[5][3] +
                  mat_A[2][6] * mat_B[6][3] +
                  mat_A[2][7] * mat_B[7][3] +
                  mat_A[2][8] * mat_B[8][3] +
                  mat_A[2][9] * mat_B[9][3] +
                  mat_A[2][10] * mat_B[10][3] +
                  mat_A[2][11] * mat_B[11][3] +
                  mat_A[2][12] * mat_B[12][3] +
                  mat_A[2][13] * mat_B[13][3] +
                  mat_A[2][14] * mat_B[14][3] +
                  mat_A[2][15] * mat_B[15][3] +
                  mat_A[2][16] * mat_B[16][3] +
                  mat_A[2][17] * mat_B[17][3] +
                  mat_A[2][18] * mat_B[18][3] +
                  mat_A[2][19] * mat_B[19][3] +
                  mat_A[2][20] * mat_B[20][3] +
                  mat_A[2][21] * mat_B[21][3] +
                  mat_A[2][22] * mat_B[22][3] +
                  mat_A[2][23] * mat_B[23][3] +
                  mat_A[2][24] * mat_B[24][3] +
                  mat_A[2][25] * mat_B[25][3] +
                  mat_A[2][26] * mat_B[26][3] +
                  mat_A[2][27] * mat_B[27][3] +
                  mat_A[2][28] * mat_B[28][3] +
                  mat_A[2][29] * mat_B[29][3] +
                  mat_A[2][30] * mat_B[30][3] +
                  mat_A[2][31] * mat_B[31][3];
    mat_C[2][4] <= 
                  mat_A[2][0] * mat_B[0][4] +
                  mat_A[2][1] * mat_B[1][4] +
                  mat_A[2][2] * mat_B[2][4] +
                  mat_A[2][3] * mat_B[3][4] +
                  mat_A[2][4] * mat_B[4][4] +
                  mat_A[2][5] * mat_B[5][4] +
                  mat_A[2][6] * mat_B[6][4] +
                  mat_A[2][7] * mat_B[7][4] +
                  mat_A[2][8] * mat_B[8][4] +
                  mat_A[2][9] * mat_B[9][4] +
                  mat_A[2][10] * mat_B[10][4] +
                  mat_A[2][11] * mat_B[11][4] +
                  mat_A[2][12] * mat_B[12][4] +
                  mat_A[2][13] * mat_B[13][4] +
                  mat_A[2][14] * mat_B[14][4] +
                  mat_A[2][15] * mat_B[15][4] +
                  mat_A[2][16] * mat_B[16][4] +
                  mat_A[2][17] * mat_B[17][4] +
                  mat_A[2][18] * mat_B[18][4] +
                  mat_A[2][19] * mat_B[19][4] +
                  mat_A[2][20] * mat_B[20][4] +
                  mat_A[2][21] * mat_B[21][4] +
                  mat_A[2][22] * mat_B[22][4] +
                  mat_A[2][23] * mat_B[23][4] +
                  mat_A[2][24] * mat_B[24][4] +
                  mat_A[2][25] * mat_B[25][4] +
                  mat_A[2][26] * mat_B[26][4] +
                  mat_A[2][27] * mat_B[27][4] +
                  mat_A[2][28] * mat_B[28][4] +
                  mat_A[2][29] * mat_B[29][4] +
                  mat_A[2][30] * mat_B[30][4] +
                  mat_A[2][31] * mat_B[31][4];
    mat_C[2][5] <= 
                  mat_A[2][0] * mat_B[0][5] +
                  mat_A[2][1] * mat_B[1][5] +
                  mat_A[2][2] * mat_B[2][5] +
                  mat_A[2][3] * mat_B[3][5] +
                  mat_A[2][4] * mat_B[4][5] +
                  mat_A[2][5] * mat_B[5][5] +
                  mat_A[2][6] * mat_B[6][5] +
                  mat_A[2][7] * mat_B[7][5] +
                  mat_A[2][8] * mat_B[8][5] +
                  mat_A[2][9] * mat_B[9][5] +
                  mat_A[2][10] * mat_B[10][5] +
                  mat_A[2][11] * mat_B[11][5] +
                  mat_A[2][12] * mat_B[12][5] +
                  mat_A[2][13] * mat_B[13][5] +
                  mat_A[2][14] * mat_B[14][5] +
                  mat_A[2][15] * mat_B[15][5] +
                  mat_A[2][16] * mat_B[16][5] +
                  mat_A[2][17] * mat_B[17][5] +
                  mat_A[2][18] * mat_B[18][5] +
                  mat_A[2][19] * mat_B[19][5] +
                  mat_A[2][20] * mat_B[20][5] +
                  mat_A[2][21] * mat_B[21][5] +
                  mat_A[2][22] * mat_B[22][5] +
                  mat_A[2][23] * mat_B[23][5] +
                  mat_A[2][24] * mat_B[24][5] +
                  mat_A[2][25] * mat_B[25][5] +
                  mat_A[2][26] * mat_B[26][5] +
                  mat_A[2][27] * mat_B[27][5] +
                  mat_A[2][28] * mat_B[28][5] +
                  mat_A[2][29] * mat_B[29][5] +
                  mat_A[2][30] * mat_B[30][5] +
                  mat_A[2][31] * mat_B[31][5];
    mat_C[2][6] <= 
                  mat_A[2][0] * mat_B[0][6] +
                  mat_A[2][1] * mat_B[1][6] +
                  mat_A[2][2] * mat_B[2][6] +
                  mat_A[2][3] * mat_B[3][6] +
                  mat_A[2][4] * mat_B[4][6] +
                  mat_A[2][5] * mat_B[5][6] +
                  mat_A[2][6] * mat_B[6][6] +
                  mat_A[2][7] * mat_B[7][6] +
                  mat_A[2][8] * mat_B[8][6] +
                  mat_A[2][9] * mat_B[9][6] +
                  mat_A[2][10] * mat_B[10][6] +
                  mat_A[2][11] * mat_B[11][6] +
                  mat_A[2][12] * mat_B[12][6] +
                  mat_A[2][13] * mat_B[13][6] +
                  mat_A[2][14] * mat_B[14][6] +
                  mat_A[2][15] * mat_B[15][6] +
                  mat_A[2][16] * mat_B[16][6] +
                  mat_A[2][17] * mat_B[17][6] +
                  mat_A[2][18] * mat_B[18][6] +
                  mat_A[2][19] * mat_B[19][6] +
                  mat_A[2][20] * mat_B[20][6] +
                  mat_A[2][21] * mat_B[21][6] +
                  mat_A[2][22] * mat_B[22][6] +
                  mat_A[2][23] * mat_B[23][6] +
                  mat_A[2][24] * mat_B[24][6] +
                  mat_A[2][25] * mat_B[25][6] +
                  mat_A[2][26] * mat_B[26][6] +
                  mat_A[2][27] * mat_B[27][6] +
                  mat_A[2][28] * mat_B[28][6] +
                  mat_A[2][29] * mat_B[29][6] +
                  mat_A[2][30] * mat_B[30][6] +
                  mat_A[2][31] * mat_B[31][6];
    mat_C[2][7] <= 
                  mat_A[2][0] * mat_B[0][7] +
                  mat_A[2][1] * mat_B[1][7] +
                  mat_A[2][2] * mat_B[2][7] +
                  mat_A[2][3] * mat_B[3][7] +
                  mat_A[2][4] * mat_B[4][7] +
                  mat_A[2][5] * mat_B[5][7] +
                  mat_A[2][6] * mat_B[6][7] +
                  mat_A[2][7] * mat_B[7][7] +
                  mat_A[2][8] * mat_B[8][7] +
                  mat_A[2][9] * mat_B[9][7] +
                  mat_A[2][10] * mat_B[10][7] +
                  mat_A[2][11] * mat_B[11][7] +
                  mat_A[2][12] * mat_B[12][7] +
                  mat_A[2][13] * mat_B[13][7] +
                  mat_A[2][14] * mat_B[14][7] +
                  mat_A[2][15] * mat_B[15][7] +
                  mat_A[2][16] * mat_B[16][7] +
                  mat_A[2][17] * mat_B[17][7] +
                  mat_A[2][18] * mat_B[18][7] +
                  mat_A[2][19] * mat_B[19][7] +
                  mat_A[2][20] * mat_B[20][7] +
                  mat_A[2][21] * mat_B[21][7] +
                  mat_A[2][22] * mat_B[22][7] +
                  mat_A[2][23] * mat_B[23][7] +
                  mat_A[2][24] * mat_B[24][7] +
                  mat_A[2][25] * mat_B[25][7] +
                  mat_A[2][26] * mat_B[26][7] +
                  mat_A[2][27] * mat_B[27][7] +
                  mat_A[2][28] * mat_B[28][7] +
                  mat_A[2][29] * mat_B[29][7] +
                  mat_A[2][30] * mat_B[30][7] +
                  mat_A[2][31] * mat_B[31][7];
    mat_C[2][8] <= 
                  mat_A[2][0] * mat_B[0][8] +
                  mat_A[2][1] * mat_B[1][8] +
                  mat_A[2][2] * mat_B[2][8] +
                  mat_A[2][3] * mat_B[3][8] +
                  mat_A[2][4] * mat_B[4][8] +
                  mat_A[2][5] * mat_B[5][8] +
                  mat_A[2][6] * mat_B[6][8] +
                  mat_A[2][7] * mat_B[7][8] +
                  mat_A[2][8] * mat_B[8][8] +
                  mat_A[2][9] * mat_B[9][8] +
                  mat_A[2][10] * mat_B[10][8] +
                  mat_A[2][11] * mat_B[11][8] +
                  mat_A[2][12] * mat_B[12][8] +
                  mat_A[2][13] * mat_B[13][8] +
                  mat_A[2][14] * mat_B[14][8] +
                  mat_A[2][15] * mat_B[15][8] +
                  mat_A[2][16] * mat_B[16][8] +
                  mat_A[2][17] * mat_B[17][8] +
                  mat_A[2][18] * mat_B[18][8] +
                  mat_A[2][19] * mat_B[19][8] +
                  mat_A[2][20] * mat_B[20][8] +
                  mat_A[2][21] * mat_B[21][8] +
                  mat_A[2][22] * mat_B[22][8] +
                  mat_A[2][23] * mat_B[23][8] +
                  mat_A[2][24] * mat_B[24][8] +
                  mat_A[2][25] * mat_B[25][8] +
                  mat_A[2][26] * mat_B[26][8] +
                  mat_A[2][27] * mat_B[27][8] +
                  mat_A[2][28] * mat_B[28][8] +
                  mat_A[2][29] * mat_B[29][8] +
                  mat_A[2][30] * mat_B[30][8] +
                  mat_A[2][31] * mat_B[31][8];
    mat_C[2][9] <= 
                  mat_A[2][0] * mat_B[0][9] +
                  mat_A[2][1] * mat_B[1][9] +
                  mat_A[2][2] * mat_B[2][9] +
                  mat_A[2][3] * mat_B[3][9] +
                  mat_A[2][4] * mat_B[4][9] +
                  mat_A[2][5] * mat_B[5][9] +
                  mat_A[2][6] * mat_B[6][9] +
                  mat_A[2][7] * mat_B[7][9] +
                  mat_A[2][8] * mat_B[8][9] +
                  mat_A[2][9] * mat_B[9][9] +
                  mat_A[2][10] * mat_B[10][9] +
                  mat_A[2][11] * mat_B[11][9] +
                  mat_A[2][12] * mat_B[12][9] +
                  mat_A[2][13] * mat_B[13][9] +
                  mat_A[2][14] * mat_B[14][9] +
                  mat_A[2][15] * mat_B[15][9] +
                  mat_A[2][16] * mat_B[16][9] +
                  mat_A[2][17] * mat_B[17][9] +
                  mat_A[2][18] * mat_B[18][9] +
                  mat_A[2][19] * mat_B[19][9] +
                  mat_A[2][20] * mat_B[20][9] +
                  mat_A[2][21] * mat_B[21][9] +
                  mat_A[2][22] * mat_B[22][9] +
                  mat_A[2][23] * mat_B[23][9] +
                  mat_A[2][24] * mat_B[24][9] +
                  mat_A[2][25] * mat_B[25][9] +
                  mat_A[2][26] * mat_B[26][9] +
                  mat_A[2][27] * mat_B[27][9] +
                  mat_A[2][28] * mat_B[28][9] +
                  mat_A[2][29] * mat_B[29][9] +
                  mat_A[2][30] * mat_B[30][9] +
                  mat_A[2][31] * mat_B[31][9];
    mat_C[2][10] <= 
                  mat_A[2][0] * mat_B[0][10] +
                  mat_A[2][1] * mat_B[1][10] +
                  mat_A[2][2] * mat_B[2][10] +
                  mat_A[2][3] * mat_B[3][10] +
                  mat_A[2][4] * mat_B[4][10] +
                  mat_A[2][5] * mat_B[5][10] +
                  mat_A[2][6] * mat_B[6][10] +
                  mat_A[2][7] * mat_B[7][10] +
                  mat_A[2][8] * mat_B[8][10] +
                  mat_A[2][9] * mat_B[9][10] +
                  mat_A[2][10] * mat_B[10][10] +
                  mat_A[2][11] * mat_B[11][10] +
                  mat_A[2][12] * mat_B[12][10] +
                  mat_A[2][13] * mat_B[13][10] +
                  mat_A[2][14] * mat_B[14][10] +
                  mat_A[2][15] * mat_B[15][10] +
                  mat_A[2][16] * mat_B[16][10] +
                  mat_A[2][17] * mat_B[17][10] +
                  mat_A[2][18] * mat_B[18][10] +
                  mat_A[2][19] * mat_B[19][10] +
                  mat_A[2][20] * mat_B[20][10] +
                  mat_A[2][21] * mat_B[21][10] +
                  mat_A[2][22] * mat_B[22][10] +
                  mat_A[2][23] * mat_B[23][10] +
                  mat_A[2][24] * mat_B[24][10] +
                  mat_A[2][25] * mat_B[25][10] +
                  mat_A[2][26] * mat_B[26][10] +
                  mat_A[2][27] * mat_B[27][10] +
                  mat_A[2][28] * mat_B[28][10] +
                  mat_A[2][29] * mat_B[29][10] +
                  mat_A[2][30] * mat_B[30][10] +
                  mat_A[2][31] * mat_B[31][10];
    mat_C[2][11] <= 
                  mat_A[2][0] * mat_B[0][11] +
                  mat_A[2][1] * mat_B[1][11] +
                  mat_A[2][2] * mat_B[2][11] +
                  mat_A[2][3] * mat_B[3][11] +
                  mat_A[2][4] * mat_B[4][11] +
                  mat_A[2][5] * mat_B[5][11] +
                  mat_A[2][6] * mat_B[6][11] +
                  mat_A[2][7] * mat_B[7][11] +
                  mat_A[2][8] * mat_B[8][11] +
                  mat_A[2][9] * mat_B[9][11] +
                  mat_A[2][10] * mat_B[10][11] +
                  mat_A[2][11] * mat_B[11][11] +
                  mat_A[2][12] * mat_B[12][11] +
                  mat_A[2][13] * mat_B[13][11] +
                  mat_A[2][14] * mat_B[14][11] +
                  mat_A[2][15] * mat_B[15][11] +
                  mat_A[2][16] * mat_B[16][11] +
                  mat_A[2][17] * mat_B[17][11] +
                  mat_A[2][18] * mat_B[18][11] +
                  mat_A[2][19] * mat_B[19][11] +
                  mat_A[2][20] * mat_B[20][11] +
                  mat_A[2][21] * mat_B[21][11] +
                  mat_A[2][22] * mat_B[22][11] +
                  mat_A[2][23] * mat_B[23][11] +
                  mat_A[2][24] * mat_B[24][11] +
                  mat_A[2][25] * mat_B[25][11] +
                  mat_A[2][26] * mat_B[26][11] +
                  mat_A[2][27] * mat_B[27][11] +
                  mat_A[2][28] * mat_B[28][11] +
                  mat_A[2][29] * mat_B[29][11] +
                  mat_A[2][30] * mat_B[30][11] +
                  mat_A[2][31] * mat_B[31][11];
    mat_C[2][12] <= 
                  mat_A[2][0] * mat_B[0][12] +
                  mat_A[2][1] * mat_B[1][12] +
                  mat_A[2][2] * mat_B[2][12] +
                  mat_A[2][3] * mat_B[3][12] +
                  mat_A[2][4] * mat_B[4][12] +
                  mat_A[2][5] * mat_B[5][12] +
                  mat_A[2][6] * mat_B[6][12] +
                  mat_A[2][7] * mat_B[7][12] +
                  mat_A[2][8] * mat_B[8][12] +
                  mat_A[2][9] * mat_B[9][12] +
                  mat_A[2][10] * mat_B[10][12] +
                  mat_A[2][11] * mat_B[11][12] +
                  mat_A[2][12] * mat_B[12][12] +
                  mat_A[2][13] * mat_B[13][12] +
                  mat_A[2][14] * mat_B[14][12] +
                  mat_A[2][15] * mat_B[15][12] +
                  mat_A[2][16] * mat_B[16][12] +
                  mat_A[2][17] * mat_B[17][12] +
                  mat_A[2][18] * mat_B[18][12] +
                  mat_A[2][19] * mat_B[19][12] +
                  mat_A[2][20] * mat_B[20][12] +
                  mat_A[2][21] * mat_B[21][12] +
                  mat_A[2][22] * mat_B[22][12] +
                  mat_A[2][23] * mat_B[23][12] +
                  mat_A[2][24] * mat_B[24][12] +
                  mat_A[2][25] * mat_B[25][12] +
                  mat_A[2][26] * mat_B[26][12] +
                  mat_A[2][27] * mat_B[27][12] +
                  mat_A[2][28] * mat_B[28][12] +
                  mat_A[2][29] * mat_B[29][12] +
                  mat_A[2][30] * mat_B[30][12] +
                  mat_A[2][31] * mat_B[31][12];
    mat_C[2][13] <= 
                  mat_A[2][0] * mat_B[0][13] +
                  mat_A[2][1] * mat_B[1][13] +
                  mat_A[2][2] * mat_B[2][13] +
                  mat_A[2][3] * mat_B[3][13] +
                  mat_A[2][4] * mat_B[4][13] +
                  mat_A[2][5] * mat_B[5][13] +
                  mat_A[2][6] * mat_B[6][13] +
                  mat_A[2][7] * mat_B[7][13] +
                  mat_A[2][8] * mat_B[8][13] +
                  mat_A[2][9] * mat_B[9][13] +
                  mat_A[2][10] * mat_B[10][13] +
                  mat_A[2][11] * mat_B[11][13] +
                  mat_A[2][12] * mat_B[12][13] +
                  mat_A[2][13] * mat_B[13][13] +
                  mat_A[2][14] * mat_B[14][13] +
                  mat_A[2][15] * mat_B[15][13] +
                  mat_A[2][16] * mat_B[16][13] +
                  mat_A[2][17] * mat_B[17][13] +
                  mat_A[2][18] * mat_B[18][13] +
                  mat_A[2][19] * mat_B[19][13] +
                  mat_A[2][20] * mat_B[20][13] +
                  mat_A[2][21] * mat_B[21][13] +
                  mat_A[2][22] * mat_B[22][13] +
                  mat_A[2][23] * mat_B[23][13] +
                  mat_A[2][24] * mat_B[24][13] +
                  mat_A[2][25] * mat_B[25][13] +
                  mat_A[2][26] * mat_B[26][13] +
                  mat_A[2][27] * mat_B[27][13] +
                  mat_A[2][28] * mat_B[28][13] +
                  mat_A[2][29] * mat_B[29][13] +
                  mat_A[2][30] * mat_B[30][13] +
                  mat_A[2][31] * mat_B[31][13];
    mat_C[2][14] <= 
                  mat_A[2][0] * mat_B[0][14] +
                  mat_A[2][1] * mat_B[1][14] +
                  mat_A[2][2] * mat_B[2][14] +
                  mat_A[2][3] * mat_B[3][14] +
                  mat_A[2][4] * mat_B[4][14] +
                  mat_A[2][5] * mat_B[5][14] +
                  mat_A[2][6] * mat_B[6][14] +
                  mat_A[2][7] * mat_B[7][14] +
                  mat_A[2][8] * mat_B[8][14] +
                  mat_A[2][9] * mat_B[9][14] +
                  mat_A[2][10] * mat_B[10][14] +
                  mat_A[2][11] * mat_B[11][14] +
                  mat_A[2][12] * mat_B[12][14] +
                  mat_A[2][13] * mat_B[13][14] +
                  mat_A[2][14] * mat_B[14][14] +
                  mat_A[2][15] * mat_B[15][14] +
                  mat_A[2][16] * mat_B[16][14] +
                  mat_A[2][17] * mat_B[17][14] +
                  mat_A[2][18] * mat_B[18][14] +
                  mat_A[2][19] * mat_B[19][14] +
                  mat_A[2][20] * mat_B[20][14] +
                  mat_A[2][21] * mat_B[21][14] +
                  mat_A[2][22] * mat_B[22][14] +
                  mat_A[2][23] * mat_B[23][14] +
                  mat_A[2][24] * mat_B[24][14] +
                  mat_A[2][25] * mat_B[25][14] +
                  mat_A[2][26] * mat_B[26][14] +
                  mat_A[2][27] * mat_B[27][14] +
                  mat_A[2][28] * mat_B[28][14] +
                  mat_A[2][29] * mat_B[29][14] +
                  mat_A[2][30] * mat_B[30][14] +
                  mat_A[2][31] * mat_B[31][14];
    mat_C[2][15] <= 
                  mat_A[2][0] * mat_B[0][15] +
                  mat_A[2][1] * mat_B[1][15] +
                  mat_A[2][2] * mat_B[2][15] +
                  mat_A[2][3] * mat_B[3][15] +
                  mat_A[2][4] * mat_B[4][15] +
                  mat_A[2][5] * mat_B[5][15] +
                  mat_A[2][6] * mat_B[6][15] +
                  mat_A[2][7] * mat_B[7][15] +
                  mat_A[2][8] * mat_B[8][15] +
                  mat_A[2][9] * mat_B[9][15] +
                  mat_A[2][10] * mat_B[10][15] +
                  mat_A[2][11] * mat_B[11][15] +
                  mat_A[2][12] * mat_B[12][15] +
                  mat_A[2][13] * mat_B[13][15] +
                  mat_A[2][14] * mat_B[14][15] +
                  mat_A[2][15] * mat_B[15][15] +
                  mat_A[2][16] * mat_B[16][15] +
                  mat_A[2][17] * mat_B[17][15] +
                  mat_A[2][18] * mat_B[18][15] +
                  mat_A[2][19] * mat_B[19][15] +
                  mat_A[2][20] * mat_B[20][15] +
                  mat_A[2][21] * mat_B[21][15] +
                  mat_A[2][22] * mat_B[22][15] +
                  mat_A[2][23] * mat_B[23][15] +
                  mat_A[2][24] * mat_B[24][15] +
                  mat_A[2][25] * mat_B[25][15] +
                  mat_A[2][26] * mat_B[26][15] +
                  mat_A[2][27] * mat_B[27][15] +
                  mat_A[2][28] * mat_B[28][15] +
                  mat_A[2][29] * mat_B[29][15] +
                  mat_A[2][30] * mat_B[30][15] +
                  mat_A[2][31] * mat_B[31][15];
    mat_C[2][16] <= 
                  mat_A[2][0] * mat_B[0][16] +
                  mat_A[2][1] * mat_B[1][16] +
                  mat_A[2][2] * mat_B[2][16] +
                  mat_A[2][3] * mat_B[3][16] +
                  mat_A[2][4] * mat_B[4][16] +
                  mat_A[2][5] * mat_B[5][16] +
                  mat_A[2][6] * mat_B[6][16] +
                  mat_A[2][7] * mat_B[7][16] +
                  mat_A[2][8] * mat_B[8][16] +
                  mat_A[2][9] * mat_B[9][16] +
                  mat_A[2][10] * mat_B[10][16] +
                  mat_A[2][11] * mat_B[11][16] +
                  mat_A[2][12] * mat_B[12][16] +
                  mat_A[2][13] * mat_B[13][16] +
                  mat_A[2][14] * mat_B[14][16] +
                  mat_A[2][15] * mat_B[15][16] +
                  mat_A[2][16] * mat_B[16][16] +
                  mat_A[2][17] * mat_B[17][16] +
                  mat_A[2][18] * mat_B[18][16] +
                  mat_A[2][19] * mat_B[19][16] +
                  mat_A[2][20] * mat_B[20][16] +
                  mat_A[2][21] * mat_B[21][16] +
                  mat_A[2][22] * mat_B[22][16] +
                  mat_A[2][23] * mat_B[23][16] +
                  mat_A[2][24] * mat_B[24][16] +
                  mat_A[2][25] * mat_B[25][16] +
                  mat_A[2][26] * mat_B[26][16] +
                  mat_A[2][27] * mat_B[27][16] +
                  mat_A[2][28] * mat_B[28][16] +
                  mat_A[2][29] * mat_B[29][16] +
                  mat_A[2][30] * mat_B[30][16] +
                  mat_A[2][31] * mat_B[31][16];
    mat_C[2][17] <= 
                  mat_A[2][0] * mat_B[0][17] +
                  mat_A[2][1] * mat_B[1][17] +
                  mat_A[2][2] * mat_B[2][17] +
                  mat_A[2][3] * mat_B[3][17] +
                  mat_A[2][4] * mat_B[4][17] +
                  mat_A[2][5] * mat_B[5][17] +
                  mat_A[2][6] * mat_B[6][17] +
                  mat_A[2][7] * mat_B[7][17] +
                  mat_A[2][8] * mat_B[8][17] +
                  mat_A[2][9] * mat_B[9][17] +
                  mat_A[2][10] * mat_B[10][17] +
                  mat_A[2][11] * mat_B[11][17] +
                  mat_A[2][12] * mat_B[12][17] +
                  mat_A[2][13] * mat_B[13][17] +
                  mat_A[2][14] * mat_B[14][17] +
                  mat_A[2][15] * mat_B[15][17] +
                  mat_A[2][16] * mat_B[16][17] +
                  mat_A[2][17] * mat_B[17][17] +
                  mat_A[2][18] * mat_B[18][17] +
                  mat_A[2][19] * mat_B[19][17] +
                  mat_A[2][20] * mat_B[20][17] +
                  mat_A[2][21] * mat_B[21][17] +
                  mat_A[2][22] * mat_B[22][17] +
                  mat_A[2][23] * mat_B[23][17] +
                  mat_A[2][24] * mat_B[24][17] +
                  mat_A[2][25] * mat_B[25][17] +
                  mat_A[2][26] * mat_B[26][17] +
                  mat_A[2][27] * mat_B[27][17] +
                  mat_A[2][28] * mat_B[28][17] +
                  mat_A[2][29] * mat_B[29][17] +
                  mat_A[2][30] * mat_B[30][17] +
                  mat_A[2][31] * mat_B[31][17];
    mat_C[2][18] <= 
                  mat_A[2][0] * mat_B[0][18] +
                  mat_A[2][1] * mat_B[1][18] +
                  mat_A[2][2] * mat_B[2][18] +
                  mat_A[2][3] * mat_B[3][18] +
                  mat_A[2][4] * mat_B[4][18] +
                  mat_A[2][5] * mat_B[5][18] +
                  mat_A[2][6] * mat_B[6][18] +
                  mat_A[2][7] * mat_B[7][18] +
                  mat_A[2][8] * mat_B[8][18] +
                  mat_A[2][9] * mat_B[9][18] +
                  mat_A[2][10] * mat_B[10][18] +
                  mat_A[2][11] * mat_B[11][18] +
                  mat_A[2][12] * mat_B[12][18] +
                  mat_A[2][13] * mat_B[13][18] +
                  mat_A[2][14] * mat_B[14][18] +
                  mat_A[2][15] * mat_B[15][18] +
                  mat_A[2][16] * mat_B[16][18] +
                  mat_A[2][17] * mat_B[17][18] +
                  mat_A[2][18] * mat_B[18][18] +
                  mat_A[2][19] * mat_B[19][18] +
                  mat_A[2][20] * mat_B[20][18] +
                  mat_A[2][21] * mat_B[21][18] +
                  mat_A[2][22] * mat_B[22][18] +
                  mat_A[2][23] * mat_B[23][18] +
                  mat_A[2][24] * mat_B[24][18] +
                  mat_A[2][25] * mat_B[25][18] +
                  mat_A[2][26] * mat_B[26][18] +
                  mat_A[2][27] * mat_B[27][18] +
                  mat_A[2][28] * mat_B[28][18] +
                  mat_A[2][29] * mat_B[29][18] +
                  mat_A[2][30] * mat_B[30][18] +
                  mat_A[2][31] * mat_B[31][18];
    mat_C[2][19] <= 
                  mat_A[2][0] * mat_B[0][19] +
                  mat_A[2][1] * mat_B[1][19] +
                  mat_A[2][2] * mat_B[2][19] +
                  mat_A[2][3] * mat_B[3][19] +
                  mat_A[2][4] * mat_B[4][19] +
                  mat_A[2][5] * mat_B[5][19] +
                  mat_A[2][6] * mat_B[6][19] +
                  mat_A[2][7] * mat_B[7][19] +
                  mat_A[2][8] * mat_B[8][19] +
                  mat_A[2][9] * mat_B[9][19] +
                  mat_A[2][10] * mat_B[10][19] +
                  mat_A[2][11] * mat_B[11][19] +
                  mat_A[2][12] * mat_B[12][19] +
                  mat_A[2][13] * mat_B[13][19] +
                  mat_A[2][14] * mat_B[14][19] +
                  mat_A[2][15] * mat_B[15][19] +
                  mat_A[2][16] * mat_B[16][19] +
                  mat_A[2][17] * mat_B[17][19] +
                  mat_A[2][18] * mat_B[18][19] +
                  mat_A[2][19] * mat_B[19][19] +
                  mat_A[2][20] * mat_B[20][19] +
                  mat_A[2][21] * mat_B[21][19] +
                  mat_A[2][22] * mat_B[22][19] +
                  mat_A[2][23] * mat_B[23][19] +
                  mat_A[2][24] * mat_B[24][19] +
                  mat_A[2][25] * mat_B[25][19] +
                  mat_A[2][26] * mat_B[26][19] +
                  mat_A[2][27] * mat_B[27][19] +
                  mat_A[2][28] * mat_B[28][19] +
                  mat_A[2][29] * mat_B[29][19] +
                  mat_A[2][30] * mat_B[30][19] +
                  mat_A[2][31] * mat_B[31][19];
    mat_C[2][20] <= 
                  mat_A[2][0] * mat_B[0][20] +
                  mat_A[2][1] * mat_B[1][20] +
                  mat_A[2][2] * mat_B[2][20] +
                  mat_A[2][3] * mat_B[3][20] +
                  mat_A[2][4] * mat_B[4][20] +
                  mat_A[2][5] * mat_B[5][20] +
                  mat_A[2][6] * mat_B[6][20] +
                  mat_A[2][7] * mat_B[7][20] +
                  mat_A[2][8] * mat_B[8][20] +
                  mat_A[2][9] * mat_B[9][20] +
                  mat_A[2][10] * mat_B[10][20] +
                  mat_A[2][11] * mat_B[11][20] +
                  mat_A[2][12] * mat_B[12][20] +
                  mat_A[2][13] * mat_B[13][20] +
                  mat_A[2][14] * mat_B[14][20] +
                  mat_A[2][15] * mat_B[15][20] +
                  mat_A[2][16] * mat_B[16][20] +
                  mat_A[2][17] * mat_B[17][20] +
                  mat_A[2][18] * mat_B[18][20] +
                  mat_A[2][19] * mat_B[19][20] +
                  mat_A[2][20] * mat_B[20][20] +
                  mat_A[2][21] * mat_B[21][20] +
                  mat_A[2][22] * mat_B[22][20] +
                  mat_A[2][23] * mat_B[23][20] +
                  mat_A[2][24] * mat_B[24][20] +
                  mat_A[2][25] * mat_B[25][20] +
                  mat_A[2][26] * mat_B[26][20] +
                  mat_A[2][27] * mat_B[27][20] +
                  mat_A[2][28] * mat_B[28][20] +
                  mat_A[2][29] * mat_B[29][20] +
                  mat_A[2][30] * mat_B[30][20] +
                  mat_A[2][31] * mat_B[31][20];
    mat_C[2][21] <= 
                  mat_A[2][0] * mat_B[0][21] +
                  mat_A[2][1] * mat_B[1][21] +
                  mat_A[2][2] * mat_B[2][21] +
                  mat_A[2][3] * mat_B[3][21] +
                  mat_A[2][4] * mat_B[4][21] +
                  mat_A[2][5] * mat_B[5][21] +
                  mat_A[2][6] * mat_B[6][21] +
                  mat_A[2][7] * mat_B[7][21] +
                  mat_A[2][8] * mat_B[8][21] +
                  mat_A[2][9] * mat_B[9][21] +
                  mat_A[2][10] * mat_B[10][21] +
                  mat_A[2][11] * mat_B[11][21] +
                  mat_A[2][12] * mat_B[12][21] +
                  mat_A[2][13] * mat_B[13][21] +
                  mat_A[2][14] * mat_B[14][21] +
                  mat_A[2][15] * mat_B[15][21] +
                  mat_A[2][16] * mat_B[16][21] +
                  mat_A[2][17] * mat_B[17][21] +
                  mat_A[2][18] * mat_B[18][21] +
                  mat_A[2][19] * mat_B[19][21] +
                  mat_A[2][20] * mat_B[20][21] +
                  mat_A[2][21] * mat_B[21][21] +
                  mat_A[2][22] * mat_B[22][21] +
                  mat_A[2][23] * mat_B[23][21] +
                  mat_A[2][24] * mat_B[24][21] +
                  mat_A[2][25] * mat_B[25][21] +
                  mat_A[2][26] * mat_B[26][21] +
                  mat_A[2][27] * mat_B[27][21] +
                  mat_A[2][28] * mat_B[28][21] +
                  mat_A[2][29] * mat_B[29][21] +
                  mat_A[2][30] * mat_B[30][21] +
                  mat_A[2][31] * mat_B[31][21];
    mat_C[2][22] <= 
                  mat_A[2][0] * mat_B[0][22] +
                  mat_A[2][1] * mat_B[1][22] +
                  mat_A[2][2] * mat_B[2][22] +
                  mat_A[2][3] * mat_B[3][22] +
                  mat_A[2][4] * mat_B[4][22] +
                  mat_A[2][5] * mat_B[5][22] +
                  mat_A[2][6] * mat_B[6][22] +
                  mat_A[2][7] * mat_B[7][22] +
                  mat_A[2][8] * mat_B[8][22] +
                  mat_A[2][9] * mat_B[9][22] +
                  mat_A[2][10] * mat_B[10][22] +
                  mat_A[2][11] * mat_B[11][22] +
                  mat_A[2][12] * mat_B[12][22] +
                  mat_A[2][13] * mat_B[13][22] +
                  mat_A[2][14] * mat_B[14][22] +
                  mat_A[2][15] * mat_B[15][22] +
                  mat_A[2][16] * mat_B[16][22] +
                  mat_A[2][17] * mat_B[17][22] +
                  mat_A[2][18] * mat_B[18][22] +
                  mat_A[2][19] * mat_B[19][22] +
                  mat_A[2][20] * mat_B[20][22] +
                  mat_A[2][21] * mat_B[21][22] +
                  mat_A[2][22] * mat_B[22][22] +
                  mat_A[2][23] * mat_B[23][22] +
                  mat_A[2][24] * mat_B[24][22] +
                  mat_A[2][25] * mat_B[25][22] +
                  mat_A[2][26] * mat_B[26][22] +
                  mat_A[2][27] * mat_B[27][22] +
                  mat_A[2][28] * mat_B[28][22] +
                  mat_A[2][29] * mat_B[29][22] +
                  mat_A[2][30] * mat_B[30][22] +
                  mat_A[2][31] * mat_B[31][22];
    mat_C[2][23] <= 
                  mat_A[2][0] * mat_B[0][23] +
                  mat_A[2][1] * mat_B[1][23] +
                  mat_A[2][2] * mat_B[2][23] +
                  mat_A[2][3] * mat_B[3][23] +
                  mat_A[2][4] * mat_B[4][23] +
                  mat_A[2][5] * mat_B[5][23] +
                  mat_A[2][6] * mat_B[6][23] +
                  mat_A[2][7] * mat_B[7][23] +
                  mat_A[2][8] * mat_B[8][23] +
                  mat_A[2][9] * mat_B[9][23] +
                  mat_A[2][10] * mat_B[10][23] +
                  mat_A[2][11] * mat_B[11][23] +
                  mat_A[2][12] * mat_B[12][23] +
                  mat_A[2][13] * mat_B[13][23] +
                  mat_A[2][14] * mat_B[14][23] +
                  mat_A[2][15] * mat_B[15][23] +
                  mat_A[2][16] * mat_B[16][23] +
                  mat_A[2][17] * mat_B[17][23] +
                  mat_A[2][18] * mat_B[18][23] +
                  mat_A[2][19] * mat_B[19][23] +
                  mat_A[2][20] * mat_B[20][23] +
                  mat_A[2][21] * mat_B[21][23] +
                  mat_A[2][22] * mat_B[22][23] +
                  mat_A[2][23] * mat_B[23][23] +
                  mat_A[2][24] * mat_B[24][23] +
                  mat_A[2][25] * mat_B[25][23] +
                  mat_A[2][26] * mat_B[26][23] +
                  mat_A[2][27] * mat_B[27][23] +
                  mat_A[2][28] * mat_B[28][23] +
                  mat_A[2][29] * mat_B[29][23] +
                  mat_A[2][30] * mat_B[30][23] +
                  mat_A[2][31] * mat_B[31][23];
    mat_C[2][24] <= 
                  mat_A[2][0] * mat_B[0][24] +
                  mat_A[2][1] * mat_B[1][24] +
                  mat_A[2][2] * mat_B[2][24] +
                  mat_A[2][3] * mat_B[3][24] +
                  mat_A[2][4] * mat_B[4][24] +
                  mat_A[2][5] * mat_B[5][24] +
                  mat_A[2][6] * mat_B[6][24] +
                  mat_A[2][7] * mat_B[7][24] +
                  mat_A[2][8] * mat_B[8][24] +
                  mat_A[2][9] * mat_B[9][24] +
                  mat_A[2][10] * mat_B[10][24] +
                  mat_A[2][11] * mat_B[11][24] +
                  mat_A[2][12] * mat_B[12][24] +
                  mat_A[2][13] * mat_B[13][24] +
                  mat_A[2][14] * mat_B[14][24] +
                  mat_A[2][15] * mat_B[15][24] +
                  mat_A[2][16] * mat_B[16][24] +
                  mat_A[2][17] * mat_B[17][24] +
                  mat_A[2][18] * mat_B[18][24] +
                  mat_A[2][19] * mat_B[19][24] +
                  mat_A[2][20] * mat_B[20][24] +
                  mat_A[2][21] * mat_B[21][24] +
                  mat_A[2][22] * mat_B[22][24] +
                  mat_A[2][23] * mat_B[23][24] +
                  mat_A[2][24] * mat_B[24][24] +
                  mat_A[2][25] * mat_B[25][24] +
                  mat_A[2][26] * mat_B[26][24] +
                  mat_A[2][27] * mat_B[27][24] +
                  mat_A[2][28] * mat_B[28][24] +
                  mat_A[2][29] * mat_B[29][24] +
                  mat_A[2][30] * mat_B[30][24] +
                  mat_A[2][31] * mat_B[31][24];
    mat_C[2][25] <= 
                  mat_A[2][0] * mat_B[0][25] +
                  mat_A[2][1] * mat_B[1][25] +
                  mat_A[2][2] * mat_B[2][25] +
                  mat_A[2][3] * mat_B[3][25] +
                  mat_A[2][4] * mat_B[4][25] +
                  mat_A[2][5] * mat_B[5][25] +
                  mat_A[2][6] * mat_B[6][25] +
                  mat_A[2][7] * mat_B[7][25] +
                  mat_A[2][8] * mat_B[8][25] +
                  mat_A[2][9] * mat_B[9][25] +
                  mat_A[2][10] * mat_B[10][25] +
                  mat_A[2][11] * mat_B[11][25] +
                  mat_A[2][12] * mat_B[12][25] +
                  mat_A[2][13] * mat_B[13][25] +
                  mat_A[2][14] * mat_B[14][25] +
                  mat_A[2][15] * mat_B[15][25] +
                  mat_A[2][16] * mat_B[16][25] +
                  mat_A[2][17] * mat_B[17][25] +
                  mat_A[2][18] * mat_B[18][25] +
                  mat_A[2][19] * mat_B[19][25] +
                  mat_A[2][20] * mat_B[20][25] +
                  mat_A[2][21] * mat_B[21][25] +
                  mat_A[2][22] * mat_B[22][25] +
                  mat_A[2][23] * mat_B[23][25] +
                  mat_A[2][24] * mat_B[24][25] +
                  mat_A[2][25] * mat_B[25][25] +
                  mat_A[2][26] * mat_B[26][25] +
                  mat_A[2][27] * mat_B[27][25] +
                  mat_A[2][28] * mat_B[28][25] +
                  mat_A[2][29] * mat_B[29][25] +
                  mat_A[2][30] * mat_B[30][25] +
                  mat_A[2][31] * mat_B[31][25];
    mat_C[2][26] <= 
                  mat_A[2][0] * mat_B[0][26] +
                  mat_A[2][1] * mat_B[1][26] +
                  mat_A[2][2] * mat_B[2][26] +
                  mat_A[2][3] * mat_B[3][26] +
                  mat_A[2][4] * mat_B[4][26] +
                  mat_A[2][5] * mat_B[5][26] +
                  mat_A[2][6] * mat_B[6][26] +
                  mat_A[2][7] * mat_B[7][26] +
                  mat_A[2][8] * mat_B[8][26] +
                  mat_A[2][9] * mat_B[9][26] +
                  mat_A[2][10] * mat_B[10][26] +
                  mat_A[2][11] * mat_B[11][26] +
                  mat_A[2][12] * mat_B[12][26] +
                  mat_A[2][13] * mat_B[13][26] +
                  mat_A[2][14] * mat_B[14][26] +
                  mat_A[2][15] * mat_B[15][26] +
                  mat_A[2][16] * mat_B[16][26] +
                  mat_A[2][17] * mat_B[17][26] +
                  mat_A[2][18] * mat_B[18][26] +
                  mat_A[2][19] * mat_B[19][26] +
                  mat_A[2][20] * mat_B[20][26] +
                  mat_A[2][21] * mat_B[21][26] +
                  mat_A[2][22] * mat_B[22][26] +
                  mat_A[2][23] * mat_B[23][26] +
                  mat_A[2][24] * mat_B[24][26] +
                  mat_A[2][25] * mat_B[25][26] +
                  mat_A[2][26] * mat_B[26][26] +
                  mat_A[2][27] * mat_B[27][26] +
                  mat_A[2][28] * mat_B[28][26] +
                  mat_A[2][29] * mat_B[29][26] +
                  mat_A[2][30] * mat_B[30][26] +
                  mat_A[2][31] * mat_B[31][26];
    mat_C[2][27] <= 
                  mat_A[2][0] * mat_B[0][27] +
                  mat_A[2][1] * mat_B[1][27] +
                  mat_A[2][2] * mat_B[2][27] +
                  mat_A[2][3] * mat_B[3][27] +
                  mat_A[2][4] * mat_B[4][27] +
                  mat_A[2][5] * mat_B[5][27] +
                  mat_A[2][6] * mat_B[6][27] +
                  mat_A[2][7] * mat_B[7][27] +
                  mat_A[2][8] * mat_B[8][27] +
                  mat_A[2][9] * mat_B[9][27] +
                  mat_A[2][10] * mat_B[10][27] +
                  mat_A[2][11] * mat_B[11][27] +
                  mat_A[2][12] * mat_B[12][27] +
                  mat_A[2][13] * mat_B[13][27] +
                  mat_A[2][14] * mat_B[14][27] +
                  mat_A[2][15] * mat_B[15][27] +
                  mat_A[2][16] * mat_B[16][27] +
                  mat_A[2][17] * mat_B[17][27] +
                  mat_A[2][18] * mat_B[18][27] +
                  mat_A[2][19] * mat_B[19][27] +
                  mat_A[2][20] * mat_B[20][27] +
                  mat_A[2][21] * mat_B[21][27] +
                  mat_A[2][22] * mat_B[22][27] +
                  mat_A[2][23] * mat_B[23][27] +
                  mat_A[2][24] * mat_B[24][27] +
                  mat_A[2][25] * mat_B[25][27] +
                  mat_A[2][26] * mat_B[26][27] +
                  mat_A[2][27] * mat_B[27][27] +
                  mat_A[2][28] * mat_B[28][27] +
                  mat_A[2][29] * mat_B[29][27] +
                  mat_A[2][30] * mat_B[30][27] +
                  mat_A[2][31] * mat_B[31][27];
    mat_C[2][28] <= 
                  mat_A[2][0] * mat_B[0][28] +
                  mat_A[2][1] * mat_B[1][28] +
                  mat_A[2][2] * mat_B[2][28] +
                  mat_A[2][3] * mat_B[3][28] +
                  mat_A[2][4] * mat_B[4][28] +
                  mat_A[2][5] * mat_B[5][28] +
                  mat_A[2][6] * mat_B[6][28] +
                  mat_A[2][7] * mat_B[7][28] +
                  mat_A[2][8] * mat_B[8][28] +
                  mat_A[2][9] * mat_B[9][28] +
                  mat_A[2][10] * mat_B[10][28] +
                  mat_A[2][11] * mat_B[11][28] +
                  mat_A[2][12] * mat_B[12][28] +
                  mat_A[2][13] * mat_B[13][28] +
                  mat_A[2][14] * mat_B[14][28] +
                  mat_A[2][15] * mat_B[15][28] +
                  mat_A[2][16] * mat_B[16][28] +
                  mat_A[2][17] * mat_B[17][28] +
                  mat_A[2][18] * mat_B[18][28] +
                  mat_A[2][19] * mat_B[19][28] +
                  mat_A[2][20] * mat_B[20][28] +
                  mat_A[2][21] * mat_B[21][28] +
                  mat_A[2][22] * mat_B[22][28] +
                  mat_A[2][23] * mat_B[23][28] +
                  mat_A[2][24] * mat_B[24][28] +
                  mat_A[2][25] * mat_B[25][28] +
                  mat_A[2][26] * mat_B[26][28] +
                  mat_A[2][27] * mat_B[27][28] +
                  mat_A[2][28] * mat_B[28][28] +
                  mat_A[2][29] * mat_B[29][28] +
                  mat_A[2][30] * mat_B[30][28] +
                  mat_A[2][31] * mat_B[31][28];
    mat_C[2][29] <= 
                  mat_A[2][0] * mat_B[0][29] +
                  mat_A[2][1] * mat_B[1][29] +
                  mat_A[2][2] * mat_B[2][29] +
                  mat_A[2][3] * mat_B[3][29] +
                  mat_A[2][4] * mat_B[4][29] +
                  mat_A[2][5] * mat_B[5][29] +
                  mat_A[2][6] * mat_B[6][29] +
                  mat_A[2][7] * mat_B[7][29] +
                  mat_A[2][8] * mat_B[8][29] +
                  mat_A[2][9] * mat_B[9][29] +
                  mat_A[2][10] * mat_B[10][29] +
                  mat_A[2][11] * mat_B[11][29] +
                  mat_A[2][12] * mat_B[12][29] +
                  mat_A[2][13] * mat_B[13][29] +
                  mat_A[2][14] * mat_B[14][29] +
                  mat_A[2][15] * mat_B[15][29] +
                  mat_A[2][16] * mat_B[16][29] +
                  mat_A[2][17] * mat_B[17][29] +
                  mat_A[2][18] * mat_B[18][29] +
                  mat_A[2][19] * mat_B[19][29] +
                  mat_A[2][20] * mat_B[20][29] +
                  mat_A[2][21] * mat_B[21][29] +
                  mat_A[2][22] * mat_B[22][29] +
                  mat_A[2][23] * mat_B[23][29] +
                  mat_A[2][24] * mat_B[24][29] +
                  mat_A[2][25] * mat_B[25][29] +
                  mat_A[2][26] * mat_B[26][29] +
                  mat_A[2][27] * mat_B[27][29] +
                  mat_A[2][28] * mat_B[28][29] +
                  mat_A[2][29] * mat_B[29][29] +
                  mat_A[2][30] * mat_B[30][29] +
                  mat_A[2][31] * mat_B[31][29];
    mat_C[2][30] <= 
                  mat_A[2][0] * mat_B[0][30] +
                  mat_A[2][1] * mat_B[1][30] +
                  mat_A[2][2] * mat_B[2][30] +
                  mat_A[2][3] * mat_B[3][30] +
                  mat_A[2][4] * mat_B[4][30] +
                  mat_A[2][5] * mat_B[5][30] +
                  mat_A[2][6] * mat_B[6][30] +
                  mat_A[2][7] * mat_B[7][30] +
                  mat_A[2][8] * mat_B[8][30] +
                  mat_A[2][9] * mat_B[9][30] +
                  mat_A[2][10] * mat_B[10][30] +
                  mat_A[2][11] * mat_B[11][30] +
                  mat_A[2][12] * mat_B[12][30] +
                  mat_A[2][13] * mat_B[13][30] +
                  mat_A[2][14] * mat_B[14][30] +
                  mat_A[2][15] * mat_B[15][30] +
                  mat_A[2][16] * mat_B[16][30] +
                  mat_A[2][17] * mat_B[17][30] +
                  mat_A[2][18] * mat_B[18][30] +
                  mat_A[2][19] * mat_B[19][30] +
                  mat_A[2][20] * mat_B[20][30] +
                  mat_A[2][21] * mat_B[21][30] +
                  mat_A[2][22] * mat_B[22][30] +
                  mat_A[2][23] * mat_B[23][30] +
                  mat_A[2][24] * mat_B[24][30] +
                  mat_A[2][25] * mat_B[25][30] +
                  mat_A[2][26] * mat_B[26][30] +
                  mat_A[2][27] * mat_B[27][30] +
                  mat_A[2][28] * mat_B[28][30] +
                  mat_A[2][29] * mat_B[29][30] +
                  mat_A[2][30] * mat_B[30][30] +
                  mat_A[2][31] * mat_B[31][30];
    mat_C[2][31] <= 
                  mat_A[2][0] * mat_B[0][31] +
                  mat_A[2][1] * mat_B[1][31] +
                  mat_A[2][2] * mat_B[2][31] +
                  mat_A[2][3] * mat_B[3][31] +
                  mat_A[2][4] * mat_B[4][31] +
                  mat_A[2][5] * mat_B[5][31] +
                  mat_A[2][6] * mat_B[6][31] +
                  mat_A[2][7] * mat_B[7][31] +
                  mat_A[2][8] * mat_B[8][31] +
                  mat_A[2][9] * mat_B[9][31] +
                  mat_A[2][10] * mat_B[10][31] +
                  mat_A[2][11] * mat_B[11][31] +
                  mat_A[2][12] * mat_B[12][31] +
                  mat_A[2][13] * mat_B[13][31] +
                  mat_A[2][14] * mat_B[14][31] +
                  mat_A[2][15] * mat_B[15][31] +
                  mat_A[2][16] * mat_B[16][31] +
                  mat_A[2][17] * mat_B[17][31] +
                  mat_A[2][18] * mat_B[18][31] +
                  mat_A[2][19] * mat_B[19][31] +
                  mat_A[2][20] * mat_B[20][31] +
                  mat_A[2][21] * mat_B[21][31] +
                  mat_A[2][22] * mat_B[22][31] +
                  mat_A[2][23] * mat_B[23][31] +
                  mat_A[2][24] * mat_B[24][31] +
                  mat_A[2][25] * mat_B[25][31] +
                  mat_A[2][26] * mat_B[26][31] +
                  mat_A[2][27] * mat_B[27][31] +
                  mat_A[2][28] * mat_B[28][31] +
                  mat_A[2][29] * mat_B[29][31] +
                  mat_A[2][30] * mat_B[30][31] +
                  mat_A[2][31] * mat_B[31][31];
    mat_C[3][0] <= 
                  mat_A[3][0] * mat_B[0][0] +
                  mat_A[3][1] * mat_B[1][0] +
                  mat_A[3][2] * mat_B[2][0] +
                  mat_A[3][3] * mat_B[3][0] +
                  mat_A[3][4] * mat_B[4][0] +
                  mat_A[3][5] * mat_B[5][0] +
                  mat_A[3][6] * mat_B[6][0] +
                  mat_A[3][7] * mat_B[7][0] +
                  mat_A[3][8] * mat_B[8][0] +
                  mat_A[3][9] * mat_B[9][0] +
                  mat_A[3][10] * mat_B[10][0] +
                  mat_A[3][11] * mat_B[11][0] +
                  mat_A[3][12] * mat_B[12][0] +
                  mat_A[3][13] * mat_B[13][0] +
                  mat_A[3][14] * mat_B[14][0] +
                  mat_A[3][15] * mat_B[15][0] +
                  mat_A[3][16] * mat_B[16][0] +
                  mat_A[3][17] * mat_B[17][0] +
                  mat_A[3][18] * mat_B[18][0] +
                  mat_A[3][19] * mat_B[19][0] +
                  mat_A[3][20] * mat_B[20][0] +
                  mat_A[3][21] * mat_B[21][0] +
                  mat_A[3][22] * mat_B[22][0] +
                  mat_A[3][23] * mat_B[23][0] +
                  mat_A[3][24] * mat_B[24][0] +
                  mat_A[3][25] * mat_B[25][0] +
                  mat_A[3][26] * mat_B[26][0] +
                  mat_A[3][27] * mat_B[27][0] +
                  mat_A[3][28] * mat_B[28][0] +
                  mat_A[3][29] * mat_B[29][0] +
                  mat_A[3][30] * mat_B[30][0] +
                  mat_A[3][31] * mat_B[31][0];
    mat_C[3][1] <= 
                  mat_A[3][0] * mat_B[0][1] +
                  mat_A[3][1] * mat_B[1][1] +
                  mat_A[3][2] * mat_B[2][1] +
                  mat_A[3][3] * mat_B[3][1] +
                  mat_A[3][4] * mat_B[4][1] +
                  mat_A[3][5] * mat_B[5][1] +
                  mat_A[3][6] * mat_B[6][1] +
                  mat_A[3][7] * mat_B[7][1] +
                  mat_A[3][8] * mat_B[8][1] +
                  mat_A[3][9] * mat_B[9][1] +
                  mat_A[3][10] * mat_B[10][1] +
                  mat_A[3][11] * mat_B[11][1] +
                  mat_A[3][12] * mat_B[12][1] +
                  mat_A[3][13] * mat_B[13][1] +
                  mat_A[3][14] * mat_B[14][1] +
                  mat_A[3][15] * mat_B[15][1] +
                  mat_A[3][16] * mat_B[16][1] +
                  mat_A[3][17] * mat_B[17][1] +
                  mat_A[3][18] * mat_B[18][1] +
                  mat_A[3][19] * mat_B[19][1] +
                  mat_A[3][20] * mat_B[20][1] +
                  mat_A[3][21] * mat_B[21][1] +
                  mat_A[3][22] * mat_B[22][1] +
                  mat_A[3][23] * mat_B[23][1] +
                  mat_A[3][24] * mat_B[24][1] +
                  mat_A[3][25] * mat_B[25][1] +
                  mat_A[3][26] * mat_B[26][1] +
                  mat_A[3][27] * mat_B[27][1] +
                  mat_A[3][28] * mat_B[28][1] +
                  mat_A[3][29] * mat_B[29][1] +
                  mat_A[3][30] * mat_B[30][1] +
                  mat_A[3][31] * mat_B[31][1];
    mat_C[3][2] <= 
                  mat_A[3][0] * mat_B[0][2] +
                  mat_A[3][1] * mat_B[1][2] +
                  mat_A[3][2] * mat_B[2][2] +
                  mat_A[3][3] * mat_B[3][2] +
                  mat_A[3][4] * mat_B[4][2] +
                  mat_A[3][5] * mat_B[5][2] +
                  mat_A[3][6] * mat_B[6][2] +
                  mat_A[3][7] * mat_B[7][2] +
                  mat_A[3][8] * mat_B[8][2] +
                  mat_A[3][9] * mat_B[9][2] +
                  mat_A[3][10] * mat_B[10][2] +
                  mat_A[3][11] * mat_B[11][2] +
                  mat_A[3][12] * mat_B[12][2] +
                  mat_A[3][13] * mat_B[13][2] +
                  mat_A[3][14] * mat_B[14][2] +
                  mat_A[3][15] * mat_B[15][2] +
                  mat_A[3][16] * mat_B[16][2] +
                  mat_A[3][17] * mat_B[17][2] +
                  mat_A[3][18] * mat_B[18][2] +
                  mat_A[3][19] * mat_B[19][2] +
                  mat_A[3][20] * mat_B[20][2] +
                  mat_A[3][21] * mat_B[21][2] +
                  mat_A[3][22] * mat_B[22][2] +
                  mat_A[3][23] * mat_B[23][2] +
                  mat_A[3][24] * mat_B[24][2] +
                  mat_A[3][25] * mat_B[25][2] +
                  mat_A[3][26] * mat_B[26][2] +
                  mat_A[3][27] * mat_B[27][2] +
                  mat_A[3][28] * mat_B[28][2] +
                  mat_A[3][29] * mat_B[29][2] +
                  mat_A[3][30] * mat_B[30][2] +
                  mat_A[3][31] * mat_B[31][2];
    mat_C[3][3] <= 
                  mat_A[3][0] * mat_B[0][3] +
                  mat_A[3][1] * mat_B[1][3] +
                  mat_A[3][2] * mat_B[2][3] +
                  mat_A[3][3] * mat_B[3][3] +
                  mat_A[3][4] * mat_B[4][3] +
                  mat_A[3][5] * mat_B[5][3] +
                  mat_A[3][6] * mat_B[6][3] +
                  mat_A[3][7] * mat_B[7][3] +
                  mat_A[3][8] * mat_B[8][3] +
                  mat_A[3][9] * mat_B[9][3] +
                  mat_A[3][10] * mat_B[10][3] +
                  mat_A[3][11] * mat_B[11][3] +
                  mat_A[3][12] * mat_B[12][3] +
                  mat_A[3][13] * mat_B[13][3] +
                  mat_A[3][14] * mat_B[14][3] +
                  mat_A[3][15] * mat_B[15][3] +
                  mat_A[3][16] * mat_B[16][3] +
                  mat_A[3][17] * mat_B[17][3] +
                  mat_A[3][18] * mat_B[18][3] +
                  mat_A[3][19] * mat_B[19][3] +
                  mat_A[3][20] * mat_B[20][3] +
                  mat_A[3][21] * mat_B[21][3] +
                  mat_A[3][22] * mat_B[22][3] +
                  mat_A[3][23] * mat_B[23][3] +
                  mat_A[3][24] * mat_B[24][3] +
                  mat_A[3][25] * mat_B[25][3] +
                  mat_A[3][26] * mat_B[26][3] +
                  mat_A[3][27] * mat_B[27][3] +
                  mat_A[3][28] * mat_B[28][3] +
                  mat_A[3][29] * mat_B[29][3] +
                  mat_A[3][30] * mat_B[30][3] +
                  mat_A[3][31] * mat_B[31][3];
    mat_C[3][4] <= 
                  mat_A[3][0] * mat_B[0][4] +
                  mat_A[3][1] * mat_B[1][4] +
                  mat_A[3][2] * mat_B[2][4] +
                  mat_A[3][3] * mat_B[3][4] +
                  mat_A[3][4] * mat_B[4][4] +
                  mat_A[3][5] * mat_B[5][4] +
                  mat_A[3][6] * mat_B[6][4] +
                  mat_A[3][7] * mat_B[7][4] +
                  mat_A[3][8] * mat_B[8][4] +
                  mat_A[3][9] * mat_B[9][4] +
                  mat_A[3][10] * mat_B[10][4] +
                  mat_A[3][11] * mat_B[11][4] +
                  mat_A[3][12] * mat_B[12][4] +
                  mat_A[3][13] * mat_B[13][4] +
                  mat_A[3][14] * mat_B[14][4] +
                  mat_A[3][15] * mat_B[15][4] +
                  mat_A[3][16] * mat_B[16][4] +
                  mat_A[3][17] * mat_B[17][4] +
                  mat_A[3][18] * mat_B[18][4] +
                  mat_A[3][19] * mat_B[19][4] +
                  mat_A[3][20] * mat_B[20][4] +
                  mat_A[3][21] * mat_B[21][4] +
                  mat_A[3][22] * mat_B[22][4] +
                  mat_A[3][23] * mat_B[23][4] +
                  mat_A[3][24] * mat_B[24][4] +
                  mat_A[3][25] * mat_B[25][4] +
                  mat_A[3][26] * mat_B[26][4] +
                  mat_A[3][27] * mat_B[27][4] +
                  mat_A[3][28] * mat_B[28][4] +
                  mat_A[3][29] * mat_B[29][4] +
                  mat_A[3][30] * mat_B[30][4] +
                  mat_A[3][31] * mat_B[31][4];
    mat_C[3][5] <= 
                  mat_A[3][0] * mat_B[0][5] +
                  mat_A[3][1] * mat_B[1][5] +
                  mat_A[3][2] * mat_B[2][5] +
                  mat_A[3][3] * mat_B[3][5] +
                  mat_A[3][4] * mat_B[4][5] +
                  mat_A[3][5] * mat_B[5][5] +
                  mat_A[3][6] * mat_B[6][5] +
                  mat_A[3][7] * mat_B[7][5] +
                  mat_A[3][8] * mat_B[8][5] +
                  mat_A[3][9] * mat_B[9][5] +
                  mat_A[3][10] * mat_B[10][5] +
                  mat_A[3][11] * mat_B[11][5] +
                  mat_A[3][12] * mat_B[12][5] +
                  mat_A[3][13] * mat_B[13][5] +
                  mat_A[3][14] * mat_B[14][5] +
                  mat_A[3][15] * mat_B[15][5] +
                  mat_A[3][16] * mat_B[16][5] +
                  mat_A[3][17] * mat_B[17][5] +
                  mat_A[3][18] * mat_B[18][5] +
                  mat_A[3][19] * mat_B[19][5] +
                  mat_A[3][20] * mat_B[20][5] +
                  mat_A[3][21] * mat_B[21][5] +
                  mat_A[3][22] * mat_B[22][5] +
                  mat_A[3][23] * mat_B[23][5] +
                  mat_A[3][24] * mat_B[24][5] +
                  mat_A[3][25] * mat_B[25][5] +
                  mat_A[3][26] * mat_B[26][5] +
                  mat_A[3][27] * mat_B[27][5] +
                  mat_A[3][28] * mat_B[28][5] +
                  mat_A[3][29] * mat_B[29][5] +
                  mat_A[3][30] * mat_B[30][5] +
                  mat_A[3][31] * mat_B[31][5];
    mat_C[3][6] <= 
                  mat_A[3][0] * mat_B[0][6] +
                  mat_A[3][1] * mat_B[1][6] +
                  mat_A[3][2] * mat_B[2][6] +
                  mat_A[3][3] * mat_B[3][6] +
                  mat_A[3][4] * mat_B[4][6] +
                  mat_A[3][5] * mat_B[5][6] +
                  mat_A[3][6] * mat_B[6][6] +
                  mat_A[3][7] * mat_B[7][6] +
                  mat_A[3][8] * mat_B[8][6] +
                  mat_A[3][9] * mat_B[9][6] +
                  mat_A[3][10] * mat_B[10][6] +
                  mat_A[3][11] * mat_B[11][6] +
                  mat_A[3][12] * mat_B[12][6] +
                  mat_A[3][13] * mat_B[13][6] +
                  mat_A[3][14] * mat_B[14][6] +
                  mat_A[3][15] * mat_B[15][6] +
                  mat_A[3][16] * mat_B[16][6] +
                  mat_A[3][17] * mat_B[17][6] +
                  mat_A[3][18] * mat_B[18][6] +
                  mat_A[3][19] * mat_B[19][6] +
                  mat_A[3][20] * mat_B[20][6] +
                  mat_A[3][21] * mat_B[21][6] +
                  mat_A[3][22] * mat_B[22][6] +
                  mat_A[3][23] * mat_B[23][6] +
                  mat_A[3][24] * mat_B[24][6] +
                  mat_A[3][25] * mat_B[25][6] +
                  mat_A[3][26] * mat_B[26][6] +
                  mat_A[3][27] * mat_B[27][6] +
                  mat_A[3][28] * mat_B[28][6] +
                  mat_A[3][29] * mat_B[29][6] +
                  mat_A[3][30] * mat_B[30][6] +
                  mat_A[3][31] * mat_B[31][6];
    mat_C[3][7] <= 
                  mat_A[3][0] * mat_B[0][7] +
                  mat_A[3][1] * mat_B[1][7] +
                  mat_A[3][2] * mat_B[2][7] +
                  mat_A[3][3] * mat_B[3][7] +
                  mat_A[3][4] * mat_B[4][7] +
                  mat_A[3][5] * mat_B[5][7] +
                  mat_A[3][6] * mat_B[6][7] +
                  mat_A[3][7] * mat_B[7][7] +
                  mat_A[3][8] * mat_B[8][7] +
                  mat_A[3][9] * mat_B[9][7] +
                  mat_A[3][10] * mat_B[10][7] +
                  mat_A[3][11] * mat_B[11][7] +
                  mat_A[3][12] * mat_B[12][7] +
                  mat_A[3][13] * mat_B[13][7] +
                  mat_A[3][14] * mat_B[14][7] +
                  mat_A[3][15] * mat_B[15][7] +
                  mat_A[3][16] * mat_B[16][7] +
                  mat_A[3][17] * mat_B[17][7] +
                  mat_A[3][18] * mat_B[18][7] +
                  mat_A[3][19] * mat_B[19][7] +
                  mat_A[3][20] * mat_B[20][7] +
                  mat_A[3][21] * mat_B[21][7] +
                  mat_A[3][22] * mat_B[22][7] +
                  mat_A[3][23] * mat_B[23][7] +
                  mat_A[3][24] * mat_B[24][7] +
                  mat_A[3][25] * mat_B[25][7] +
                  mat_A[3][26] * mat_B[26][7] +
                  mat_A[3][27] * mat_B[27][7] +
                  mat_A[3][28] * mat_B[28][7] +
                  mat_A[3][29] * mat_B[29][7] +
                  mat_A[3][30] * mat_B[30][7] +
                  mat_A[3][31] * mat_B[31][7];
    mat_C[3][8] <= 
                  mat_A[3][0] * mat_B[0][8] +
                  mat_A[3][1] * mat_B[1][8] +
                  mat_A[3][2] * mat_B[2][8] +
                  mat_A[3][3] * mat_B[3][8] +
                  mat_A[3][4] * mat_B[4][8] +
                  mat_A[3][5] * mat_B[5][8] +
                  mat_A[3][6] * mat_B[6][8] +
                  mat_A[3][7] * mat_B[7][8] +
                  mat_A[3][8] * mat_B[8][8] +
                  mat_A[3][9] * mat_B[9][8] +
                  mat_A[3][10] * mat_B[10][8] +
                  mat_A[3][11] * mat_B[11][8] +
                  mat_A[3][12] * mat_B[12][8] +
                  mat_A[3][13] * mat_B[13][8] +
                  mat_A[3][14] * mat_B[14][8] +
                  mat_A[3][15] * mat_B[15][8] +
                  mat_A[3][16] * mat_B[16][8] +
                  mat_A[3][17] * mat_B[17][8] +
                  mat_A[3][18] * mat_B[18][8] +
                  mat_A[3][19] * mat_B[19][8] +
                  mat_A[3][20] * mat_B[20][8] +
                  mat_A[3][21] * mat_B[21][8] +
                  mat_A[3][22] * mat_B[22][8] +
                  mat_A[3][23] * mat_B[23][8] +
                  mat_A[3][24] * mat_B[24][8] +
                  mat_A[3][25] * mat_B[25][8] +
                  mat_A[3][26] * mat_B[26][8] +
                  mat_A[3][27] * mat_B[27][8] +
                  mat_A[3][28] * mat_B[28][8] +
                  mat_A[3][29] * mat_B[29][8] +
                  mat_A[3][30] * mat_B[30][8] +
                  mat_A[3][31] * mat_B[31][8];
    mat_C[3][9] <= 
                  mat_A[3][0] * mat_B[0][9] +
                  mat_A[3][1] * mat_B[1][9] +
                  mat_A[3][2] * mat_B[2][9] +
                  mat_A[3][3] * mat_B[3][9] +
                  mat_A[3][4] * mat_B[4][9] +
                  mat_A[3][5] * mat_B[5][9] +
                  mat_A[3][6] * mat_B[6][9] +
                  mat_A[3][7] * mat_B[7][9] +
                  mat_A[3][8] * mat_B[8][9] +
                  mat_A[3][9] * mat_B[9][9] +
                  mat_A[3][10] * mat_B[10][9] +
                  mat_A[3][11] * mat_B[11][9] +
                  mat_A[3][12] * mat_B[12][9] +
                  mat_A[3][13] * mat_B[13][9] +
                  mat_A[3][14] * mat_B[14][9] +
                  mat_A[3][15] * mat_B[15][9] +
                  mat_A[3][16] * mat_B[16][9] +
                  mat_A[3][17] * mat_B[17][9] +
                  mat_A[3][18] * mat_B[18][9] +
                  mat_A[3][19] * mat_B[19][9] +
                  mat_A[3][20] * mat_B[20][9] +
                  mat_A[3][21] * mat_B[21][9] +
                  mat_A[3][22] * mat_B[22][9] +
                  mat_A[3][23] * mat_B[23][9] +
                  mat_A[3][24] * mat_B[24][9] +
                  mat_A[3][25] * mat_B[25][9] +
                  mat_A[3][26] * mat_B[26][9] +
                  mat_A[3][27] * mat_B[27][9] +
                  mat_A[3][28] * mat_B[28][9] +
                  mat_A[3][29] * mat_B[29][9] +
                  mat_A[3][30] * mat_B[30][9] +
                  mat_A[3][31] * mat_B[31][9];
    mat_C[3][10] <= 
                  mat_A[3][0] * mat_B[0][10] +
                  mat_A[3][1] * mat_B[1][10] +
                  mat_A[3][2] * mat_B[2][10] +
                  mat_A[3][3] * mat_B[3][10] +
                  mat_A[3][4] * mat_B[4][10] +
                  mat_A[3][5] * mat_B[5][10] +
                  mat_A[3][6] * mat_B[6][10] +
                  mat_A[3][7] * mat_B[7][10] +
                  mat_A[3][8] * mat_B[8][10] +
                  mat_A[3][9] * mat_B[9][10] +
                  mat_A[3][10] * mat_B[10][10] +
                  mat_A[3][11] * mat_B[11][10] +
                  mat_A[3][12] * mat_B[12][10] +
                  mat_A[3][13] * mat_B[13][10] +
                  mat_A[3][14] * mat_B[14][10] +
                  mat_A[3][15] * mat_B[15][10] +
                  mat_A[3][16] * mat_B[16][10] +
                  mat_A[3][17] * mat_B[17][10] +
                  mat_A[3][18] * mat_B[18][10] +
                  mat_A[3][19] * mat_B[19][10] +
                  mat_A[3][20] * mat_B[20][10] +
                  mat_A[3][21] * mat_B[21][10] +
                  mat_A[3][22] * mat_B[22][10] +
                  mat_A[3][23] * mat_B[23][10] +
                  mat_A[3][24] * mat_B[24][10] +
                  mat_A[3][25] * mat_B[25][10] +
                  mat_A[3][26] * mat_B[26][10] +
                  mat_A[3][27] * mat_B[27][10] +
                  mat_A[3][28] * mat_B[28][10] +
                  mat_A[3][29] * mat_B[29][10] +
                  mat_A[3][30] * mat_B[30][10] +
                  mat_A[3][31] * mat_B[31][10];
    mat_C[3][11] <= 
                  mat_A[3][0] * mat_B[0][11] +
                  mat_A[3][1] * mat_B[1][11] +
                  mat_A[3][2] * mat_B[2][11] +
                  mat_A[3][3] * mat_B[3][11] +
                  mat_A[3][4] * mat_B[4][11] +
                  mat_A[3][5] * mat_B[5][11] +
                  mat_A[3][6] * mat_B[6][11] +
                  mat_A[3][7] * mat_B[7][11] +
                  mat_A[3][8] * mat_B[8][11] +
                  mat_A[3][9] * mat_B[9][11] +
                  mat_A[3][10] * mat_B[10][11] +
                  mat_A[3][11] * mat_B[11][11] +
                  mat_A[3][12] * mat_B[12][11] +
                  mat_A[3][13] * mat_B[13][11] +
                  mat_A[3][14] * mat_B[14][11] +
                  mat_A[3][15] * mat_B[15][11] +
                  mat_A[3][16] * mat_B[16][11] +
                  mat_A[3][17] * mat_B[17][11] +
                  mat_A[3][18] * mat_B[18][11] +
                  mat_A[3][19] * mat_B[19][11] +
                  mat_A[3][20] * mat_B[20][11] +
                  mat_A[3][21] * mat_B[21][11] +
                  mat_A[3][22] * mat_B[22][11] +
                  mat_A[3][23] * mat_B[23][11] +
                  mat_A[3][24] * mat_B[24][11] +
                  mat_A[3][25] * mat_B[25][11] +
                  mat_A[3][26] * mat_B[26][11] +
                  mat_A[3][27] * mat_B[27][11] +
                  mat_A[3][28] * mat_B[28][11] +
                  mat_A[3][29] * mat_B[29][11] +
                  mat_A[3][30] * mat_B[30][11] +
                  mat_A[3][31] * mat_B[31][11];
    mat_C[3][12] <= 
                  mat_A[3][0] * mat_B[0][12] +
                  mat_A[3][1] * mat_B[1][12] +
                  mat_A[3][2] * mat_B[2][12] +
                  mat_A[3][3] * mat_B[3][12] +
                  mat_A[3][4] * mat_B[4][12] +
                  mat_A[3][5] * mat_B[5][12] +
                  mat_A[3][6] * mat_B[6][12] +
                  mat_A[3][7] * mat_B[7][12] +
                  mat_A[3][8] * mat_B[8][12] +
                  mat_A[3][9] * mat_B[9][12] +
                  mat_A[3][10] * mat_B[10][12] +
                  mat_A[3][11] * mat_B[11][12] +
                  mat_A[3][12] * mat_B[12][12] +
                  mat_A[3][13] * mat_B[13][12] +
                  mat_A[3][14] * mat_B[14][12] +
                  mat_A[3][15] * mat_B[15][12] +
                  mat_A[3][16] * mat_B[16][12] +
                  mat_A[3][17] * mat_B[17][12] +
                  mat_A[3][18] * mat_B[18][12] +
                  mat_A[3][19] * mat_B[19][12] +
                  mat_A[3][20] * mat_B[20][12] +
                  mat_A[3][21] * mat_B[21][12] +
                  mat_A[3][22] * mat_B[22][12] +
                  mat_A[3][23] * mat_B[23][12] +
                  mat_A[3][24] * mat_B[24][12] +
                  mat_A[3][25] * mat_B[25][12] +
                  mat_A[3][26] * mat_B[26][12] +
                  mat_A[3][27] * mat_B[27][12] +
                  mat_A[3][28] * mat_B[28][12] +
                  mat_A[3][29] * mat_B[29][12] +
                  mat_A[3][30] * mat_B[30][12] +
                  mat_A[3][31] * mat_B[31][12];
    mat_C[3][13] <= 
                  mat_A[3][0] * mat_B[0][13] +
                  mat_A[3][1] * mat_B[1][13] +
                  mat_A[3][2] * mat_B[2][13] +
                  mat_A[3][3] * mat_B[3][13] +
                  mat_A[3][4] * mat_B[4][13] +
                  mat_A[3][5] * mat_B[5][13] +
                  mat_A[3][6] * mat_B[6][13] +
                  mat_A[3][7] * mat_B[7][13] +
                  mat_A[3][8] * mat_B[8][13] +
                  mat_A[3][9] * mat_B[9][13] +
                  mat_A[3][10] * mat_B[10][13] +
                  mat_A[3][11] * mat_B[11][13] +
                  mat_A[3][12] * mat_B[12][13] +
                  mat_A[3][13] * mat_B[13][13] +
                  mat_A[3][14] * mat_B[14][13] +
                  mat_A[3][15] * mat_B[15][13] +
                  mat_A[3][16] * mat_B[16][13] +
                  mat_A[3][17] * mat_B[17][13] +
                  mat_A[3][18] * mat_B[18][13] +
                  mat_A[3][19] * mat_B[19][13] +
                  mat_A[3][20] * mat_B[20][13] +
                  mat_A[3][21] * mat_B[21][13] +
                  mat_A[3][22] * mat_B[22][13] +
                  mat_A[3][23] * mat_B[23][13] +
                  mat_A[3][24] * mat_B[24][13] +
                  mat_A[3][25] * mat_B[25][13] +
                  mat_A[3][26] * mat_B[26][13] +
                  mat_A[3][27] * mat_B[27][13] +
                  mat_A[3][28] * mat_B[28][13] +
                  mat_A[3][29] * mat_B[29][13] +
                  mat_A[3][30] * mat_B[30][13] +
                  mat_A[3][31] * mat_B[31][13];
    mat_C[3][14] <= 
                  mat_A[3][0] * mat_B[0][14] +
                  mat_A[3][1] * mat_B[1][14] +
                  mat_A[3][2] * mat_B[2][14] +
                  mat_A[3][3] * mat_B[3][14] +
                  mat_A[3][4] * mat_B[4][14] +
                  mat_A[3][5] * mat_B[5][14] +
                  mat_A[3][6] * mat_B[6][14] +
                  mat_A[3][7] * mat_B[7][14] +
                  mat_A[3][8] * mat_B[8][14] +
                  mat_A[3][9] * mat_B[9][14] +
                  mat_A[3][10] * mat_B[10][14] +
                  mat_A[3][11] * mat_B[11][14] +
                  mat_A[3][12] * mat_B[12][14] +
                  mat_A[3][13] * mat_B[13][14] +
                  mat_A[3][14] * mat_B[14][14] +
                  mat_A[3][15] * mat_B[15][14] +
                  mat_A[3][16] * mat_B[16][14] +
                  mat_A[3][17] * mat_B[17][14] +
                  mat_A[3][18] * mat_B[18][14] +
                  mat_A[3][19] * mat_B[19][14] +
                  mat_A[3][20] * mat_B[20][14] +
                  mat_A[3][21] * mat_B[21][14] +
                  mat_A[3][22] * mat_B[22][14] +
                  mat_A[3][23] * mat_B[23][14] +
                  mat_A[3][24] * mat_B[24][14] +
                  mat_A[3][25] * mat_B[25][14] +
                  mat_A[3][26] * mat_B[26][14] +
                  mat_A[3][27] * mat_B[27][14] +
                  mat_A[3][28] * mat_B[28][14] +
                  mat_A[3][29] * mat_B[29][14] +
                  mat_A[3][30] * mat_B[30][14] +
                  mat_A[3][31] * mat_B[31][14];
    mat_C[3][15] <= 
                  mat_A[3][0] * mat_B[0][15] +
                  mat_A[3][1] * mat_B[1][15] +
                  mat_A[3][2] * mat_B[2][15] +
                  mat_A[3][3] * mat_B[3][15] +
                  mat_A[3][4] * mat_B[4][15] +
                  mat_A[3][5] * mat_B[5][15] +
                  mat_A[3][6] * mat_B[6][15] +
                  mat_A[3][7] * mat_B[7][15] +
                  mat_A[3][8] * mat_B[8][15] +
                  mat_A[3][9] * mat_B[9][15] +
                  mat_A[3][10] * mat_B[10][15] +
                  mat_A[3][11] * mat_B[11][15] +
                  mat_A[3][12] * mat_B[12][15] +
                  mat_A[3][13] * mat_B[13][15] +
                  mat_A[3][14] * mat_B[14][15] +
                  mat_A[3][15] * mat_B[15][15] +
                  mat_A[3][16] * mat_B[16][15] +
                  mat_A[3][17] * mat_B[17][15] +
                  mat_A[3][18] * mat_B[18][15] +
                  mat_A[3][19] * mat_B[19][15] +
                  mat_A[3][20] * mat_B[20][15] +
                  mat_A[3][21] * mat_B[21][15] +
                  mat_A[3][22] * mat_B[22][15] +
                  mat_A[3][23] * mat_B[23][15] +
                  mat_A[3][24] * mat_B[24][15] +
                  mat_A[3][25] * mat_B[25][15] +
                  mat_A[3][26] * mat_B[26][15] +
                  mat_A[3][27] * mat_B[27][15] +
                  mat_A[3][28] * mat_B[28][15] +
                  mat_A[3][29] * mat_B[29][15] +
                  mat_A[3][30] * mat_B[30][15] +
                  mat_A[3][31] * mat_B[31][15];
    mat_C[3][16] <= 
                  mat_A[3][0] * mat_B[0][16] +
                  mat_A[3][1] * mat_B[1][16] +
                  mat_A[3][2] * mat_B[2][16] +
                  mat_A[3][3] * mat_B[3][16] +
                  mat_A[3][4] * mat_B[4][16] +
                  mat_A[3][5] * mat_B[5][16] +
                  mat_A[3][6] * mat_B[6][16] +
                  mat_A[3][7] * mat_B[7][16] +
                  mat_A[3][8] * mat_B[8][16] +
                  mat_A[3][9] * mat_B[9][16] +
                  mat_A[3][10] * mat_B[10][16] +
                  mat_A[3][11] * mat_B[11][16] +
                  mat_A[3][12] * mat_B[12][16] +
                  mat_A[3][13] * mat_B[13][16] +
                  mat_A[3][14] * mat_B[14][16] +
                  mat_A[3][15] * mat_B[15][16] +
                  mat_A[3][16] * mat_B[16][16] +
                  mat_A[3][17] * mat_B[17][16] +
                  mat_A[3][18] * mat_B[18][16] +
                  mat_A[3][19] * mat_B[19][16] +
                  mat_A[3][20] * mat_B[20][16] +
                  mat_A[3][21] * mat_B[21][16] +
                  mat_A[3][22] * mat_B[22][16] +
                  mat_A[3][23] * mat_B[23][16] +
                  mat_A[3][24] * mat_B[24][16] +
                  mat_A[3][25] * mat_B[25][16] +
                  mat_A[3][26] * mat_B[26][16] +
                  mat_A[3][27] * mat_B[27][16] +
                  mat_A[3][28] * mat_B[28][16] +
                  mat_A[3][29] * mat_B[29][16] +
                  mat_A[3][30] * mat_B[30][16] +
                  mat_A[3][31] * mat_B[31][16];
    mat_C[3][17] <= 
                  mat_A[3][0] * mat_B[0][17] +
                  mat_A[3][1] * mat_B[1][17] +
                  mat_A[3][2] * mat_B[2][17] +
                  mat_A[3][3] * mat_B[3][17] +
                  mat_A[3][4] * mat_B[4][17] +
                  mat_A[3][5] * mat_B[5][17] +
                  mat_A[3][6] * mat_B[6][17] +
                  mat_A[3][7] * mat_B[7][17] +
                  mat_A[3][8] * mat_B[8][17] +
                  mat_A[3][9] * mat_B[9][17] +
                  mat_A[3][10] * mat_B[10][17] +
                  mat_A[3][11] * mat_B[11][17] +
                  mat_A[3][12] * mat_B[12][17] +
                  mat_A[3][13] * mat_B[13][17] +
                  mat_A[3][14] * mat_B[14][17] +
                  mat_A[3][15] * mat_B[15][17] +
                  mat_A[3][16] * mat_B[16][17] +
                  mat_A[3][17] * mat_B[17][17] +
                  mat_A[3][18] * mat_B[18][17] +
                  mat_A[3][19] * mat_B[19][17] +
                  mat_A[3][20] * mat_B[20][17] +
                  mat_A[3][21] * mat_B[21][17] +
                  mat_A[3][22] * mat_B[22][17] +
                  mat_A[3][23] * mat_B[23][17] +
                  mat_A[3][24] * mat_B[24][17] +
                  mat_A[3][25] * mat_B[25][17] +
                  mat_A[3][26] * mat_B[26][17] +
                  mat_A[3][27] * mat_B[27][17] +
                  mat_A[3][28] * mat_B[28][17] +
                  mat_A[3][29] * mat_B[29][17] +
                  mat_A[3][30] * mat_B[30][17] +
                  mat_A[3][31] * mat_B[31][17];
    mat_C[3][18] <= 
                  mat_A[3][0] * mat_B[0][18] +
                  mat_A[3][1] * mat_B[1][18] +
                  mat_A[3][2] * mat_B[2][18] +
                  mat_A[3][3] * mat_B[3][18] +
                  mat_A[3][4] * mat_B[4][18] +
                  mat_A[3][5] * mat_B[5][18] +
                  mat_A[3][6] * mat_B[6][18] +
                  mat_A[3][7] * mat_B[7][18] +
                  mat_A[3][8] * mat_B[8][18] +
                  mat_A[3][9] * mat_B[9][18] +
                  mat_A[3][10] * mat_B[10][18] +
                  mat_A[3][11] * mat_B[11][18] +
                  mat_A[3][12] * mat_B[12][18] +
                  mat_A[3][13] * mat_B[13][18] +
                  mat_A[3][14] * mat_B[14][18] +
                  mat_A[3][15] * mat_B[15][18] +
                  mat_A[3][16] * mat_B[16][18] +
                  mat_A[3][17] * mat_B[17][18] +
                  mat_A[3][18] * mat_B[18][18] +
                  mat_A[3][19] * mat_B[19][18] +
                  mat_A[3][20] * mat_B[20][18] +
                  mat_A[3][21] * mat_B[21][18] +
                  mat_A[3][22] * mat_B[22][18] +
                  mat_A[3][23] * mat_B[23][18] +
                  mat_A[3][24] * mat_B[24][18] +
                  mat_A[3][25] * mat_B[25][18] +
                  mat_A[3][26] * mat_B[26][18] +
                  mat_A[3][27] * mat_B[27][18] +
                  mat_A[3][28] * mat_B[28][18] +
                  mat_A[3][29] * mat_B[29][18] +
                  mat_A[3][30] * mat_B[30][18] +
                  mat_A[3][31] * mat_B[31][18];
    mat_C[3][19] <= 
                  mat_A[3][0] * mat_B[0][19] +
                  mat_A[3][1] * mat_B[1][19] +
                  mat_A[3][2] * mat_B[2][19] +
                  mat_A[3][3] * mat_B[3][19] +
                  mat_A[3][4] * mat_B[4][19] +
                  mat_A[3][5] * mat_B[5][19] +
                  mat_A[3][6] * mat_B[6][19] +
                  mat_A[3][7] * mat_B[7][19] +
                  mat_A[3][8] * mat_B[8][19] +
                  mat_A[3][9] * mat_B[9][19] +
                  mat_A[3][10] * mat_B[10][19] +
                  mat_A[3][11] * mat_B[11][19] +
                  mat_A[3][12] * mat_B[12][19] +
                  mat_A[3][13] * mat_B[13][19] +
                  mat_A[3][14] * mat_B[14][19] +
                  mat_A[3][15] * mat_B[15][19] +
                  mat_A[3][16] * mat_B[16][19] +
                  mat_A[3][17] * mat_B[17][19] +
                  mat_A[3][18] * mat_B[18][19] +
                  mat_A[3][19] * mat_B[19][19] +
                  mat_A[3][20] * mat_B[20][19] +
                  mat_A[3][21] * mat_B[21][19] +
                  mat_A[3][22] * mat_B[22][19] +
                  mat_A[3][23] * mat_B[23][19] +
                  mat_A[3][24] * mat_B[24][19] +
                  mat_A[3][25] * mat_B[25][19] +
                  mat_A[3][26] * mat_B[26][19] +
                  mat_A[3][27] * mat_B[27][19] +
                  mat_A[3][28] * mat_B[28][19] +
                  mat_A[3][29] * mat_B[29][19] +
                  mat_A[3][30] * mat_B[30][19] +
                  mat_A[3][31] * mat_B[31][19];
    mat_C[3][20] <= 
                  mat_A[3][0] * mat_B[0][20] +
                  mat_A[3][1] * mat_B[1][20] +
                  mat_A[3][2] * mat_B[2][20] +
                  mat_A[3][3] * mat_B[3][20] +
                  mat_A[3][4] * mat_B[4][20] +
                  mat_A[3][5] * mat_B[5][20] +
                  mat_A[3][6] * mat_B[6][20] +
                  mat_A[3][7] * mat_B[7][20] +
                  mat_A[3][8] * mat_B[8][20] +
                  mat_A[3][9] * mat_B[9][20] +
                  mat_A[3][10] * mat_B[10][20] +
                  mat_A[3][11] * mat_B[11][20] +
                  mat_A[3][12] * mat_B[12][20] +
                  mat_A[3][13] * mat_B[13][20] +
                  mat_A[3][14] * mat_B[14][20] +
                  mat_A[3][15] * mat_B[15][20] +
                  mat_A[3][16] * mat_B[16][20] +
                  mat_A[3][17] * mat_B[17][20] +
                  mat_A[3][18] * mat_B[18][20] +
                  mat_A[3][19] * mat_B[19][20] +
                  mat_A[3][20] * mat_B[20][20] +
                  mat_A[3][21] * mat_B[21][20] +
                  mat_A[3][22] * mat_B[22][20] +
                  mat_A[3][23] * mat_B[23][20] +
                  mat_A[3][24] * mat_B[24][20] +
                  mat_A[3][25] * mat_B[25][20] +
                  mat_A[3][26] * mat_B[26][20] +
                  mat_A[3][27] * mat_B[27][20] +
                  mat_A[3][28] * mat_B[28][20] +
                  mat_A[3][29] * mat_B[29][20] +
                  mat_A[3][30] * mat_B[30][20] +
                  mat_A[3][31] * mat_B[31][20];
    mat_C[3][21] <= 
                  mat_A[3][0] * mat_B[0][21] +
                  mat_A[3][1] * mat_B[1][21] +
                  mat_A[3][2] * mat_B[2][21] +
                  mat_A[3][3] * mat_B[3][21] +
                  mat_A[3][4] * mat_B[4][21] +
                  mat_A[3][5] * mat_B[5][21] +
                  mat_A[3][6] * mat_B[6][21] +
                  mat_A[3][7] * mat_B[7][21] +
                  mat_A[3][8] * mat_B[8][21] +
                  mat_A[3][9] * mat_B[9][21] +
                  mat_A[3][10] * mat_B[10][21] +
                  mat_A[3][11] * mat_B[11][21] +
                  mat_A[3][12] * mat_B[12][21] +
                  mat_A[3][13] * mat_B[13][21] +
                  mat_A[3][14] * mat_B[14][21] +
                  mat_A[3][15] * mat_B[15][21] +
                  mat_A[3][16] * mat_B[16][21] +
                  mat_A[3][17] * mat_B[17][21] +
                  mat_A[3][18] * mat_B[18][21] +
                  mat_A[3][19] * mat_B[19][21] +
                  mat_A[3][20] * mat_B[20][21] +
                  mat_A[3][21] * mat_B[21][21] +
                  mat_A[3][22] * mat_B[22][21] +
                  mat_A[3][23] * mat_B[23][21] +
                  mat_A[3][24] * mat_B[24][21] +
                  mat_A[3][25] * mat_B[25][21] +
                  mat_A[3][26] * mat_B[26][21] +
                  mat_A[3][27] * mat_B[27][21] +
                  mat_A[3][28] * mat_B[28][21] +
                  mat_A[3][29] * mat_B[29][21] +
                  mat_A[3][30] * mat_B[30][21] +
                  mat_A[3][31] * mat_B[31][21];
    mat_C[3][22] <= 
                  mat_A[3][0] * mat_B[0][22] +
                  mat_A[3][1] * mat_B[1][22] +
                  mat_A[3][2] * mat_B[2][22] +
                  mat_A[3][3] * mat_B[3][22] +
                  mat_A[3][4] * mat_B[4][22] +
                  mat_A[3][5] * mat_B[5][22] +
                  mat_A[3][6] * mat_B[6][22] +
                  mat_A[3][7] * mat_B[7][22] +
                  mat_A[3][8] * mat_B[8][22] +
                  mat_A[3][9] * mat_B[9][22] +
                  mat_A[3][10] * mat_B[10][22] +
                  mat_A[3][11] * mat_B[11][22] +
                  mat_A[3][12] * mat_B[12][22] +
                  mat_A[3][13] * mat_B[13][22] +
                  mat_A[3][14] * mat_B[14][22] +
                  mat_A[3][15] * mat_B[15][22] +
                  mat_A[3][16] * mat_B[16][22] +
                  mat_A[3][17] * mat_B[17][22] +
                  mat_A[3][18] * mat_B[18][22] +
                  mat_A[3][19] * mat_B[19][22] +
                  mat_A[3][20] * mat_B[20][22] +
                  mat_A[3][21] * mat_B[21][22] +
                  mat_A[3][22] * mat_B[22][22] +
                  mat_A[3][23] * mat_B[23][22] +
                  mat_A[3][24] * mat_B[24][22] +
                  mat_A[3][25] * mat_B[25][22] +
                  mat_A[3][26] * mat_B[26][22] +
                  mat_A[3][27] * mat_B[27][22] +
                  mat_A[3][28] * mat_B[28][22] +
                  mat_A[3][29] * mat_B[29][22] +
                  mat_A[3][30] * mat_B[30][22] +
                  mat_A[3][31] * mat_B[31][22];
    mat_C[3][23] <= 
                  mat_A[3][0] * mat_B[0][23] +
                  mat_A[3][1] * mat_B[1][23] +
                  mat_A[3][2] * mat_B[2][23] +
                  mat_A[3][3] * mat_B[3][23] +
                  mat_A[3][4] * mat_B[4][23] +
                  mat_A[3][5] * mat_B[5][23] +
                  mat_A[3][6] * mat_B[6][23] +
                  mat_A[3][7] * mat_B[7][23] +
                  mat_A[3][8] * mat_B[8][23] +
                  mat_A[3][9] * mat_B[9][23] +
                  mat_A[3][10] * mat_B[10][23] +
                  mat_A[3][11] * mat_B[11][23] +
                  mat_A[3][12] * mat_B[12][23] +
                  mat_A[3][13] * mat_B[13][23] +
                  mat_A[3][14] * mat_B[14][23] +
                  mat_A[3][15] * mat_B[15][23] +
                  mat_A[3][16] * mat_B[16][23] +
                  mat_A[3][17] * mat_B[17][23] +
                  mat_A[3][18] * mat_B[18][23] +
                  mat_A[3][19] * mat_B[19][23] +
                  mat_A[3][20] * mat_B[20][23] +
                  mat_A[3][21] * mat_B[21][23] +
                  mat_A[3][22] * mat_B[22][23] +
                  mat_A[3][23] * mat_B[23][23] +
                  mat_A[3][24] * mat_B[24][23] +
                  mat_A[3][25] * mat_B[25][23] +
                  mat_A[3][26] * mat_B[26][23] +
                  mat_A[3][27] * mat_B[27][23] +
                  mat_A[3][28] * mat_B[28][23] +
                  mat_A[3][29] * mat_B[29][23] +
                  mat_A[3][30] * mat_B[30][23] +
                  mat_A[3][31] * mat_B[31][23];
    mat_C[3][24] <= 
                  mat_A[3][0] * mat_B[0][24] +
                  mat_A[3][1] * mat_B[1][24] +
                  mat_A[3][2] * mat_B[2][24] +
                  mat_A[3][3] * mat_B[3][24] +
                  mat_A[3][4] * mat_B[4][24] +
                  mat_A[3][5] * mat_B[5][24] +
                  mat_A[3][6] * mat_B[6][24] +
                  mat_A[3][7] * mat_B[7][24] +
                  mat_A[3][8] * mat_B[8][24] +
                  mat_A[3][9] * mat_B[9][24] +
                  mat_A[3][10] * mat_B[10][24] +
                  mat_A[3][11] * mat_B[11][24] +
                  mat_A[3][12] * mat_B[12][24] +
                  mat_A[3][13] * mat_B[13][24] +
                  mat_A[3][14] * mat_B[14][24] +
                  mat_A[3][15] * mat_B[15][24] +
                  mat_A[3][16] * mat_B[16][24] +
                  mat_A[3][17] * mat_B[17][24] +
                  mat_A[3][18] * mat_B[18][24] +
                  mat_A[3][19] * mat_B[19][24] +
                  mat_A[3][20] * mat_B[20][24] +
                  mat_A[3][21] * mat_B[21][24] +
                  mat_A[3][22] * mat_B[22][24] +
                  mat_A[3][23] * mat_B[23][24] +
                  mat_A[3][24] * mat_B[24][24] +
                  mat_A[3][25] * mat_B[25][24] +
                  mat_A[3][26] * mat_B[26][24] +
                  mat_A[3][27] * mat_B[27][24] +
                  mat_A[3][28] * mat_B[28][24] +
                  mat_A[3][29] * mat_B[29][24] +
                  mat_A[3][30] * mat_B[30][24] +
                  mat_A[3][31] * mat_B[31][24];
    mat_C[3][25] <= 
                  mat_A[3][0] * mat_B[0][25] +
                  mat_A[3][1] * mat_B[1][25] +
                  mat_A[3][2] * mat_B[2][25] +
                  mat_A[3][3] * mat_B[3][25] +
                  mat_A[3][4] * mat_B[4][25] +
                  mat_A[3][5] * mat_B[5][25] +
                  mat_A[3][6] * mat_B[6][25] +
                  mat_A[3][7] * mat_B[7][25] +
                  mat_A[3][8] * mat_B[8][25] +
                  mat_A[3][9] * mat_B[9][25] +
                  mat_A[3][10] * mat_B[10][25] +
                  mat_A[3][11] * mat_B[11][25] +
                  mat_A[3][12] * mat_B[12][25] +
                  mat_A[3][13] * mat_B[13][25] +
                  mat_A[3][14] * mat_B[14][25] +
                  mat_A[3][15] * mat_B[15][25] +
                  mat_A[3][16] * mat_B[16][25] +
                  mat_A[3][17] * mat_B[17][25] +
                  mat_A[3][18] * mat_B[18][25] +
                  mat_A[3][19] * mat_B[19][25] +
                  mat_A[3][20] * mat_B[20][25] +
                  mat_A[3][21] * mat_B[21][25] +
                  mat_A[3][22] * mat_B[22][25] +
                  mat_A[3][23] * mat_B[23][25] +
                  mat_A[3][24] * mat_B[24][25] +
                  mat_A[3][25] * mat_B[25][25] +
                  mat_A[3][26] * mat_B[26][25] +
                  mat_A[3][27] * mat_B[27][25] +
                  mat_A[3][28] * mat_B[28][25] +
                  mat_A[3][29] * mat_B[29][25] +
                  mat_A[3][30] * mat_B[30][25] +
                  mat_A[3][31] * mat_B[31][25];
    mat_C[3][26] <= 
                  mat_A[3][0] * mat_B[0][26] +
                  mat_A[3][1] * mat_B[1][26] +
                  mat_A[3][2] * mat_B[2][26] +
                  mat_A[3][3] * mat_B[3][26] +
                  mat_A[3][4] * mat_B[4][26] +
                  mat_A[3][5] * mat_B[5][26] +
                  mat_A[3][6] * mat_B[6][26] +
                  mat_A[3][7] * mat_B[7][26] +
                  mat_A[3][8] * mat_B[8][26] +
                  mat_A[3][9] * mat_B[9][26] +
                  mat_A[3][10] * mat_B[10][26] +
                  mat_A[3][11] * mat_B[11][26] +
                  mat_A[3][12] * mat_B[12][26] +
                  mat_A[3][13] * mat_B[13][26] +
                  mat_A[3][14] * mat_B[14][26] +
                  mat_A[3][15] * mat_B[15][26] +
                  mat_A[3][16] * mat_B[16][26] +
                  mat_A[3][17] * mat_B[17][26] +
                  mat_A[3][18] * mat_B[18][26] +
                  mat_A[3][19] * mat_B[19][26] +
                  mat_A[3][20] * mat_B[20][26] +
                  mat_A[3][21] * mat_B[21][26] +
                  mat_A[3][22] * mat_B[22][26] +
                  mat_A[3][23] * mat_B[23][26] +
                  mat_A[3][24] * mat_B[24][26] +
                  mat_A[3][25] * mat_B[25][26] +
                  mat_A[3][26] * mat_B[26][26] +
                  mat_A[3][27] * mat_B[27][26] +
                  mat_A[3][28] * mat_B[28][26] +
                  mat_A[3][29] * mat_B[29][26] +
                  mat_A[3][30] * mat_B[30][26] +
                  mat_A[3][31] * mat_B[31][26];
    mat_C[3][27] <= 
                  mat_A[3][0] * mat_B[0][27] +
                  mat_A[3][1] * mat_B[1][27] +
                  mat_A[3][2] * mat_B[2][27] +
                  mat_A[3][3] * mat_B[3][27] +
                  mat_A[3][4] * mat_B[4][27] +
                  mat_A[3][5] * mat_B[5][27] +
                  mat_A[3][6] * mat_B[6][27] +
                  mat_A[3][7] * mat_B[7][27] +
                  mat_A[3][8] * mat_B[8][27] +
                  mat_A[3][9] * mat_B[9][27] +
                  mat_A[3][10] * mat_B[10][27] +
                  mat_A[3][11] * mat_B[11][27] +
                  mat_A[3][12] * mat_B[12][27] +
                  mat_A[3][13] * mat_B[13][27] +
                  mat_A[3][14] * mat_B[14][27] +
                  mat_A[3][15] * mat_B[15][27] +
                  mat_A[3][16] * mat_B[16][27] +
                  mat_A[3][17] * mat_B[17][27] +
                  mat_A[3][18] * mat_B[18][27] +
                  mat_A[3][19] * mat_B[19][27] +
                  mat_A[3][20] * mat_B[20][27] +
                  mat_A[3][21] * mat_B[21][27] +
                  mat_A[3][22] * mat_B[22][27] +
                  mat_A[3][23] * mat_B[23][27] +
                  mat_A[3][24] * mat_B[24][27] +
                  mat_A[3][25] * mat_B[25][27] +
                  mat_A[3][26] * mat_B[26][27] +
                  mat_A[3][27] * mat_B[27][27] +
                  mat_A[3][28] * mat_B[28][27] +
                  mat_A[3][29] * mat_B[29][27] +
                  mat_A[3][30] * mat_B[30][27] +
                  mat_A[3][31] * mat_B[31][27];
    mat_C[3][28] <= 
                  mat_A[3][0] * mat_B[0][28] +
                  mat_A[3][1] * mat_B[1][28] +
                  mat_A[3][2] * mat_B[2][28] +
                  mat_A[3][3] * mat_B[3][28] +
                  mat_A[3][4] * mat_B[4][28] +
                  mat_A[3][5] * mat_B[5][28] +
                  mat_A[3][6] * mat_B[6][28] +
                  mat_A[3][7] * mat_B[7][28] +
                  mat_A[3][8] * mat_B[8][28] +
                  mat_A[3][9] * mat_B[9][28] +
                  mat_A[3][10] * mat_B[10][28] +
                  mat_A[3][11] * mat_B[11][28] +
                  mat_A[3][12] * mat_B[12][28] +
                  mat_A[3][13] * mat_B[13][28] +
                  mat_A[3][14] * mat_B[14][28] +
                  mat_A[3][15] * mat_B[15][28] +
                  mat_A[3][16] * mat_B[16][28] +
                  mat_A[3][17] * mat_B[17][28] +
                  mat_A[3][18] * mat_B[18][28] +
                  mat_A[3][19] * mat_B[19][28] +
                  mat_A[3][20] * mat_B[20][28] +
                  mat_A[3][21] * mat_B[21][28] +
                  mat_A[3][22] * mat_B[22][28] +
                  mat_A[3][23] * mat_B[23][28] +
                  mat_A[3][24] * mat_B[24][28] +
                  mat_A[3][25] * mat_B[25][28] +
                  mat_A[3][26] * mat_B[26][28] +
                  mat_A[3][27] * mat_B[27][28] +
                  mat_A[3][28] * mat_B[28][28] +
                  mat_A[3][29] * mat_B[29][28] +
                  mat_A[3][30] * mat_B[30][28] +
                  mat_A[3][31] * mat_B[31][28];
    mat_C[3][29] <= 
                  mat_A[3][0] * mat_B[0][29] +
                  mat_A[3][1] * mat_B[1][29] +
                  mat_A[3][2] * mat_B[2][29] +
                  mat_A[3][3] * mat_B[3][29] +
                  mat_A[3][4] * mat_B[4][29] +
                  mat_A[3][5] * mat_B[5][29] +
                  mat_A[3][6] * mat_B[6][29] +
                  mat_A[3][7] * mat_B[7][29] +
                  mat_A[3][8] * mat_B[8][29] +
                  mat_A[3][9] * mat_B[9][29] +
                  mat_A[3][10] * mat_B[10][29] +
                  mat_A[3][11] * mat_B[11][29] +
                  mat_A[3][12] * mat_B[12][29] +
                  mat_A[3][13] * mat_B[13][29] +
                  mat_A[3][14] * mat_B[14][29] +
                  mat_A[3][15] * mat_B[15][29] +
                  mat_A[3][16] * mat_B[16][29] +
                  mat_A[3][17] * mat_B[17][29] +
                  mat_A[3][18] * mat_B[18][29] +
                  mat_A[3][19] * mat_B[19][29] +
                  mat_A[3][20] * mat_B[20][29] +
                  mat_A[3][21] * mat_B[21][29] +
                  mat_A[3][22] * mat_B[22][29] +
                  mat_A[3][23] * mat_B[23][29] +
                  mat_A[3][24] * mat_B[24][29] +
                  mat_A[3][25] * mat_B[25][29] +
                  mat_A[3][26] * mat_B[26][29] +
                  mat_A[3][27] * mat_B[27][29] +
                  mat_A[3][28] * mat_B[28][29] +
                  mat_A[3][29] * mat_B[29][29] +
                  mat_A[3][30] * mat_B[30][29] +
                  mat_A[3][31] * mat_B[31][29];
    mat_C[3][30] <= 
                  mat_A[3][0] * mat_B[0][30] +
                  mat_A[3][1] * mat_B[1][30] +
                  mat_A[3][2] * mat_B[2][30] +
                  mat_A[3][3] * mat_B[3][30] +
                  mat_A[3][4] * mat_B[4][30] +
                  mat_A[3][5] * mat_B[5][30] +
                  mat_A[3][6] * mat_B[6][30] +
                  mat_A[3][7] * mat_B[7][30] +
                  mat_A[3][8] * mat_B[8][30] +
                  mat_A[3][9] * mat_B[9][30] +
                  mat_A[3][10] * mat_B[10][30] +
                  mat_A[3][11] * mat_B[11][30] +
                  mat_A[3][12] * mat_B[12][30] +
                  mat_A[3][13] * mat_B[13][30] +
                  mat_A[3][14] * mat_B[14][30] +
                  mat_A[3][15] * mat_B[15][30] +
                  mat_A[3][16] * mat_B[16][30] +
                  mat_A[3][17] * mat_B[17][30] +
                  mat_A[3][18] * mat_B[18][30] +
                  mat_A[3][19] * mat_B[19][30] +
                  mat_A[3][20] * mat_B[20][30] +
                  mat_A[3][21] * mat_B[21][30] +
                  mat_A[3][22] * mat_B[22][30] +
                  mat_A[3][23] * mat_B[23][30] +
                  mat_A[3][24] * mat_B[24][30] +
                  mat_A[3][25] * mat_B[25][30] +
                  mat_A[3][26] * mat_B[26][30] +
                  mat_A[3][27] * mat_B[27][30] +
                  mat_A[3][28] * mat_B[28][30] +
                  mat_A[3][29] * mat_B[29][30] +
                  mat_A[3][30] * mat_B[30][30] +
                  mat_A[3][31] * mat_B[31][30];
    mat_C[3][31] <= 
                  mat_A[3][0] * mat_B[0][31] +
                  mat_A[3][1] * mat_B[1][31] +
                  mat_A[3][2] * mat_B[2][31] +
                  mat_A[3][3] * mat_B[3][31] +
                  mat_A[3][4] * mat_B[4][31] +
                  mat_A[3][5] * mat_B[5][31] +
                  mat_A[3][6] * mat_B[6][31] +
                  mat_A[3][7] * mat_B[7][31] +
                  mat_A[3][8] * mat_B[8][31] +
                  mat_A[3][9] * mat_B[9][31] +
                  mat_A[3][10] * mat_B[10][31] +
                  mat_A[3][11] * mat_B[11][31] +
                  mat_A[3][12] * mat_B[12][31] +
                  mat_A[3][13] * mat_B[13][31] +
                  mat_A[3][14] * mat_B[14][31] +
                  mat_A[3][15] * mat_B[15][31] +
                  mat_A[3][16] * mat_B[16][31] +
                  mat_A[3][17] * mat_B[17][31] +
                  mat_A[3][18] * mat_B[18][31] +
                  mat_A[3][19] * mat_B[19][31] +
                  mat_A[3][20] * mat_B[20][31] +
                  mat_A[3][21] * mat_B[21][31] +
                  mat_A[3][22] * mat_B[22][31] +
                  mat_A[3][23] * mat_B[23][31] +
                  mat_A[3][24] * mat_B[24][31] +
                  mat_A[3][25] * mat_B[25][31] +
                  mat_A[3][26] * mat_B[26][31] +
                  mat_A[3][27] * mat_B[27][31] +
                  mat_A[3][28] * mat_B[28][31] +
                  mat_A[3][29] * mat_B[29][31] +
                  mat_A[3][30] * mat_B[30][31] +
                  mat_A[3][31] * mat_B[31][31];
    mat_C[4][0] <= 
                  mat_A[4][0] * mat_B[0][0] +
                  mat_A[4][1] * mat_B[1][0] +
                  mat_A[4][2] * mat_B[2][0] +
                  mat_A[4][3] * mat_B[3][0] +
                  mat_A[4][4] * mat_B[4][0] +
                  mat_A[4][5] * mat_B[5][0] +
                  mat_A[4][6] * mat_B[6][0] +
                  mat_A[4][7] * mat_B[7][0] +
                  mat_A[4][8] * mat_B[8][0] +
                  mat_A[4][9] * mat_B[9][0] +
                  mat_A[4][10] * mat_B[10][0] +
                  mat_A[4][11] * mat_B[11][0] +
                  mat_A[4][12] * mat_B[12][0] +
                  mat_A[4][13] * mat_B[13][0] +
                  mat_A[4][14] * mat_B[14][0] +
                  mat_A[4][15] * mat_B[15][0] +
                  mat_A[4][16] * mat_B[16][0] +
                  mat_A[4][17] * mat_B[17][0] +
                  mat_A[4][18] * mat_B[18][0] +
                  mat_A[4][19] * mat_B[19][0] +
                  mat_A[4][20] * mat_B[20][0] +
                  mat_A[4][21] * mat_B[21][0] +
                  mat_A[4][22] * mat_B[22][0] +
                  mat_A[4][23] * mat_B[23][0] +
                  mat_A[4][24] * mat_B[24][0] +
                  mat_A[4][25] * mat_B[25][0] +
                  mat_A[4][26] * mat_B[26][0] +
                  mat_A[4][27] * mat_B[27][0] +
                  mat_A[4][28] * mat_B[28][0] +
                  mat_A[4][29] * mat_B[29][0] +
                  mat_A[4][30] * mat_B[30][0] +
                  mat_A[4][31] * mat_B[31][0];
    mat_C[4][1] <= 
                  mat_A[4][0] * mat_B[0][1] +
                  mat_A[4][1] * mat_B[1][1] +
                  mat_A[4][2] * mat_B[2][1] +
                  mat_A[4][3] * mat_B[3][1] +
                  mat_A[4][4] * mat_B[4][1] +
                  mat_A[4][5] * mat_B[5][1] +
                  mat_A[4][6] * mat_B[6][1] +
                  mat_A[4][7] * mat_B[7][1] +
                  mat_A[4][8] * mat_B[8][1] +
                  mat_A[4][9] * mat_B[9][1] +
                  mat_A[4][10] * mat_B[10][1] +
                  mat_A[4][11] * mat_B[11][1] +
                  mat_A[4][12] * mat_B[12][1] +
                  mat_A[4][13] * mat_B[13][1] +
                  mat_A[4][14] * mat_B[14][1] +
                  mat_A[4][15] * mat_B[15][1] +
                  mat_A[4][16] * mat_B[16][1] +
                  mat_A[4][17] * mat_B[17][1] +
                  mat_A[4][18] * mat_B[18][1] +
                  mat_A[4][19] * mat_B[19][1] +
                  mat_A[4][20] * mat_B[20][1] +
                  mat_A[4][21] * mat_B[21][1] +
                  mat_A[4][22] * mat_B[22][1] +
                  mat_A[4][23] * mat_B[23][1] +
                  mat_A[4][24] * mat_B[24][1] +
                  mat_A[4][25] * mat_B[25][1] +
                  mat_A[4][26] * mat_B[26][1] +
                  mat_A[4][27] * mat_B[27][1] +
                  mat_A[4][28] * mat_B[28][1] +
                  mat_A[4][29] * mat_B[29][1] +
                  mat_A[4][30] * mat_B[30][1] +
                  mat_A[4][31] * mat_B[31][1];
    mat_C[4][2] <= 
                  mat_A[4][0] * mat_B[0][2] +
                  mat_A[4][1] * mat_B[1][2] +
                  mat_A[4][2] * mat_B[2][2] +
                  mat_A[4][3] * mat_B[3][2] +
                  mat_A[4][4] * mat_B[4][2] +
                  mat_A[4][5] * mat_B[5][2] +
                  mat_A[4][6] * mat_B[6][2] +
                  mat_A[4][7] * mat_B[7][2] +
                  mat_A[4][8] * mat_B[8][2] +
                  mat_A[4][9] * mat_B[9][2] +
                  mat_A[4][10] * mat_B[10][2] +
                  mat_A[4][11] * mat_B[11][2] +
                  mat_A[4][12] * mat_B[12][2] +
                  mat_A[4][13] * mat_B[13][2] +
                  mat_A[4][14] * mat_B[14][2] +
                  mat_A[4][15] * mat_B[15][2] +
                  mat_A[4][16] * mat_B[16][2] +
                  mat_A[4][17] * mat_B[17][2] +
                  mat_A[4][18] * mat_B[18][2] +
                  mat_A[4][19] * mat_B[19][2] +
                  mat_A[4][20] * mat_B[20][2] +
                  mat_A[4][21] * mat_B[21][2] +
                  mat_A[4][22] * mat_B[22][2] +
                  mat_A[4][23] * mat_B[23][2] +
                  mat_A[4][24] * mat_B[24][2] +
                  mat_A[4][25] * mat_B[25][2] +
                  mat_A[4][26] * mat_B[26][2] +
                  mat_A[4][27] * mat_B[27][2] +
                  mat_A[4][28] * mat_B[28][2] +
                  mat_A[4][29] * mat_B[29][2] +
                  mat_A[4][30] * mat_B[30][2] +
                  mat_A[4][31] * mat_B[31][2];
    mat_C[4][3] <= 
                  mat_A[4][0] * mat_B[0][3] +
                  mat_A[4][1] * mat_B[1][3] +
                  mat_A[4][2] * mat_B[2][3] +
                  mat_A[4][3] * mat_B[3][3] +
                  mat_A[4][4] * mat_B[4][3] +
                  mat_A[4][5] * mat_B[5][3] +
                  mat_A[4][6] * mat_B[6][3] +
                  mat_A[4][7] * mat_B[7][3] +
                  mat_A[4][8] * mat_B[8][3] +
                  mat_A[4][9] * mat_B[9][3] +
                  mat_A[4][10] * mat_B[10][3] +
                  mat_A[4][11] * mat_B[11][3] +
                  mat_A[4][12] * mat_B[12][3] +
                  mat_A[4][13] * mat_B[13][3] +
                  mat_A[4][14] * mat_B[14][3] +
                  mat_A[4][15] * mat_B[15][3] +
                  mat_A[4][16] * mat_B[16][3] +
                  mat_A[4][17] * mat_B[17][3] +
                  mat_A[4][18] * mat_B[18][3] +
                  mat_A[4][19] * mat_B[19][3] +
                  mat_A[4][20] * mat_B[20][3] +
                  mat_A[4][21] * mat_B[21][3] +
                  mat_A[4][22] * mat_B[22][3] +
                  mat_A[4][23] * mat_B[23][3] +
                  mat_A[4][24] * mat_B[24][3] +
                  mat_A[4][25] * mat_B[25][3] +
                  mat_A[4][26] * mat_B[26][3] +
                  mat_A[4][27] * mat_B[27][3] +
                  mat_A[4][28] * mat_B[28][3] +
                  mat_A[4][29] * mat_B[29][3] +
                  mat_A[4][30] * mat_B[30][3] +
                  mat_A[4][31] * mat_B[31][3];
    mat_C[4][4] <= 
                  mat_A[4][0] * mat_B[0][4] +
                  mat_A[4][1] * mat_B[1][4] +
                  mat_A[4][2] * mat_B[2][4] +
                  mat_A[4][3] * mat_B[3][4] +
                  mat_A[4][4] * mat_B[4][4] +
                  mat_A[4][5] * mat_B[5][4] +
                  mat_A[4][6] * mat_B[6][4] +
                  mat_A[4][7] * mat_B[7][4] +
                  mat_A[4][8] * mat_B[8][4] +
                  mat_A[4][9] * mat_B[9][4] +
                  mat_A[4][10] * mat_B[10][4] +
                  mat_A[4][11] * mat_B[11][4] +
                  mat_A[4][12] * mat_B[12][4] +
                  mat_A[4][13] * mat_B[13][4] +
                  mat_A[4][14] * mat_B[14][4] +
                  mat_A[4][15] * mat_B[15][4] +
                  mat_A[4][16] * mat_B[16][4] +
                  mat_A[4][17] * mat_B[17][4] +
                  mat_A[4][18] * mat_B[18][4] +
                  mat_A[4][19] * mat_B[19][4] +
                  mat_A[4][20] * mat_B[20][4] +
                  mat_A[4][21] * mat_B[21][4] +
                  mat_A[4][22] * mat_B[22][4] +
                  mat_A[4][23] * mat_B[23][4] +
                  mat_A[4][24] * mat_B[24][4] +
                  mat_A[4][25] * mat_B[25][4] +
                  mat_A[4][26] * mat_B[26][4] +
                  mat_A[4][27] * mat_B[27][4] +
                  mat_A[4][28] * mat_B[28][4] +
                  mat_A[4][29] * mat_B[29][4] +
                  mat_A[4][30] * mat_B[30][4] +
                  mat_A[4][31] * mat_B[31][4];
    mat_C[4][5] <= 
                  mat_A[4][0] * mat_B[0][5] +
                  mat_A[4][1] * mat_B[1][5] +
                  mat_A[4][2] * mat_B[2][5] +
                  mat_A[4][3] * mat_B[3][5] +
                  mat_A[4][4] * mat_B[4][5] +
                  mat_A[4][5] * mat_B[5][5] +
                  mat_A[4][6] * mat_B[6][5] +
                  mat_A[4][7] * mat_B[7][5] +
                  mat_A[4][8] * mat_B[8][5] +
                  mat_A[4][9] * mat_B[9][5] +
                  mat_A[4][10] * mat_B[10][5] +
                  mat_A[4][11] * mat_B[11][5] +
                  mat_A[4][12] * mat_B[12][5] +
                  mat_A[4][13] * mat_B[13][5] +
                  mat_A[4][14] * mat_B[14][5] +
                  mat_A[4][15] * mat_B[15][5] +
                  mat_A[4][16] * mat_B[16][5] +
                  mat_A[4][17] * mat_B[17][5] +
                  mat_A[4][18] * mat_B[18][5] +
                  mat_A[4][19] * mat_B[19][5] +
                  mat_A[4][20] * mat_B[20][5] +
                  mat_A[4][21] * mat_B[21][5] +
                  mat_A[4][22] * mat_B[22][5] +
                  mat_A[4][23] * mat_B[23][5] +
                  mat_A[4][24] * mat_B[24][5] +
                  mat_A[4][25] * mat_B[25][5] +
                  mat_A[4][26] * mat_B[26][5] +
                  mat_A[4][27] * mat_B[27][5] +
                  mat_A[4][28] * mat_B[28][5] +
                  mat_A[4][29] * mat_B[29][5] +
                  mat_A[4][30] * mat_B[30][5] +
                  mat_A[4][31] * mat_B[31][5];
    mat_C[4][6] <= 
                  mat_A[4][0] * mat_B[0][6] +
                  mat_A[4][1] * mat_B[1][6] +
                  mat_A[4][2] * mat_B[2][6] +
                  mat_A[4][3] * mat_B[3][6] +
                  mat_A[4][4] * mat_B[4][6] +
                  mat_A[4][5] * mat_B[5][6] +
                  mat_A[4][6] * mat_B[6][6] +
                  mat_A[4][7] * mat_B[7][6] +
                  mat_A[4][8] * mat_B[8][6] +
                  mat_A[4][9] * mat_B[9][6] +
                  mat_A[4][10] * mat_B[10][6] +
                  mat_A[4][11] * mat_B[11][6] +
                  mat_A[4][12] * mat_B[12][6] +
                  mat_A[4][13] * mat_B[13][6] +
                  mat_A[4][14] * mat_B[14][6] +
                  mat_A[4][15] * mat_B[15][6] +
                  mat_A[4][16] * mat_B[16][6] +
                  mat_A[4][17] * mat_B[17][6] +
                  mat_A[4][18] * mat_B[18][6] +
                  mat_A[4][19] * mat_B[19][6] +
                  mat_A[4][20] * mat_B[20][6] +
                  mat_A[4][21] * mat_B[21][6] +
                  mat_A[4][22] * mat_B[22][6] +
                  mat_A[4][23] * mat_B[23][6] +
                  mat_A[4][24] * mat_B[24][6] +
                  mat_A[4][25] * mat_B[25][6] +
                  mat_A[4][26] * mat_B[26][6] +
                  mat_A[4][27] * mat_B[27][6] +
                  mat_A[4][28] * mat_B[28][6] +
                  mat_A[4][29] * mat_B[29][6] +
                  mat_A[4][30] * mat_B[30][6] +
                  mat_A[4][31] * mat_B[31][6];
    mat_C[4][7] <= 
                  mat_A[4][0] * mat_B[0][7] +
                  mat_A[4][1] * mat_B[1][7] +
                  mat_A[4][2] * mat_B[2][7] +
                  mat_A[4][3] * mat_B[3][7] +
                  mat_A[4][4] * mat_B[4][7] +
                  mat_A[4][5] * mat_B[5][7] +
                  mat_A[4][6] * mat_B[6][7] +
                  mat_A[4][7] * mat_B[7][7] +
                  mat_A[4][8] * mat_B[8][7] +
                  mat_A[4][9] * mat_B[9][7] +
                  mat_A[4][10] * mat_B[10][7] +
                  mat_A[4][11] * mat_B[11][7] +
                  mat_A[4][12] * mat_B[12][7] +
                  mat_A[4][13] * mat_B[13][7] +
                  mat_A[4][14] * mat_B[14][7] +
                  mat_A[4][15] * mat_B[15][7] +
                  mat_A[4][16] * mat_B[16][7] +
                  mat_A[4][17] * mat_B[17][7] +
                  mat_A[4][18] * mat_B[18][7] +
                  mat_A[4][19] * mat_B[19][7] +
                  mat_A[4][20] * mat_B[20][7] +
                  mat_A[4][21] * mat_B[21][7] +
                  mat_A[4][22] * mat_B[22][7] +
                  mat_A[4][23] * mat_B[23][7] +
                  mat_A[4][24] * mat_B[24][7] +
                  mat_A[4][25] * mat_B[25][7] +
                  mat_A[4][26] * mat_B[26][7] +
                  mat_A[4][27] * mat_B[27][7] +
                  mat_A[4][28] * mat_B[28][7] +
                  mat_A[4][29] * mat_B[29][7] +
                  mat_A[4][30] * mat_B[30][7] +
                  mat_A[4][31] * mat_B[31][7];
    mat_C[4][8] <= 
                  mat_A[4][0] * mat_B[0][8] +
                  mat_A[4][1] * mat_B[1][8] +
                  mat_A[4][2] * mat_B[2][8] +
                  mat_A[4][3] * mat_B[3][8] +
                  mat_A[4][4] * mat_B[4][8] +
                  mat_A[4][5] * mat_B[5][8] +
                  mat_A[4][6] * mat_B[6][8] +
                  mat_A[4][7] * mat_B[7][8] +
                  mat_A[4][8] * mat_B[8][8] +
                  mat_A[4][9] * mat_B[9][8] +
                  mat_A[4][10] * mat_B[10][8] +
                  mat_A[4][11] * mat_B[11][8] +
                  mat_A[4][12] * mat_B[12][8] +
                  mat_A[4][13] * mat_B[13][8] +
                  mat_A[4][14] * mat_B[14][8] +
                  mat_A[4][15] * mat_B[15][8] +
                  mat_A[4][16] * mat_B[16][8] +
                  mat_A[4][17] * mat_B[17][8] +
                  mat_A[4][18] * mat_B[18][8] +
                  mat_A[4][19] * mat_B[19][8] +
                  mat_A[4][20] * mat_B[20][8] +
                  mat_A[4][21] * mat_B[21][8] +
                  mat_A[4][22] * mat_B[22][8] +
                  mat_A[4][23] * mat_B[23][8] +
                  mat_A[4][24] * mat_B[24][8] +
                  mat_A[4][25] * mat_B[25][8] +
                  mat_A[4][26] * mat_B[26][8] +
                  mat_A[4][27] * mat_B[27][8] +
                  mat_A[4][28] * mat_B[28][8] +
                  mat_A[4][29] * mat_B[29][8] +
                  mat_A[4][30] * mat_B[30][8] +
                  mat_A[4][31] * mat_B[31][8];
    mat_C[4][9] <= 
                  mat_A[4][0] * mat_B[0][9] +
                  mat_A[4][1] * mat_B[1][9] +
                  mat_A[4][2] * mat_B[2][9] +
                  mat_A[4][3] * mat_B[3][9] +
                  mat_A[4][4] * mat_B[4][9] +
                  mat_A[4][5] * mat_B[5][9] +
                  mat_A[4][6] * mat_B[6][9] +
                  mat_A[4][7] * mat_B[7][9] +
                  mat_A[4][8] * mat_B[8][9] +
                  mat_A[4][9] * mat_B[9][9] +
                  mat_A[4][10] * mat_B[10][9] +
                  mat_A[4][11] * mat_B[11][9] +
                  mat_A[4][12] * mat_B[12][9] +
                  mat_A[4][13] * mat_B[13][9] +
                  mat_A[4][14] * mat_B[14][9] +
                  mat_A[4][15] * mat_B[15][9] +
                  mat_A[4][16] * mat_B[16][9] +
                  mat_A[4][17] * mat_B[17][9] +
                  mat_A[4][18] * mat_B[18][9] +
                  mat_A[4][19] * mat_B[19][9] +
                  mat_A[4][20] * mat_B[20][9] +
                  mat_A[4][21] * mat_B[21][9] +
                  mat_A[4][22] * mat_B[22][9] +
                  mat_A[4][23] * mat_B[23][9] +
                  mat_A[4][24] * mat_B[24][9] +
                  mat_A[4][25] * mat_B[25][9] +
                  mat_A[4][26] * mat_B[26][9] +
                  mat_A[4][27] * mat_B[27][9] +
                  mat_A[4][28] * mat_B[28][9] +
                  mat_A[4][29] * mat_B[29][9] +
                  mat_A[4][30] * mat_B[30][9] +
                  mat_A[4][31] * mat_B[31][9];
    mat_C[4][10] <= 
                  mat_A[4][0] * mat_B[0][10] +
                  mat_A[4][1] * mat_B[1][10] +
                  mat_A[4][2] * mat_B[2][10] +
                  mat_A[4][3] * mat_B[3][10] +
                  mat_A[4][4] * mat_B[4][10] +
                  mat_A[4][5] * mat_B[5][10] +
                  mat_A[4][6] * mat_B[6][10] +
                  mat_A[4][7] * mat_B[7][10] +
                  mat_A[4][8] * mat_B[8][10] +
                  mat_A[4][9] * mat_B[9][10] +
                  mat_A[4][10] * mat_B[10][10] +
                  mat_A[4][11] * mat_B[11][10] +
                  mat_A[4][12] * mat_B[12][10] +
                  mat_A[4][13] * mat_B[13][10] +
                  mat_A[4][14] * mat_B[14][10] +
                  mat_A[4][15] * mat_B[15][10] +
                  mat_A[4][16] * mat_B[16][10] +
                  mat_A[4][17] * mat_B[17][10] +
                  mat_A[4][18] * mat_B[18][10] +
                  mat_A[4][19] * mat_B[19][10] +
                  mat_A[4][20] * mat_B[20][10] +
                  mat_A[4][21] * mat_B[21][10] +
                  mat_A[4][22] * mat_B[22][10] +
                  mat_A[4][23] * mat_B[23][10] +
                  mat_A[4][24] * mat_B[24][10] +
                  mat_A[4][25] * mat_B[25][10] +
                  mat_A[4][26] * mat_B[26][10] +
                  mat_A[4][27] * mat_B[27][10] +
                  mat_A[4][28] * mat_B[28][10] +
                  mat_A[4][29] * mat_B[29][10] +
                  mat_A[4][30] * mat_B[30][10] +
                  mat_A[4][31] * mat_B[31][10];
    mat_C[4][11] <= 
                  mat_A[4][0] * mat_B[0][11] +
                  mat_A[4][1] * mat_B[1][11] +
                  mat_A[4][2] * mat_B[2][11] +
                  mat_A[4][3] * mat_B[3][11] +
                  mat_A[4][4] * mat_B[4][11] +
                  mat_A[4][5] * mat_B[5][11] +
                  mat_A[4][6] * mat_B[6][11] +
                  mat_A[4][7] * mat_B[7][11] +
                  mat_A[4][8] * mat_B[8][11] +
                  mat_A[4][9] * mat_B[9][11] +
                  mat_A[4][10] * mat_B[10][11] +
                  mat_A[4][11] * mat_B[11][11] +
                  mat_A[4][12] * mat_B[12][11] +
                  mat_A[4][13] * mat_B[13][11] +
                  mat_A[4][14] * mat_B[14][11] +
                  mat_A[4][15] * mat_B[15][11] +
                  mat_A[4][16] * mat_B[16][11] +
                  mat_A[4][17] * mat_B[17][11] +
                  mat_A[4][18] * mat_B[18][11] +
                  mat_A[4][19] * mat_B[19][11] +
                  mat_A[4][20] * mat_B[20][11] +
                  mat_A[4][21] * mat_B[21][11] +
                  mat_A[4][22] * mat_B[22][11] +
                  mat_A[4][23] * mat_B[23][11] +
                  mat_A[4][24] * mat_B[24][11] +
                  mat_A[4][25] * mat_B[25][11] +
                  mat_A[4][26] * mat_B[26][11] +
                  mat_A[4][27] * mat_B[27][11] +
                  mat_A[4][28] * mat_B[28][11] +
                  mat_A[4][29] * mat_B[29][11] +
                  mat_A[4][30] * mat_B[30][11] +
                  mat_A[4][31] * mat_B[31][11];
    mat_C[4][12] <= 
                  mat_A[4][0] * mat_B[0][12] +
                  mat_A[4][1] * mat_B[1][12] +
                  mat_A[4][2] * mat_B[2][12] +
                  mat_A[4][3] * mat_B[3][12] +
                  mat_A[4][4] * mat_B[4][12] +
                  mat_A[4][5] * mat_B[5][12] +
                  mat_A[4][6] * mat_B[6][12] +
                  mat_A[4][7] * mat_B[7][12] +
                  mat_A[4][8] * mat_B[8][12] +
                  mat_A[4][9] * mat_B[9][12] +
                  mat_A[4][10] * mat_B[10][12] +
                  mat_A[4][11] * mat_B[11][12] +
                  mat_A[4][12] * mat_B[12][12] +
                  mat_A[4][13] * mat_B[13][12] +
                  mat_A[4][14] * mat_B[14][12] +
                  mat_A[4][15] * mat_B[15][12] +
                  mat_A[4][16] * mat_B[16][12] +
                  mat_A[4][17] * mat_B[17][12] +
                  mat_A[4][18] * mat_B[18][12] +
                  mat_A[4][19] * mat_B[19][12] +
                  mat_A[4][20] * mat_B[20][12] +
                  mat_A[4][21] * mat_B[21][12] +
                  mat_A[4][22] * mat_B[22][12] +
                  mat_A[4][23] * mat_B[23][12] +
                  mat_A[4][24] * mat_B[24][12] +
                  mat_A[4][25] * mat_B[25][12] +
                  mat_A[4][26] * mat_B[26][12] +
                  mat_A[4][27] * mat_B[27][12] +
                  mat_A[4][28] * mat_B[28][12] +
                  mat_A[4][29] * mat_B[29][12] +
                  mat_A[4][30] * mat_B[30][12] +
                  mat_A[4][31] * mat_B[31][12];
    mat_C[4][13] <= 
                  mat_A[4][0] * mat_B[0][13] +
                  mat_A[4][1] * mat_B[1][13] +
                  mat_A[4][2] * mat_B[2][13] +
                  mat_A[4][3] * mat_B[3][13] +
                  mat_A[4][4] * mat_B[4][13] +
                  mat_A[4][5] * mat_B[5][13] +
                  mat_A[4][6] * mat_B[6][13] +
                  mat_A[4][7] * mat_B[7][13] +
                  mat_A[4][8] * mat_B[8][13] +
                  mat_A[4][9] * mat_B[9][13] +
                  mat_A[4][10] * mat_B[10][13] +
                  mat_A[4][11] * mat_B[11][13] +
                  mat_A[4][12] * mat_B[12][13] +
                  mat_A[4][13] * mat_B[13][13] +
                  mat_A[4][14] * mat_B[14][13] +
                  mat_A[4][15] * mat_B[15][13] +
                  mat_A[4][16] * mat_B[16][13] +
                  mat_A[4][17] * mat_B[17][13] +
                  mat_A[4][18] * mat_B[18][13] +
                  mat_A[4][19] * mat_B[19][13] +
                  mat_A[4][20] * mat_B[20][13] +
                  mat_A[4][21] * mat_B[21][13] +
                  mat_A[4][22] * mat_B[22][13] +
                  mat_A[4][23] * mat_B[23][13] +
                  mat_A[4][24] * mat_B[24][13] +
                  mat_A[4][25] * mat_B[25][13] +
                  mat_A[4][26] * mat_B[26][13] +
                  mat_A[4][27] * mat_B[27][13] +
                  mat_A[4][28] * mat_B[28][13] +
                  mat_A[4][29] * mat_B[29][13] +
                  mat_A[4][30] * mat_B[30][13] +
                  mat_A[4][31] * mat_B[31][13];
    mat_C[4][14] <= 
                  mat_A[4][0] * mat_B[0][14] +
                  mat_A[4][1] * mat_B[1][14] +
                  mat_A[4][2] * mat_B[2][14] +
                  mat_A[4][3] * mat_B[3][14] +
                  mat_A[4][4] * mat_B[4][14] +
                  mat_A[4][5] * mat_B[5][14] +
                  mat_A[4][6] * mat_B[6][14] +
                  mat_A[4][7] * mat_B[7][14] +
                  mat_A[4][8] * mat_B[8][14] +
                  mat_A[4][9] * mat_B[9][14] +
                  mat_A[4][10] * mat_B[10][14] +
                  mat_A[4][11] * mat_B[11][14] +
                  mat_A[4][12] * mat_B[12][14] +
                  mat_A[4][13] * mat_B[13][14] +
                  mat_A[4][14] * mat_B[14][14] +
                  mat_A[4][15] * mat_B[15][14] +
                  mat_A[4][16] * mat_B[16][14] +
                  mat_A[4][17] * mat_B[17][14] +
                  mat_A[4][18] * mat_B[18][14] +
                  mat_A[4][19] * mat_B[19][14] +
                  mat_A[4][20] * mat_B[20][14] +
                  mat_A[4][21] * mat_B[21][14] +
                  mat_A[4][22] * mat_B[22][14] +
                  mat_A[4][23] * mat_B[23][14] +
                  mat_A[4][24] * mat_B[24][14] +
                  mat_A[4][25] * mat_B[25][14] +
                  mat_A[4][26] * mat_B[26][14] +
                  mat_A[4][27] * mat_B[27][14] +
                  mat_A[4][28] * mat_B[28][14] +
                  mat_A[4][29] * mat_B[29][14] +
                  mat_A[4][30] * mat_B[30][14] +
                  mat_A[4][31] * mat_B[31][14];
    mat_C[4][15] <= 
                  mat_A[4][0] * mat_B[0][15] +
                  mat_A[4][1] * mat_B[1][15] +
                  mat_A[4][2] * mat_B[2][15] +
                  mat_A[4][3] * mat_B[3][15] +
                  mat_A[4][4] * mat_B[4][15] +
                  mat_A[4][5] * mat_B[5][15] +
                  mat_A[4][6] * mat_B[6][15] +
                  mat_A[4][7] * mat_B[7][15] +
                  mat_A[4][8] * mat_B[8][15] +
                  mat_A[4][9] * mat_B[9][15] +
                  mat_A[4][10] * mat_B[10][15] +
                  mat_A[4][11] * mat_B[11][15] +
                  mat_A[4][12] * mat_B[12][15] +
                  mat_A[4][13] * mat_B[13][15] +
                  mat_A[4][14] * mat_B[14][15] +
                  mat_A[4][15] * mat_B[15][15] +
                  mat_A[4][16] * mat_B[16][15] +
                  mat_A[4][17] * mat_B[17][15] +
                  mat_A[4][18] * mat_B[18][15] +
                  mat_A[4][19] * mat_B[19][15] +
                  mat_A[4][20] * mat_B[20][15] +
                  mat_A[4][21] * mat_B[21][15] +
                  mat_A[4][22] * mat_B[22][15] +
                  mat_A[4][23] * mat_B[23][15] +
                  mat_A[4][24] * mat_B[24][15] +
                  mat_A[4][25] * mat_B[25][15] +
                  mat_A[4][26] * mat_B[26][15] +
                  mat_A[4][27] * mat_B[27][15] +
                  mat_A[4][28] * mat_B[28][15] +
                  mat_A[4][29] * mat_B[29][15] +
                  mat_A[4][30] * mat_B[30][15] +
                  mat_A[4][31] * mat_B[31][15];
    mat_C[4][16] <= 
                  mat_A[4][0] * mat_B[0][16] +
                  mat_A[4][1] * mat_B[1][16] +
                  mat_A[4][2] * mat_B[2][16] +
                  mat_A[4][3] * mat_B[3][16] +
                  mat_A[4][4] * mat_B[4][16] +
                  mat_A[4][5] * mat_B[5][16] +
                  mat_A[4][6] * mat_B[6][16] +
                  mat_A[4][7] * mat_B[7][16] +
                  mat_A[4][8] * mat_B[8][16] +
                  mat_A[4][9] * mat_B[9][16] +
                  mat_A[4][10] * mat_B[10][16] +
                  mat_A[4][11] * mat_B[11][16] +
                  mat_A[4][12] * mat_B[12][16] +
                  mat_A[4][13] * mat_B[13][16] +
                  mat_A[4][14] * mat_B[14][16] +
                  mat_A[4][15] * mat_B[15][16] +
                  mat_A[4][16] * mat_B[16][16] +
                  mat_A[4][17] * mat_B[17][16] +
                  mat_A[4][18] * mat_B[18][16] +
                  mat_A[4][19] * mat_B[19][16] +
                  mat_A[4][20] * mat_B[20][16] +
                  mat_A[4][21] * mat_B[21][16] +
                  mat_A[4][22] * mat_B[22][16] +
                  mat_A[4][23] * mat_B[23][16] +
                  mat_A[4][24] * mat_B[24][16] +
                  mat_A[4][25] * mat_B[25][16] +
                  mat_A[4][26] * mat_B[26][16] +
                  mat_A[4][27] * mat_B[27][16] +
                  mat_A[4][28] * mat_B[28][16] +
                  mat_A[4][29] * mat_B[29][16] +
                  mat_A[4][30] * mat_B[30][16] +
                  mat_A[4][31] * mat_B[31][16];
    mat_C[4][17] <= 
                  mat_A[4][0] * mat_B[0][17] +
                  mat_A[4][1] * mat_B[1][17] +
                  mat_A[4][2] * mat_B[2][17] +
                  mat_A[4][3] * mat_B[3][17] +
                  mat_A[4][4] * mat_B[4][17] +
                  mat_A[4][5] * mat_B[5][17] +
                  mat_A[4][6] * mat_B[6][17] +
                  mat_A[4][7] * mat_B[7][17] +
                  mat_A[4][8] * mat_B[8][17] +
                  mat_A[4][9] * mat_B[9][17] +
                  mat_A[4][10] * mat_B[10][17] +
                  mat_A[4][11] * mat_B[11][17] +
                  mat_A[4][12] * mat_B[12][17] +
                  mat_A[4][13] * mat_B[13][17] +
                  mat_A[4][14] * mat_B[14][17] +
                  mat_A[4][15] * mat_B[15][17] +
                  mat_A[4][16] * mat_B[16][17] +
                  mat_A[4][17] * mat_B[17][17] +
                  mat_A[4][18] * mat_B[18][17] +
                  mat_A[4][19] * mat_B[19][17] +
                  mat_A[4][20] * mat_B[20][17] +
                  mat_A[4][21] * mat_B[21][17] +
                  mat_A[4][22] * mat_B[22][17] +
                  mat_A[4][23] * mat_B[23][17] +
                  mat_A[4][24] * mat_B[24][17] +
                  mat_A[4][25] * mat_B[25][17] +
                  mat_A[4][26] * mat_B[26][17] +
                  mat_A[4][27] * mat_B[27][17] +
                  mat_A[4][28] * mat_B[28][17] +
                  mat_A[4][29] * mat_B[29][17] +
                  mat_A[4][30] * mat_B[30][17] +
                  mat_A[4][31] * mat_B[31][17];
    mat_C[4][18] <= 
                  mat_A[4][0] * mat_B[0][18] +
                  mat_A[4][1] * mat_B[1][18] +
                  mat_A[4][2] * mat_B[2][18] +
                  mat_A[4][3] * mat_B[3][18] +
                  mat_A[4][4] * mat_B[4][18] +
                  mat_A[4][5] * mat_B[5][18] +
                  mat_A[4][6] * mat_B[6][18] +
                  mat_A[4][7] * mat_B[7][18] +
                  mat_A[4][8] * mat_B[8][18] +
                  mat_A[4][9] * mat_B[9][18] +
                  mat_A[4][10] * mat_B[10][18] +
                  mat_A[4][11] * mat_B[11][18] +
                  mat_A[4][12] * mat_B[12][18] +
                  mat_A[4][13] * mat_B[13][18] +
                  mat_A[4][14] * mat_B[14][18] +
                  mat_A[4][15] * mat_B[15][18] +
                  mat_A[4][16] * mat_B[16][18] +
                  mat_A[4][17] * mat_B[17][18] +
                  mat_A[4][18] * mat_B[18][18] +
                  mat_A[4][19] * mat_B[19][18] +
                  mat_A[4][20] * mat_B[20][18] +
                  mat_A[4][21] * mat_B[21][18] +
                  mat_A[4][22] * mat_B[22][18] +
                  mat_A[4][23] * mat_B[23][18] +
                  mat_A[4][24] * mat_B[24][18] +
                  mat_A[4][25] * mat_B[25][18] +
                  mat_A[4][26] * mat_B[26][18] +
                  mat_A[4][27] * mat_B[27][18] +
                  mat_A[4][28] * mat_B[28][18] +
                  mat_A[4][29] * mat_B[29][18] +
                  mat_A[4][30] * mat_B[30][18] +
                  mat_A[4][31] * mat_B[31][18];
    mat_C[4][19] <= 
                  mat_A[4][0] * mat_B[0][19] +
                  mat_A[4][1] * mat_B[1][19] +
                  mat_A[4][2] * mat_B[2][19] +
                  mat_A[4][3] * mat_B[3][19] +
                  mat_A[4][4] * mat_B[4][19] +
                  mat_A[4][5] * mat_B[5][19] +
                  mat_A[4][6] * mat_B[6][19] +
                  mat_A[4][7] * mat_B[7][19] +
                  mat_A[4][8] * mat_B[8][19] +
                  mat_A[4][9] * mat_B[9][19] +
                  mat_A[4][10] * mat_B[10][19] +
                  mat_A[4][11] * mat_B[11][19] +
                  mat_A[4][12] * mat_B[12][19] +
                  mat_A[4][13] * mat_B[13][19] +
                  mat_A[4][14] * mat_B[14][19] +
                  mat_A[4][15] * mat_B[15][19] +
                  mat_A[4][16] * mat_B[16][19] +
                  mat_A[4][17] * mat_B[17][19] +
                  mat_A[4][18] * mat_B[18][19] +
                  mat_A[4][19] * mat_B[19][19] +
                  mat_A[4][20] * mat_B[20][19] +
                  mat_A[4][21] * mat_B[21][19] +
                  mat_A[4][22] * mat_B[22][19] +
                  mat_A[4][23] * mat_B[23][19] +
                  mat_A[4][24] * mat_B[24][19] +
                  mat_A[4][25] * mat_B[25][19] +
                  mat_A[4][26] * mat_B[26][19] +
                  mat_A[4][27] * mat_B[27][19] +
                  mat_A[4][28] * mat_B[28][19] +
                  mat_A[4][29] * mat_B[29][19] +
                  mat_A[4][30] * mat_B[30][19] +
                  mat_A[4][31] * mat_B[31][19];
    mat_C[4][20] <= 
                  mat_A[4][0] * mat_B[0][20] +
                  mat_A[4][1] * mat_B[1][20] +
                  mat_A[4][2] * mat_B[2][20] +
                  mat_A[4][3] * mat_B[3][20] +
                  mat_A[4][4] * mat_B[4][20] +
                  mat_A[4][5] * mat_B[5][20] +
                  mat_A[4][6] * mat_B[6][20] +
                  mat_A[4][7] * mat_B[7][20] +
                  mat_A[4][8] * mat_B[8][20] +
                  mat_A[4][9] * mat_B[9][20] +
                  mat_A[4][10] * mat_B[10][20] +
                  mat_A[4][11] * mat_B[11][20] +
                  mat_A[4][12] * mat_B[12][20] +
                  mat_A[4][13] * mat_B[13][20] +
                  mat_A[4][14] * mat_B[14][20] +
                  mat_A[4][15] * mat_B[15][20] +
                  mat_A[4][16] * mat_B[16][20] +
                  mat_A[4][17] * mat_B[17][20] +
                  mat_A[4][18] * mat_B[18][20] +
                  mat_A[4][19] * mat_B[19][20] +
                  mat_A[4][20] * mat_B[20][20] +
                  mat_A[4][21] * mat_B[21][20] +
                  mat_A[4][22] * mat_B[22][20] +
                  mat_A[4][23] * mat_B[23][20] +
                  mat_A[4][24] * mat_B[24][20] +
                  mat_A[4][25] * mat_B[25][20] +
                  mat_A[4][26] * mat_B[26][20] +
                  mat_A[4][27] * mat_B[27][20] +
                  mat_A[4][28] * mat_B[28][20] +
                  mat_A[4][29] * mat_B[29][20] +
                  mat_A[4][30] * mat_B[30][20] +
                  mat_A[4][31] * mat_B[31][20];
    mat_C[4][21] <= 
                  mat_A[4][0] * mat_B[0][21] +
                  mat_A[4][1] * mat_B[1][21] +
                  mat_A[4][2] * mat_B[2][21] +
                  mat_A[4][3] * mat_B[3][21] +
                  mat_A[4][4] * mat_B[4][21] +
                  mat_A[4][5] * mat_B[5][21] +
                  mat_A[4][6] * mat_B[6][21] +
                  mat_A[4][7] * mat_B[7][21] +
                  mat_A[4][8] * mat_B[8][21] +
                  mat_A[4][9] * mat_B[9][21] +
                  mat_A[4][10] * mat_B[10][21] +
                  mat_A[4][11] * mat_B[11][21] +
                  mat_A[4][12] * mat_B[12][21] +
                  mat_A[4][13] * mat_B[13][21] +
                  mat_A[4][14] * mat_B[14][21] +
                  mat_A[4][15] * mat_B[15][21] +
                  mat_A[4][16] * mat_B[16][21] +
                  mat_A[4][17] * mat_B[17][21] +
                  mat_A[4][18] * mat_B[18][21] +
                  mat_A[4][19] * mat_B[19][21] +
                  mat_A[4][20] * mat_B[20][21] +
                  mat_A[4][21] * mat_B[21][21] +
                  mat_A[4][22] * mat_B[22][21] +
                  mat_A[4][23] * mat_B[23][21] +
                  mat_A[4][24] * mat_B[24][21] +
                  mat_A[4][25] * mat_B[25][21] +
                  mat_A[4][26] * mat_B[26][21] +
                  mat_A[4][27] * mat_B[27][21] +
                  mat_A[4][28] * mat_B[28][21] +
                  mat_A[4][29] * mat_B[29][21] +
                  mat_A[4][30] * mat_B[30][21] +
                  mat_A[4][31] * mat_B[31][21];
    mat_C[4][22] <= 
                  mat_A[4][0] * mat_B[0][22] +
                  mat_A[4][1] * mat_B[1][22] +
                  mat_A[4][2] * mat_B[2][22] +
                  mat_A[4][3] * mat_B[3][22] +
                  mat_A[4][4] * mat_B[4][22] +
                  mat_A[4][5] * mat_B[5][22] +
                  mat_A[4][6] * mat_B[6][22] +
                  mat_A[4][7] * mat_B[7][22] +
                  mat_A[4][8] * mat_B[8][22] +
                  mat_A[4][9] * mat_B[9][22] +
                  mat_A[4][10] * mat_B[10][22] +
                  mat_A[4][11] * mat_B[11][22] +
                  mat_A[4][12] * mat_B[12][22] +
                  mat_A[4][13] * mat_B[13][22] +
                  mat_A[4][14] * mat_B[14][22] +
                  mat_A[4][15] * mat_B[15][22] +
                  mat_A[4][16] * mat_B[16][22] +
                  mat_A[4][17] * mat_B[17][22] +
                  mat_A[4][18] * mat_B[18][22] +
                  mat_A[4][19] * mat_B[19][22] +
                  mat_A[4][20] * mat_B[20][22] +
                  mat_A[4][21] * mat_B[21][22] +
                  mat_A[4][22] * mat_B[22][22] +
                  mat_A[4][23] * mat_B[23][22] +
                  mat_A[4][24] * mat_B[24][22] +
                  mat_A[4][25] * mat_B[25][22] +
                  mat_A[4][26] * mat_B[26][22] +
                  mat_A[4][27] * mat_B[27][22] +
                  mat_A[4][28] * mat_B[28][22] +
                  mat_A[4][29] * mat_B[29][22] +
                  mat_A[4][30] * mat_B[30][22] +
                  mat_A[4][31] * mat_B[31][22];
    mat_C[4][23] <= 
                  mat_A[4][0] * mat_B[0][23] +
                  mat_A[4][1] * mat_B[1][23] +
                  mat_A[4][2] * mat_B[2][23] +
                  mat_A[4][3] * mat_B[3][23] +
                  mat_A[4][4] * mat_B[4][23] +
                  mat_A[4][5] * mat_B[5][23] +
                  mat_A[4][6] * mat_B[6][23] +
                  mat_A[4][7] * mat_B[7][23] +
                  mat_A[4][8] * mat_B[8][23] +
                  mat_A[4][9] * mat_B[9][23] +
                  mat_A[4][10] * mat_B[10][23] +
                  mat_A[4][11] * mat_B[11][23] +
                  mat_A[4][12] * mat_B[12][23] +
                  mat_A[4][13] * mat_B[13][23] +
                  mat_A[4][14] * mat_B[14][23] +
                  mat_A[4][15] * mat_B[15][23] +
                  mat_A[4][16] * mat_B[16][23] +
                  mat_A[4][17] * mat_B[17][23] +
                  mat_A[4][18] * mat_B[18][23] +
                  mat_A[4][19] * mat_B[19][23] +
                  mat_A[4][20] * mat_B[20][23] +
                  mat_A[4][21] * mat_B[21][23] +
                  mat_A[4][22] * mat_B[22][23] +
                  mat_A[4][23] * mat_B[23][23] +
                  mat_A[4][24] * mat_B[24][23] +
                  mat_A[4][25] * mat_B[25][23] +
                  mat_A[4][26] * mat_B[26][23] +
                  mat_A[4][27] * mat_B[27][23] +
                  mat_A[4][28] * mat_B[28][23] +
                  mat_A[4][29] * mat_B[29][23] +
                  mat_A[4][30] * mat_B[30][23] +
                  mat_A[4][31] * mat_B[31][23];
    mat_C[4][24] <= 
                  mat_A[4][0] * mat_B[0][24] +
                  mat_A[4][1] * mat_B[1][24] +
                  mat_A[4][2] * mat_B[2][24] +
                  mat_A[4][3] * mat_B[3][24] +
                  mat_A[4][4] * mat_B[4][24] +
                  mat_A[4][5] * mat_B[5][24] +
                  mat_A[4][6] * mat_B[6][24] +
                  mat_A[4][7] * mat_B[7][24] +
                  mat_A[4][8] * mat_B[8][24] +
                  mat_A[4][9] * mat_B[9][24] +
                  mat_A[4][10] * mat_B[10][24] +
                  mat_A[4][11] * mat_B[11][24] +
                  mat_A[4][12] * mat_B[12][24] +
                  mat_A[4][13] * mat_B[13][24] +
                  mat_A[4][14] * mat_B[14][24] +
                  mat_A[4][15] * mat_B[15][24] +
                  mat_A[4][16] * mat_B[16][24] +
                  mat_A[4][17] * mat_B[17][24] +
                  mat_A[4][18] * mat_B[18][24] +
                  mat_A[4][19] * mat_B[19][24] +
                  mat_A[4][20] * mat_B[20][24] +
                  mat_A[4][21] * mat_B[21][24] +
                  mat_A[4][22] * mat_B[22][24] +
                  mat_A[4][23] * mat_B[23][24] +
                  mat_A[4][24] * mat_B[24][24] +
                  mat_A[4][25] * mat_B[25][24] +
                  mat_A[4][26] * mat_B[26][24] +
                  mat_A[4][27] * mat_B[27][24] +
                  mat_A[4][28] * mat_B[28][24] +
                  mat_A[4][29] * mat_B[29][24] +
                  mat_A[4][30] * mat_B[30][24] +
                  mat_A[4][31] * mat_B[31][24];
    mat_C[4][25] <= 
                  mat_A[4][0] * mat_B[0][25] +
                  mat_A[4][1] * mat_B[1][25] +
                  mat_A[4][2] * mat_B[2][25] +
                  mat_A[4][3] * mat_B[3][25] +
                  mat_A[4][4] * mat_B[4][25] +
                  mat_A[4][5] * mat_B[5][25] +
                  mat_A[4][6] * mat_B[6][25] +
                  mat_A[4][7] * mat_B[7][25] +
                  mat_A[4][8] * mat_B[8][25] +
                  mat_A[4][9] * mat_B[9][25] +
                  mat_A[4][10] * mat_B[10][25] +
                  mat_A[4][11] * mat_B[11][25] +
                  mat_A[4][12] * mat_B[12][25] +
                  mat_A[4][13] * mat_B[13][25] +
                  mat_A[4][14] * mat_B[14][25] +
                  mat_A[4][15] * mat_B[15][25] +
                  mat_A[4][16] * mat_B[16][25] +
                  mat_A[4][17] * mat_B[17][25] +
                  mat_A[4][18] * mat_B[18][25] +
                  mat_A[4][19] * mat_B[19][25] +
                  mat_A[4][20] * mat_B[20][25] +
                  mat_A[4][21] * mat_B[21][25] +
                  mat_A[4][22] * mat_B[22][25] +
                  mat_A[4][23] * mat_B[23][25] +
                  mat_A[4][24] * mat_B[24][25] +
                  mat_A[4][25] * mat_B[25][25] +
                  mat_A[4][26] * mat_B[26][25] +
                  mat_A[4][27] * mat_B[27][25] +
                  mat_A[4][28] * mat_B[28][25] +
                  mat_A[4][29] * mat_B[29][25] +
                  mat_A[4][30] * mat_B[30][25] +
                  mat_A[4][31] * mat_B[31][25];
    mat_C[4][26] <= 
                  mat_A[4][0] * mat_B[0][26] +
                  mat_A[4][1] * mat_B[1][26] +
                  mat_A[4][2] * mat_B[2][26] +
                  mat_A[4][3] * mat_B[3][26] +
                  mat_A[4][4] * mat_B[4][26] +
                  mat_A[4][5] * mat_B[5][26] +
                  mat_A[4][6] * mat_B[6][26] +
                  mat_A[4][7] * mat_B[7][26] +
                  mat_A[4][8] * mat_B[8][26] +
                  mat_A[4][9] * mat_B[9][26] +
                  mat_A[4][10] * mat_B[10][26] +
                  mat_A[4][11] * mat_B[11][26] +
                  mat_A[4][12] * mat_B[12][26] +
                  mat_A[4][13] * mat_B[13][26] +
                  mat_A[4][14] * mat_B[14][26] +
                  mat_A[4][15] * mat_B[15][26] +
                  mat_A[4][16] * mat_B[16][26] +
                  mat_A[4][17] * mat_B[17][26] +
                  mat_A[4][18] * mat_B[18][26] +
                  mat_A[4][19] * mat_B[19][26] +
                  mat_A[4][20] * mat_B[20][26] +
                  mat_A[4][21] * mat_B[21][26] +
                  mat_A[4][22] * mat_B[22][26] +
                  mat_A[4][23] * mat_B[23][26] +
                  mat_A[4][24] * mat_B[24][26] +
                  mat_A[4][25] * mat_B[25][26] +
                  mat_A[4][26] * mat_B[26][26] +
                  mat_A[4][27] * mat_B[27][26] +
                  mat_A[4][28] * mat_B[28][26] +
                  mat_A[4][29] * mat_B[29][26] +
                  mat_A[4][30] * mat_B[30][26] +
                  mat_A[4][31] * mat_B[31][26];
    mat_C[4][27] <= 
                  mat_A[4][0] * mat_B[0][27] +
                  mat_A[4][1] * mat_B[1][27] +
                  mat_A[4][2] * mat_B[2][27] +
                  mat_A[4][3] * mat_B[3][27] +
                  mat_A[4][4] * mat_B[4][27] +
                  mat_A[4][5] * mat_B[5][27] +
                  mat_A[4][6] * mat_B[6][27] +
                  mat_A[4][7] * mat_B[7][27] +
                  mat_A[4][8] * mat_B[8][27] +
                  mat_A[4][9] * mat_B[9][27] +
                  mat_A[4][10] * mat_B[10][27] +
                  mat_A[4][11] * mat_B[11][27] +
                  mat_A[4][12] * mat_B[12][27] +
                  mat_A[4][13] * mat_B[13][27] +
                  mat_A[4][14] * mat_B[14][27] +
                  mat_A[4][15] * mat_B[15][27] +
                  mat_A[4][16] * mat_B[16][27] +
                  mat_A[4][17] * mat_B[17][27] +
                  mat_A[4][18] * mat_B[18][27] +
                  mat_A[4][19] * mat_B[19][27] +
                  mat_A[4][20] * mat_B[20][27] +
                  mat_A[4][21] * mat_B[21][27] +
                  mat_A[4][22] * mat_B[22][27] +
                  mat_A[4][23] * mat_B[23][27] +
                  mat_A[4][24] * mat_B[24][27] +
                  mat_A[4][25] * mat_B[25][27] +
                  mat_A[4][26] * mat_B[26][27] +
                  mat_A[4][27] * mat_B[27][27] +
                  mat_A[4][28] * mat_B[28][27] +
                  mat_A[4][29] * mat_B[29][27] +
                  mat_A[4][30] * mat_B[30][27] +
                  mat_A[4][31] * mat_B[31][27];
    mat_C[4][28] <= 
                  mat_A[4][0] * mat_B[0][28] +
                  mat_A[4][1] * mat_B[1][28] +
                  mat_A[4][2] * mat_B[2][28] +
                  mat_A[4][3] * mat_B[3][28] +
                  mat_A[4][4] * mat_B[4][28] +
                  mat_A[4][5] * mat_B[5][28] +
                  mat_A[4][6] * mat_B[6][28] +
                  mat_A[4][7] * mat_B[7][28] +
                  mat_A[4][8] * mat_B[8][28] +
                  mat_A[4][9] * mat_B[9][28] +
                  mat_A[4][10] * mat_B[10][28] +
                  mat_A[4][11] * mat_B[11][28] +
                  mat_A[4][12] * mat_B[12][28] +
                  mat_A[4][13] * mat_B[13][28] +
                  mat_A[4][14] * mat_B[14][28] +
                  mat_A[4][15] * mat_B[15][28] +
                  mat_A[4][16] * mat_B[16][28] +
                  mat_A[4][17] * mat_B[17][28] +
                  mat_A[4][18] * mat_B[18][28] +
                  mat_A[4][19] * mat_B[19][28] +
                  mat_A[4][20] * mat_B[20][28] +
                  mat_A[4][21] * mat_B[21][28] +
                  mat_A[4][22] * mat_B[22][28] +
                  mat_A[4][23] * mat_B[23][28] +
                  mat_A[4][24] * mat_B[24][28] +
                  mat_A[4][25] * mat_B[25][28] +
                  mat_A[4][26] * mat_B[26][28] +
                  mat_A[4][27] * mat_B[27][28] +
                  mat_A[4][28] * mat_B[28][28] +
                  mat_A[4][29] * mat_B[29][28] +
                  mat_A[4][30] * mat_B[30][28] +
                  mat_A[4][31] * mat_B[31][28];
    mat_C[4][29] <= 
                  mat_A[4][0] * mat_B[0][29] +
                  mat_A[4][1] * mat_B[1][29] +
                  mat_A[4][2] * mat_B[2][29] +
                  mat_A[4][3] * mat_B[3][29] +
                  mat_A[4][4] * mat_B[4][29] +
                  mat_A[4][5] * mat_B[5][29] +
                  mat_A[4][6] * mat_B[6][29] +
                  mat_A[4][7] * mat_B[7][29] +
                  mat_A[4][8] * mat_B[8][29] +
                  mat_A[4][9] * mat_B[9][29] +
                  mat_A[4][10] * mat_B[10][29] +
                  mat_A[4][11] * mat_B[11][29] +
                  mat_A[4][12] * mat_B[12][29] +
                  mat_A[4][13] * mat_B[13][29] +
                  mat_A[4][14] * mat_B[14][29] +
                  mat_A[4][15] * mat_B[15][29] +
                  mat_A[4][16] * mat_B[16][29] +
                  mat_A[4][17] * mat_B[17][29] +
                  mat_A[4][18] * mat_B[18][29] +
                  mat_A[4][19] * mat_B[19][29] +
                  mat_A[4][20] * mat_B[20][29] +
                  mat_A[4][21] * mat_B[21][29] +
                  mat_A[4][22] * mat_B[22][29] +
                  mat_A[4][23] * mat_B[23][29] +
                  mat_A[4][24] * mat_B[24][29] +
                  mat_A[4][25] * mat_B[25][29] +
                  mat_A[4][26] * mat_B[26][29] +
                  mat_A[4][27] * mat_B[27][29] +
                  mat_A[4][28] * mat_B[28][29] +
                  mat_A[4][29] * mat_B[29][29] +
                  mat_A[4][30] * mat_B[30][29] +
                  mat_A[4][31] * mat_B[31][29];
    mat_C[4][30] <= 
                  mat_A[4][0] * mat_B[0][30] +
                  mat_A[4][1] * mat_B[1][30] +
                  mat_A[4][2] * mat_B[2][30] +
                  mat_A[4][3] * mat_B[3][30] +
                  mat_A[4][4] * mat_B[4][30] +
                  mat_A[4][5] * mat_B[5][30] +
                  mat_A[4][6] * mat_B[6][30] +
                  mat_A[4][7] * mat_B[7][30] +
                  mat_A[4][8] * mat_B[8][30] +
                  mat_A[4][9] * mat_B[9][30] +
                  mat_A[4][10] * mat_B[10][30] +
                  mat_A[4][11] * mat_B[11][30] +
                  mat_A[4][12] * mat_B[12][30] +
                  mat_A[4][13] * mat_B[13][30] +
                  mat_A[4][14] * mat_B[14][30] +
                  mat_A[4][15] * mat_B[15][30] +
                  mat_A[4][16] * mat_B[16][30] +
                  mat_A[4][17] * mat_B[17][30] +
                  mat_A[4][18] * mat_B[18][30] +
                  mat_A[4][19] * mat_B[19][30] +
                  mat_A[4][20] * mat_B[20][30] +
                  mat_A[4][21] * mat_B[21][30] +
                  mat_A[4][22] * mat_B[22][30] +
                  mat_A[4][23] * mat_B[23][30] +
                  mat_A[4][24] * mat_B[24][30] +
                  mat_A[4][25] * mat_B[25][30] +
                  mat_A[4][26] * mat_B[26][30] +
                  mat_A[4][27] * mat_B[27][30] +
                  mat_A[4][28] * mat_B[28][30] +
                  mat_A[4][29] * mat_B[29][30] +
                  mat_A[4][30] * mat_B[30][30] +
                  mat_A[4][31] * mat_B[31][30];
    mat_C[4][31] <= 
                  mat_A[4][0] * mat_B[0][31] +
                  mat_A[4][1] * mat_B[1][31] +
                  mat_A[4][2] * mat_B[2][31] +
                  mat_A[4][3] * mat_B[3][31] +
                  mat_A[4][4] * mat_B[4][31] +
                  mat_A[4][5] * mat_B[5][31] +
                  mat_A[4][6] * mat_B[6][31] +
                  mat_A[4][7] * mat_B[7][31] +
                  mat_A[4][8] * mat_B[8][31] +
                  mat_A[4][9] * mat_B[9][31] +
                  mat_A[4][10] * mat_B[10][31] +
                  mat_A[4][11] * mat_B[11][31] +
                  mat_A[4][12] * mat_B[12][31] +
                  mat_A[4][13] * mat_B[13][31] +
                  mat_A[4][14] * mat_B[14][31] +
                  mat_A[4][15] * mat_B[15][31] +
                  mat_A[4][16] * mat_B[16][31] +
                  mat_A[4][17] * mat_B[17][31] +
                  mat_A[4][18] * mat_B[18][31] +
                  mat_A[4][19] * mat_B[19][31] +
                  mat_A[4][20] * mat_B[20][31] +
                  mat_A[4][21] * mat_B[21][31] +
                  mat_A[4][22] * mat_B[22][31] +
                  mat_A[4][23] * mat_B[23][31] +
                  mat_A[4][24] * mat_B[24][31] +
                  mat_A[4][25] * mat_B[25][31] +
                  mat_A[4][26] * mat_B[26][31] +
                  mat_A[4][27] * mat_B[27][31] +
                  mat_A[4][28] * mat_B[28][31] +
                  mat_A[4][29] * mat_B[29][31] +
                  mat_A[4][30] * mat_B[30][31] +
                  mat_A[4][31] * mat_B[31][31];
    mat_C[5][0] <= 
                  mat_A[5][0] * mat_B[0][0] +
                  mat_A[5][1] * mat_B[1][0] +
                  mat_A[5][2] * mat_B[2][0] +
                  mat_A[5][3] * mat_B[3][0] +
                  mat_A[5][4] * mat_B[4][0] +
                  mat_A[5][5] * mat_B[5][0] +
                  mat_A[5][6] * mat_B[6][0] +
                  mat_A[5][7] * mat_B[7][0] +
                  mat_A[5][8] * mat_B[8][0] +
                  mat_A[5][9] * mat_B[9][0] +
                  mat_A[5][10] * mat_B[10][0] +
                  mat_A[5][11] * mat_B[11][0] +
                  mat_A[5][12] * mat_B[12][0] +
                  mat_A[5][13] * mat_B[13][0] +
                  mat_A[5][14] * mat_B[14][0] +
                  mat_A[5][15] * mat_B[15][0] +
                  mat_A[5][16] * mat_B[16][0] +
                  mat_A[5][17] * mat_B[17][0] +
                  mat_A[5][18] * mat_B[18][0] +
                  mat_A[5][19] * mat_B[19][0] +
                  mat_A[5][20] * mat_B[20][0] +
                  mat_A[5][21] * mat_B[21][0] +
                  mat_A[5][22] * mat_B[22][0] +
                  mat_A[5][23] * mat_B[23][0] +
                  mat_A[5][24] * mat_B[24][0] +
                  mat_A[5][25] * mat_B[25][0] +
                  mat_A[5][26] * mat_B[26][0] +
                  mat_A[5][27] * mat_B[27][0] +
                  mat_A[5][28] * mat_B[28][0] +
                  mat_A[5][29] * mat_B[29][0] +
                  mat_A[5][30] * mat_B[30][0] +
                  mat_A[5][31] * mat_B[31][0];
    mat_C[5][1] <= 
                  mat_A[5][0] * mat_B[0][1] +
                  mat_A[5][1] * mat_B[1][1] +
                  mat_A[5][2] * mat_B[2][1] +
                  mat_A[5][3] * mat_B[3][1] +
                  mat_A[5][4] * mat_B[4][1] +
                  mat_A[5][5] * mat_B[5][1] +
                  mat_A[5][6] * mat_B[6][1] +
                  mat_A[5][7] * mat_B[7][1] +
                  mat_A[5][8] * mat_B[8][1] +
                  mat_A[5][9] * mat_B[9][1] +
                  mat_A[5][10] * mat_B[10][1] +
                  mat_A[5][11] * mat_B[11][1] +
                  mat_A[5][12] * mat_B[12][1] +
                  mat_A[5][13] * mat_B[13][1] +
                  mat_A[5][14] * mat_B[14][1] +
                  mat_A[5][15] * mat_B[15][1] +
                  mat_A[5][16] * mat_B[16][1] +
                  mat_A[5][17] * mat_B[17][1] +
                  mat_A[5][18] * mat_B[18][1] +
                  mat_A[5][19] * mat_B[19][1] +
                  mat_A[5][20] * mat_B[20][1] +
                  mat_A[5][21] * mat_B[21][1] +
                  mat_A[5][22] * mat_B[22][1] +
                  mat_A[5][23] * mat_B[23][1] +
                  mat_A[5][24] * mat_B[24][1] +
                  mat_A[5][25] * mat_B[25][1] +
                  mat_A[5][26] * mat_B[26][1] +
                  mat_A[5][27] * mat_B[27][1] +
                  mat_A[5][28] * mat_B[28][1] +
                  mat_A[5][29] * mat_B[29][1] +
                  mat_A[5][30] * mat_B[30][1] +
                  mat_A[5][31] * mat_B[31][1];
    mat_C[5][2] <= 
                  mat_A[5][0] * mat_B[0][2] +
                  mat_A[5][1] * mat_B[1][2] +
                  mat_A[5][2] * mat_B[2][2] +
                  mat_A[5][3] * mat_B[3][2] +
                  mat_A[5][4] * mat_B[4][2] +
                  mat_A[5][5] * mat_B[5][2] +
                  mat_A[5][6] * mat_B[6][2] +
                  mat_A[5][7] * mat_B[7][2] +
                  mat_A[5][8] * mat_B[8][2] +
                  mat_A[5][9] * mat_B[9][2] +
                  mat_A[5][10] * mat_B[10][2] +
                  mat_A[5][11] * mat_B[11][2] +
                  mat_A[5][12] * mat_B[12][2] +
                  mat_A[5][13] * mat_B[13][2] +
                  mat_A[5][14] * mat_B[14][2] +
                  mat_A[5][15] * mat_B[15][2] +
                  mat_A[5][16] * mat_B[16][2] +
                  mat_A[5][17] * mat_B[17][2] +
                  mat_A[5][18] * mat_B[18][2] +
                  mat_A[5][19] * mat_B[19][2] +
                  mat_A[5][20] * mat_B[20][2] +
                  mat_A[5][21] * mat_B[21][2] +
                  mat_A[5][22] * mat_B[22][2] +
                  mat_A[5][23] * mat_B[23][2] +
                  mat_A[5][24] * mat_B[24][2] +
                  mat_A[5][25] * mat_B[25][2] +
                  mat_A[5][26] * mat_B[26][2] +
                  mat_A[5][27] * mat_B[27][2] +
                  mat_A[5][28] * mat_B[28][2] +
                  mat_A[5][29] * mat_B[29][2] +
                  mat_A[5][30] * mat_B[30][2] +
                  mat_A[5][31] * mat_B[31][2];
    mat_C[5][3] <= 
                  mat_A[5][0] * mat_B[0][3] +
                  mat_A[5][1] * mat_B[1][3] +
                  mat_A[5][2] * mat_B[2][3] +
                  mat_A[5][3] * mat_B[3][3] +
                  mat_A[5][4] * mat_B[4][3] +
                  mat_A[5][5] * mat_B[5][3] +
                  mat_A[5][6] * mat_B[6][3] +
                  mat_A[5][7] * mat_B[7][3] +
                  mat_A[5][8] * mat_B[8][3] +
                  mat_A[5][9] * mat_B[9][3] +
                  mat_A[5][10] * mat_B[10][3] +
                  mat_A[5][11] * mat_B[11][3] +
                  mat_A[5][12] * mat_B[12][3] +
                  mat_A[5][13] * mat_B[13][3] +
                  mat_A[5][14] * mat_B[14][3] +
                  mat_A[5][15] * mat_B[15][3] +
                  mat_A[5][16] * mat_B[16][3] +
                  mat_A[5][17] * mat_B[17][3] +
                  mat_A[5][18] * mat_B[18][3] +
                  mat_A[5][19] * mat_B[19][3] +
                  mat_A[5][20] * mat_B[20][3] +
                  mat_A[5][21] * mat_B[21][3] +
                  mat_A[5][22] * mat_B[22][3] +
                  mat_A[5][23] * mat_B[23][3] +
                  mat_A[5][24] * mat_B[24][3] +
                  mat_A[5][25] * mat_B[25][3] +
                  mat_A[5][26] * mat_B[26][3] +
                  mat_A[5][27] * mat_B[27][3] +
                  mat_A[5][28] * mat_B[28][3] +
                  mat_A[5][29] * mat_B[29][3] +
                  mat_A[5][30] * mat_B[30][3] +
                  mat_A[5][31] * mat_B[31][3];
    mat_C[5][4] <= 
                  mat_A[5][0] * mat_B[0][4] +
                  mat_A[5][1] * mat_B[1][4] +
                  mat_A[5][2] * mat_B[2][4] +
                  mat_A[5][3] * mat_B[3][4] +
                  mat_A[5][4] * mat_B[4][4] +
                  mat_A[5][5] * mat_B[5][4] +
                  mat_A[5][6] * mat_B[6][4] +
                  mat_A[5][7] * mat_B[7][4] +
                  mat_A[5][8] * mat_B[8][4] +
                  mat_A[5][9] * mat_B[9][4] +
                  mat_A[5][10] * mat_B[10][4] +
                  mat_A[5][11] * mat_B[11][4] +
                  mat_A[5][12] * mat_B[12][4] +
                  mat_A[5][13] * mat_B[13][4] +
                  mat_A[5][14] * mat_B[14][4] +
                  mat_A[5][15] * mat_B[15][4] +
                  mat_A[5][16] * mat_B[16][4] +
                  mat_A[5][17] * mat_B[17][4] +
                  mat_A[5][18] * mat_B[18][4] +
                  mat_A[5][19] * mat_B[19][4] +
                  mat_A[5][20] * mat_B[20][4] +
                  mat_A[5][21] * mat_B[21][4] +
                  mat_A[5][22] * mat_B[22][4] +
                  mat_A[5][23] * mat_B[23][4] +
                  mat_A[5][24] * mat_B[24][4] +
                  mat_A[5][25] * mat_B[25][4] +
                  mat_A[5][26] * mat_B[26][4] +
                  mat_A[5][27] * mat_B[27][4] +
                  mat_A[5][28] * mat_B[28][4] +
                  mat_A[5][29] * mat_B[29][4] +
                  mat_A[5][30] * mat_B[30][4] +
                  mat_A[5][31] * mat_B[31][4];
    mat_C[5][5] <= 
                  mat_A[5][0] * mat_B[0][5] +
                  mat_A[5][1] * mat_B[1][5] +
                  mat_A[5][2] * mat_B[2][5] +
                  mat_A[5][3] * mat_B[3][5] +
                  mat_A[5][4] * mat_B[4][5] +
                  mat_A[5][5] * mat_B[5][5] +
                  mat_A[5][6] * mat_B[6][5] +
                  mat_A[5][7] * mat_B[7][5] +
                  mat_A[5][8] * mat_B[8][5] +
                  mat_A[5][9] * mat_B[9][5] +
                  mat_A[5][10] * mat_B[10][5] +
                  mat_A[5][11] * mat_B[11][5] +
                  mat_A[5][12] * mat_B[12][5] +
                  mat_A[5][13] * mat_B[13][5] +
                  mat_A[5][14] * mat_B[14][5] +
                  mat_A[5][15] * mat_B[15][5] +
                  mat_A[5][16] * mat_B[16][5] +
                  mat_A[5][17] * mat_B[17][5] +
                  mat_A[5][18] * mat_B[18][5] +
                  mat_A[5][19] * mat_B[19][5] +
                  mat_A[5][20] * mat_B[20][5] +
                  mat_A[5][21] * mat_B[21][5] +
                  mat_A[5][22] * mat_B[22][5] +
                  mat_A[5][23] * mat_B[23][5] +
                  mat_A[5][24] * mat_B[24][5] +
                  mat_A[5][25] * mat_B[25][5] +
                  mat_A[5][26] * mat_B[26][5] +
                  mat_A[5][27] * mat_B[27][5] +
                  mat_A[5][28] * mat_B[28][5] +
                  mat_A[5][29] * mat_B[29][5] +
                  mat_A[5][30] * mat_B[30][5] +
                  mat_A[5][31] * mat_B[31][5];
    mat_C[5][6] <= 
                  mat_A[5][0] * mat_B[0][6] +
                  mat_A[5][1] * mat_B[1][6] +
                  mat_A[5][2] * mat_B[2][6] +
                  mat_A[5][3] * mat_B[3][6] +
                  mat_A[5][4] * mat_B[4][6] +
                  mat_A[5][5] * mat_B[5][6] +
                  mat_A[5][6] * mat_B[6][6] +
                  mat_A[5][7] * mat_B[7][6] +
                  mat_A[5][8] * mat_B[8][6] +
                  mat_A[5][9] * mat_B[9][6] +
                  mat_A[5][10] * mat_B[10][6] +
                  mat_A[5][11] * mat_B[11][6] +
                  mat_A[5][12] * mat_B[12][6] +
                  mat_A[5][13] * mat_B[13][6] +
                  mat_A[5][14] * mat_B[14][6] +
                  mat_A[5][15] * mat_B[15][6] +
                  mat_A[5][16] * mat_B[16][6] +
                  mat_A[5][17] * mat_B[17][6] +
                  mat_A[5][18] * mat_B[18][6] +
                  mat_A[5][19] * mat_B[19][6] +
                  mat_A[5][20] * mat_B[20][6] +
                  mat_A[5][21] * mat_B[21][6] +
                  mat_A[5][22] * mat_B[22][6] +
                  mat_A[5][23] * mat_B[23][6] +
                  mat_A[5][24] * mat_B[24][6] +
                  mat_A[5][25] * mat_B[25][6] +
                  mat_A[5][26] * mat_B[26][6] +
                  mat_A[5][27] * mat_B[27][6] +
                  mat_A[5][28] * mat_B[28][6] +
                  mat_A[5][29] * mat_B[29][6] +
                  mat_A[5][30] * mat_B[30][6] +
                  mat_A[5][31] * mat_B[31][6];
    mat_C[5][7] <= 
                  mat_A[5][0] * mat_B[0][7] +
                  mat_A[5][1] * mat_B[1][7] +
                  mat_A[5][2] * mat_B[2][7] +
                  mat_A[5][3] * mat_B[3][7] +
                  mat_A[5][4] * mat_B[4][7] +
                  mat_A[5][5] * mat_B[5][7] +
                  mat_A[5][6] * mat_B[6][7] +
                  mat_A[5][7] * mat_B[7][7] +
                  mat_A[5][8] * mat_B[8][7] +
                  mat_A[5][9] * mat_B[9][7] +
                  mat_A[5][10] * mat_B[10][7] +
                  mat_A[5][11] * mat_B[11][7] +
                  mat_A[5][12] * mat_B[12][7] +
                  mat_A[5][13] * mat_B[13][7] +
                  mat_A[5][14] * mat_B[14][7] +
                  mat_A[5][15] * mat_B[15][7] +
                  mat_A[5][16] * mat_B[16][7] +
                  mat_A[5][17] * mat_B[17][7] +
                  mat_A[5][18] * mat_B[18][7] +
                  mat_A[5][19] * mat_B[19][7] +
                  mat_A[5][20] * mat_B[20][7] +
                  mat_A[5][21] * mat_B[21][7] +
                  mat_A[5][22] * mat_B[22][7] +
                  mat_A[5][23] * mat_B[23][7] +
                  mat_A[5][24] * mat_B[24][7] +
                  mat_A[5][25] * mat_B[25][7] +
                  mat_A[5][26] * mat_B[26][7] +
                  mat_A[5][27] * mat_B[27][7] +
                  mat_A[5][28] * mat_B[28][7] +
                  mat_A[5][29] * mat_B[29][7] +
                  mat_A[5][30] * mat_B[30][7] +
                  mat_A[5][31] * mat_B[31][7];
    mat_C[5][8] <= 
                  mat_A[5][0] * mat_B[0][8] +
                  mat_A[5][1] * mat_B[1][8] +
                  mat_A[5][2] * mat_B[2][8] +
                  mat_A[5][3] * mat_B[3][8] +
                  mat_A[5][4] * mat_B[4][8] +
                  mat_A[5][5] * mat_B[5][8] +
                  mat_A[5][6] * mat_B[6][8] +
                  mat_A[5][7] * mat_B[7][8] +
                  mat_A[5][8] * mat_B[8][8] +
                  mat_A[5][9] * mat_B[9][8] +
                  mat_A[5][10] * mat_B[10][8] +
                  mat_A[5][11] * mat_B[11][8] +
                  mat_A[5][12] * mat_B[12][8] +
                  mat_A[5][13] * mat_B[13][8] +
                  mat_A[5][14] * mat_B[14][8] +
                  mat_A[5][15] * mat_B[15][8] +
                  mat_A[5][16] * mat_B[16][8] +
                  mat_A[5][17] * mat_B[17][8] +
                  mat_A[5][18] * mat_B[18][8] +
                  mat_A[5][19] * mat_B[19][8] +
                  mat_A[5][20] * mat_B[20][8] +
                  mat_A[5][21] * mat_B[21][8] +
                  mat_A[5][22] * mat_B[22][8] +
                  mat_A[5][23] * mat_B[23][8] +
                  mat_A[5][24] * mat_B[24][8] +
                  mat_A[5][25] * mat_B[25][8] +
                  mat_A[5][26] * mat_B[26][8] +
                  mat_A[5][27] * mat_B[27][8] +
                  mat_A[5][28] * mat_B[28][8] +
                  mat_A[5][29] * mat_B[29][8] +
                  mat_A[5][30] * mat_B[30][8] +
                  mat_A[5][31] * mat_B[31][8];
    mat_C[5][9] <= 
                  mat_A[5][0] * mat_B[0][9] +
                  mat_A[5][1] * mat_B[1][9] +
                  mat_A[5][2] * mat_B[2][9] +
                  mat_A[5][3] * mat_B[3][9] +
                  mat_A[5][4] * mat_B[4][9] +
                  mat_A[5][5] * mat_B[5][9] +
                  mat_A[5][6] * mat_B[6][9] +
                  mat_A[5][7] * mat_B[7][9] +
                  mat_A[5][8] * mat_B[8][9] +
                  mat_A[5][9] * mat_B[9][9] +
                  mat_A[5][10] * mat_B[10][9] +
                  mat_A[5][11] * mat_B[11][9] +
                  mat_A[5][12] * mat_B[12][9] +
                  mat_A[5][13] * mat_B[13][9] +
                  mat_A[5][14] * mat_B[14][9] +
                  mat_A[5][15] * mat_B[15][9] +
                  mat_A[5][16] * mat_B[16][9] +
                  mat_A[5][17] * mat_B[17][9] +
                  mat_A[5][18] * mat_B[18][9] +
                  mat_A[5][19] * mat_B[19][9] +
                  mat_A[5][20] * mat_B[20][9] +
                  mat_A[5][21] * mat_B[21][9] +
                  mat_A[5][22] * mat_B[22][9] +
                  mat_A[5][23] * mat_B[23][9] +
                  mat_A[5][24] * mat_B[24][9] +
                  mat_A[5][25] * mat_B[25][9] +
                  mat_A[5][26] * mat_B[26][9] +
                  mat_A[5][27] * mat_B[27][9] +
                  mat_A[5][28] * mat_B[28][9] +
                  mat_A[5][29] * mat_B[29][9] +
                  mat_A[5][30] * mat_B[30][9] +
                  mat_A[5][31] * mat_B[31][9];
    mat_C[5][10] <= 
                  mat_A[5][0] * mat_B[0][10] +
                  mat_A[5][1] * mat_B[1][10] +
                  mat_A[5][2] * mat_B[2][10] +
                  mat_A[5][3] * mat_B[3][10] +
                  mat_A[5][4] * mat_B[4][10] +
                  mat_A[5][5] * mat_B[5][10] +
                  mat_A[5][6] * mat_B[6][10] +
                  mat_A[5][7] * mat_B[7][10] +
                  mat_A[5][8] * mat_B[8][10] +
                  mat_A[5][9] * mat_B[9][10] +
                  mat_A[5][10] * mat_B[10][10] +
                  mat_A[5][11] * mat_B[11][10] +
                  mat_A[5][12] * mat_B[12][10] +
                  mat_A[5][13] * mat_B[13][10] +
                  mat_A[5][14] * mat_B[14][10] +
                  mat_A[5][15] * mat_B[15][10] +
                  mat_A[5][16] * mat_B[16][10] +
                  mat_A[5][17] * mat_B[17][10] +
                  mat_A[5][18] * mat_B[18][10] +
                  mat_A[5][19] * mat_B[19][10] +
                  mat_A[5][20] * mat_B[20][10] +
                  mat_A[5][21] * mat_B[21][10] +
                  mat_A[5][22] * mat_B[22][10] +
                  mat_A[5][23] * mat_B[23][10] +
                  mat_A[5][24] * mat_B[24][10] +
                  mat_A[5][25] * mat_B[25][10] +
                  mat_A[5][26] * mat_B[26][10] +
                  mat_A[5][27] * mat_B[27][10] +
                  mat_A[5][28] * mat_B[28][10] +
                  mat_A[5][29] * mat_B[29][10] +
                  mat_A[5][30] * mat_B[30][10] +
                  mat_A[5][31] * mat_B[31][10];
    mat_C[5][11] <= 
                  mat_A[5][0] * mat_B[0][11] +
                  mat_A[5][1] * mat_B[1][11] +
                  mat_A[5][2] * mat_B[2][11] +
                  mat_A[5][3] * mat_B[3][11] +
                  mat_A[5][4] * mat_B[4][11] +
                  mat_A[5][5] * mat_B[5][11] +
                  mat_A[5][6] * mat_B[6][11] +
                  mat_A[5][7] * mat_B[7][11] +
                  mat_A[5][8] * mat_B[8][11] +
                  mat_A[5][9] * mat_B[9][11] +
                  mat_A[5][10] * mat_B[10][11] +
                  mat_A[5][11] * mat_B[11][11] +
                  mat_A[5][12] * mat_B[12][11] +
                  mat_A[5][13] * mat_B[13][11] +
                  mat_A[5][14] * mat_B[14][11] +
                  mat_A[5][15] * mat_B[15][11] +
                  mat_A[5][16] * mat_B[16][11] +
                  mat_A[5][17] * mat_B[17][11] +
                  mat_A[5][18] * mat_B[18][11] +
                  mat_A[5][19] * mat_B[19][11] +
                  mat_A[5][20] * mat_B[20][11] +
                  mat_A[5][21] * mat_B[21][11] +
                  mat_A[5][22] * mat_B[22][11] +
                  mat_A[5][23] * mat_B[23][11] +
                  mat_A[5][24] * mat_B[24][11] +
                  mat_A[5][25] * mat_B[25][11] +
                  mat_A[5][26] * mat_B[26][11] +
                  mat_A[5][27] * mat_B[27][11] +
                  mat_A[5][28] * mat_B[28][11] +
                  mat_A[5][29] * mat_B[29][11] +
                  mat_A[5][30] * mat_B[30][11] +
                  mat_A[5][31] * mat_B[31][11];
    mat_C[5][12] <= 
                  mat_A[5][0] * mat_B[0][12] +
                  mat_A[5][1] * mat_B[1][12] +
                  mat_A[5][2] * mat_B[2][12] +
                  mat_A[5][3] * mat_B[3][12] +
                  mat_A[5][4] * mat_B[4][12] +
                  mat_A[5][5] * mat_B[5][12] +
                  mat_A[5][6] * mat_B[6][12] +
                  mat_A[5][7] * mat_B[7][12] +
                  mat_A[5][8] * mat_B[8][12] +
                  mat_A[5][9] * mat_B[9][12] +
                  mat_A[5][10] * mat_B[10][12] +
                  mat_A[5][11] * mat_B[11][12] +
                  mat_A[5][12] * mat_B[12][12] +
                  mat_A[5][13] * mat_B[13][12] +
                  mat_A[5][14] * mat_B[14][12] +
                  mat_A[5][15] * mat_B[15][12] +
                  mat_A[5][16] * mat_B[16][12] +
                  mat_A[5][17] * mat_B[17][12] +
                  mat_A[5][18] * mat_B[18][12] +
                  mat_A[5][19] * mat_B[19][12] +
                  mat_A[5][20] * mat_B[20][12] +
                  mat_A[5][21] * mat_B[21][12] +
                  mat_A[5][22] * mat_B[22][12] +
                  mat_A[5][23] * mat_B[23][12] +
                  mat_A[5][24] * mat_B[24][12] +
                  mat_A[5][25] * mat_B[25][12] +
                  mat_A[5][26] * mat_B[26][12] +
                  mat_A[5][27] * mat_B[27][12] +
                  mat_A[5][28] * mat_B[28][12] +
                  mat_A[5][29] * mat_B[29][12] +
                  mat_A[5][30] * mat_B[30][12] +
                  mat_A[5][31] * mat_B[31][12];
    mat_C[5][13] <= 
                  mat_A[5][0] * mat_B[0][13] +
                  mat_A[5][1] * mat_B[1][13] +
                  mat_A[5][2] * mat_B[2][13] +
                  mat_A[5][3] * mat_B[3][13] +
                  mat_A[5][4] * mat_B[4][13] +
                  mat_A[5][5] * mat_B[5][13] +
                  mat_A[5][6] * mat_B[6][13] +
                  mat_A[5][7] * mat_B[7][13] +
                  mat_A[5][8] * mat_B[8][13] +
                  mat_A[5][9] * mat_B[9][13] +
                  mat_A[5][10] * mat_B[10][13] +
                  mat_A[5][11] * mat_B[11][13] +
                  mat_A[5][12] * mat_B[12][13] +
                  mat_A[5][13] * mat_B[13][13] +
                  mat_A[5][14] * mat_B[14][13] +
                  mat_A[5][15] * mat_B[15][13] +
                  mat_A[5][16] * mat_B[16][13] +
                  mat_A[5][17] * mat_B[17][13] +
                  mat_A[5][18] * mat_B[18][13] +
                  mat_A[5][19] * mat_B[19][13] +
                  mat_A[5][20] * mat_B[20][13] +
                  mat_A[5][21] * mat_B[21][13] +
                  mat_A[5][22] * mat_B[22][13] +
                  mat_A[5][23] * mat_B[23][13] +
                  mat_A[5][24] * mat_B[24][13] +
                  mat_A[5][25] * mat_B[25][13] +
                  mat_A[5][26] * mat_B[26][13] +
                  mat_A[5][27] * mat_B[27][13] +
                  mat_A[5][28] * mat_B[28][13] +
                  mat_A[5][29] * mat_B[29][13] +
                  mat_A[5][30] * mat_B[30][13] +
                  mat_A[5][31] * mat_B[31][13];
    mat_C[5][14] <= 
                  mat_A[5][0] * mat_B[0][14] +
                  mat_A[5][1] * mat_B[1][14] +
                  mat_A[5][2] * mat_B[2][14] +
                  mat_A[5][3] * mat_B[3][14] +
                  mat_A[5][4] * mat_B[4][14] +
                  mat_A[5][5] * mat_B[5][14] +
                  mat_A[5][6] * mat_B[6][14] +
                  mat_A[5][7] * mat_B[7][14] +
                  mat_A[5][8] * mat_B[8][14] +
                  mat_A[5][9] * mat_B[9][14] +
                  mat_A[5][10] * mat_B[10][14] +
                  mat_A[5][11] * mat_B[11][14] +
                  mat_A[5][12] * mat_B[12][14] +
                  mat_A[5][13] * mat_B[13][14] +
                  mat_A[5][14] * mat_B[14][14] +
                  mat_A[5][15] * mat_B[15][14] +
                  mat_A[5][16] * mat_B[16][14] +
                  mat_A[5][17] * mat_B[17][14] +
                  mat_A[5][18] * mat_B[18][14] +
                  mat_A[5][19] * mat_B[19][14] +
                  mat_A[5][20] * mat_B[20][14] +
                  mat_A[5][21] * mat_B[21][14] +
                  mat_A[5][22] * mat_B[22][14] +
                  mat_A[5][23] * mat_B[23][14] +
                  mat_A[5][24] * mat_B[24][14] +
                  mat_A[5][25] * mat_B[25][14] +
                  mat_A[5][26] * mat_B[26][14] +
                  mat_A[5][27] * mat_B[27][14] +
                  mat_A[5][28] * mat_B[28][14] +
                  mat_A[5][29] * mat_B[29][14] +
                  mat_A[5][30] * mat_B[30][14] +
                  mat_A[5][31] * mat_B[31][14];
    mat_C[5][15] <= 
                  mat_A[5][0] * mat_B[0][15] +
                  mat_A[5][1] * mat_B[1][15] +
                  mat_A[5][2] * mat_B[2][15] +
                  mat_A[5][3] * mat_B[3][15] +
                  mat_A[5][4] * mat_B[4][15] +
                  mat_A[5][5] * mat_B[5][15] +
                  mat_A[5][6] * mat_B[6][15] +
                  mat_A[5][7] * mat_B[7][15] +
                  mat_A[5][8] * mat_B[8][15] +
                  mat_A[5][9] * mat_B[9][15] +
                  mat_A[5][10] * mat_B[10][15] +
                  mat_A[5][11] * mat_B[11][15] +
                  mat_A[5][12] * mat_B[12][15] +
                  mat_A[5][13] * mat_B[13][15] +
                  mat_A[5][14] * mat_B[14][15] +
                  mat_A[5][15] * mat_B[15][15] +
                  mat_A[5][16] * mat_B[16][15] +
                  mat_A[5][17] * mat_B[17][15] +
                  mat_A[5][18] * mat_B[18][15] +
                  mat_A[5][19] * mat_B[19][15] +
                  mat_A[5][20] * mat_B[20][15] +
                  mat_A[5][21] * mat_B[21][15] +
                  mat_A[5][22] * mat_B[22][15] +
                  mat_A[5][23] * mat_B[23][15] +
                  mat_A[5][24] * mat_B[24][15] +
                  mat_A[5][25] * mat_B[25][15] +
                  mat_A[5][26] * mat_B[26][15] +
                  mat_A[5][27] * mat_B[27][15] +
                  mat_A[5][28] * mat_B[28][15] +
                  mat_A[5][29] * mat_B[29][15] +
                  mat_A[5][30] * mat_B[30][15] +
                  mat_A[5][31] * mat_B[31][15];
    mat_C[5][16] <= 
                  mat_A[5][0] * mat_B[0][16] +
                  mat_A[5][1] * mat_B[1][16] +
                  mat_A[5][2] * mat_B[2][16] +
                  mat_A[5][3] * mat_B[3][16] +
                  mat_A[5][4] * mat_B[4][16] +
                  mat_A[5][5] * mat_B[5][16] +
                  mat_A[5][6] * mat_B[6][16] +
                  mat_A[5][7] * mat_B[7][16] +
                  mat_A[5][8] * mat_B[8][16] +
                  mat_A[5][9] * mat_B[9][16] +
                  mat_A[5][10] * mat_B[10][16] +
                  mat_A[5][11] * mat_B[11][16] +
                  mat_A[5][12] * mat_B[12][16] +
                  mat_A[5][13] * mat_B[13][16] +
                  mat_A[5][14] * mat_B[14][16] +
                  mat_A[5][15] * mat_B[15][16] +
                  mat_A[5][16] * mat_B[16][16] +
                  mat_A[5][17] * mat_B[17][16] +
                  mat_A[5][18] * mat_B[18][16] +
                  mat_A[5][19] * mat_B[19][16] +
                  mat_A[5][20] * mat_B[20][16] +
                  mat_A[5][21] * mat_B[21][16] +
                  mat_A[5][22] * mat_B[22][16] +
                  mat_A[5][23] * mat_B[23][16] +
                  mat_A[5][24] * mat_B[24][16] +
                  mat_A[5][25] * mat_B[25][16] +
                  mat_A[5][26] * mat_B[26][16] +
                  mat_A[5][27] * mat_B[27][16] +
                  mat_A[5][28] * mat_B[28][16] +
                  mat_A[5][29] * mat_B[29][16] +
                  mat_A[5][30] * mat_B[30][16] +
                  mat_A[5][31] * mat_B[31][16];
    mat_C[5][17] <= 
                  mat_A[5][0] * mat_B[0][17] +
                  mat_A[5][1] * mat_B[1][17] +
                  mat_A[5][2] * mat_B[2][17] +
                  mat_A[5][3] * mat_B[3][17] +
                  mat_A[5][4] * mat_B[4][17] +
                  mat_A[5][5] * mat_B[5][17] +
                  mat_A[5][6] * mat_B[6][17] +
                  mat_A[5][7] * mat_B[7][17] +
                  mat_A[5][8] * mat_B[8][17] +
                  mat_A[5][9] * mat_B[9][17] +
                  mat_A[5][10] * mat_B[10][17] +
                  mat_A[5][11] * mat_B[11][17] +
                  mat_A[5][12] * mat_B[12][17] +
                  mat_A[5][13] * mat_B[13][17] +
                  mat_A[5][14] * mat_B[14][17] +
                  mat_A[5][15] * mat_B[15][17] +
                  mat_A[5][16] * mat_B[16][17] +
                  mat_A[5][17] * mat_B[17][17] +
                  mat_A[5][18] * mat_B[18][17] +
                  mat_A[5][19] * mat_B[19][17] +
                  mat_A[5][20] * mat_B[20][17] +
                  mat_A[5][21] * mat_B[21][17] +
                  mat_A[5][22] * mat_B[22][17] +
                  mat_A[5][23] * mat_B[23][17] +
                  mat_A[5][24] * mat_B[24][17] +
                  mat_A[5][25] * mat_B[25][17] +
                  mat_A[5][26] * mat_B[26][17] +
                  mat_A[5][27] * mat_B[27][17] +
                  mat_A[5][28] * mat_B[28][17] +
                  mat_A[5][29] * mat_B[29][17] +
                  mat_A[5][30] * mat_B[30][17] +
                  mat_A[5][31] * mat_B[31][17];
    mat_C[5][18] <= 
                  mat_A[5][0] * mat_B[0][18] +
                  mat_A[5][1] * mat_B[1][18] +
                  mat_A[5][2] * mat_B[2][18] +
                  mat_A[5][3] * mat_B[3][18] +
                  mat_A[5][4] * mat_B[4][18] +
                  mat_A[5][5] * mat_B[5][18] +
                  mat_A[5][6] * mat_B[6][18] +
                  mat_A[5][7] * mat_B[7][18] +
                  mat_A[5][8] * mat_B[8][18] +
                  mat_A[5][9] * mat_B[9][18] +
                  mat_A[5][10] * mat_B[10][18] +
                  mat_A[5][11] * mat_B[11][18] +
                  mat_A[5][12] * mat_B[12][18] +
                  mat_A[5][13] * mat_B[13][18] +
                  mat_A[5][14] * mat_B[14][18] +
                  mat_A[5][15] * mat_B[15][18] +
                  mat_A[5][16] * mat_B[16][18] +
                  mat_A[5][17] * mat_B[17][18] +
                  mat_A[5][18] * mat_B[18][18] +
                  mat_A[5][19] * mat_B[19][18] +
                  mat_A[5][20] * mat_B[20][18] +
                  mat_A[5][21] * mat_B[21][18] +
                  mat_A[5][22] * mat_B[22][18] +
                  mat_A[5][23] * mat_B[23][18] +
                  mat_A[5][24] * mat_B[24][18] +
                  mat_A[5][25] * mat_B[25][18] +
                  mat_A[5][26] * mat_B[26][18] +
                  mat_A[5][27] * mat_B[27][18] +
                  mat_A[5][28] * mat_B[28][18] +
                  mat_A[5][29] * mat_B[29][18] +
                  mat_A[5][30] * mat_B[30][18] +
                  mat_A[5][31] * mat_B[31][18];
    mat_C[5][19] <= 
                  mat_A[5][0] * mat_B[0][19] +
                  mat_A[5][1] * mat_B[1][19] +
                  mat_A[5][2] * mat_B[2][19] +
                  mat_A[5][3] * mat_B[3][19] +
                  mat_A[5][4] * mat_B[4][19] +
                  mat_A[5][5] * mat_B[5][19] +
                  mat_A[5][6] * mat_B[6][19] +
                  mat_A[5][7] * mat_B[7][19] +
                  mat_A[5][8] * mat_B[8][19] +
                  mat_A[5][9] * mat_B[9][19] +
                  mat_A[5][10] * mat_B[10][19] +
                  mat_A[5][11] * mat_B[11][19] +
                  mat_A[5][12] * mat_B[12][19] +
                  mat_A[5][13] * mat_B[13][19] +
                  mat_A[5][14] * mat_B[14][19] +
                  mat_A[5][15] * mat_B[15][19] +
                  mat_A[5][16] * mat_B[16][19] +
                  mat_A[5][17] * mat_B[17][19] +
                  mat_A[5][18] * mat_B[18][19] +
                  mat_A[5][19] * mat_B[19][19] +
                  mat_A[5][20] * mat_B[20][19] +
                  mat_A[5][21] * mat_B[21][19] +
                  mat_A[5][22] * mat_B[22][19] +
                  mat_A[5][23] * mat_B[23][19] +
                  mat_A[5][24] * mat_B[24][19] +
                  mat_A[5][25] * mat_B[25][19] +
                  mat_A[5][26] * mat_B[26][19] +
                  mat_A[5][27] * mat_B[27][19] +
                  mat_A[5][28] * mat_B[28][19] +
                  mat_A[5][29] * mat_B[29][19] +
                  mat_A[5][30] * mat_B[30][19] +
                  mat_A[5][31] * mat_B[31][19];
    mat_C[5][20] <= 
                  mat_A[5][0] * mat_B[0][20] +
                  mat_A[5][1] * mat_B[1][20] +
                  mat_A[5][2] * mat_B[2][20] +
                  mat_A[5][3] * mat_B[3][20] +
                  mat_A[5][4] * mat_B[4][20] +
                  mat_A[5][5] * mat_B[5][20] +
                  mat_A[5][6] * mat_B[6][20] +
                  mat_A[5][7] * mat_B[7][20] +
                  mat_A[5][8] * mat_B[8][20] +
                  mat_A[5][9] * mat_B[9][20] +
                  mat_A[5][10] * mat_B[10][20] +
                  mat_A[5][11] * mat_B[11][20] +
                  mat_A[5][12] * mat_B[12][20] +
                  mat_A[5][13] * mat_B[13][20] +
                  mat_A[5][14] * mat_B[14][20] +
                  mat_A[5][15] * mat_B[15][20] +
                  mat_A[5][16] * mat_B[16][20] +
                  mat_A[5][17] * mat_B[17][20] +
                  mat_A[5][18] * mat_B[18][20] +
                  mat_A[5][19] * mat_B[19][20] +
                  mat_A[5][20] * mat_B[20][20] +
                  mat_A[5][21] * mat_B[21][20] +
                  mat_A[5][22] * mat_B[22][20] +
                  mat_A[5][23] * mat_B[23][20] +
                  mat_A[5][24] * mat_B[24][20] +
                  mat_A[5][25] * mat_B[25][20] +
                  mat_A[5][26] * mat_B[26][20] +
                  mat_A[5][27] * mat_B[27][20] +
                  mat_A[5][28] * mat_B[28][20] +
                  mat_A[5][29] * mat_B[29][20] +
                  mat_A[5][30] * mat_B[30][20] +
                  mat_A[5][31] * mat_B[31][20];
    mat_C[5][21] <= 
                  mat_A[5][0] * mat_B[0][21] +
                  mat_A[5][1] * mat_B[1][21] +
                  mat_A[5][2] * mat_B[2][21] +
                  mat_A[5][3] * mat_B[3][21] +
                  mat_A[5][4] * mat_B[4][21] +
                  mat_A[5][5] * mat_B[5][21] +
                  mat_A[5][6] * mat_B[6][21] +
                  mat_A[5][7] * mat_B[7][21] +
                  mat_A[5][8] * mat_B[8][21] +
                  mat_A[5][9] * mat_B[9][21] +
                  mat_A[5][10] * mat_B[10][21] +
                  mat_A[5][11] * mat_B[11][21] +
                  mat_A[5][12] * mat_B[12][21] +
                  mat_A[5][13] * mat_B[13][21] +
                  mat_A[5][14] * mat_B[14][21] +
                  mat_A[5][15] * mat_B[15][21] +
                  mat_A[5][16] * mat_B[16][21] +
                  mat_A[5][17] * mat_B[17][21] +
                  mat_A[5][18] * mat_B[18][21] +
                  mat_A[5][19] * mat_B[19][21] +
                  mat_A[5][20] * mat_B[20][21] +
                  mat_A[5][21] * mat_B[21][21] +
                  mat_A[5][22] * mat_B[22][21] +
                  mat_A[5][23] * mat_B[23][21] +
                  mat_A[5][24] * mat_B[24][21] +
                  mat_A[5][25] * mat_B[25][21] +
                  mat_A[5][26] * mat_B[26][21] +
                  mat_A[5][27] * mat_B[27][21] +
                  mat_A[5][28] * mat_B[28][21] +
                  mat_A[5][29] * mat_B[29][21] +
                  mat_A[5][30] * mat_B[30][21] +
                  mat_A[5][31] * mat_B[31][21];
    mat_C[5][22] <= 
                  mat_A[5][0] * mat_B[0][22] +
                  mat_A[5][1] * mat_B[1][22] +
                  mat_A[5][2] * mat_B[2][22] +
                  mat_A[5][3] * mat_B[3][22] +
                  mat_A[5][4] * mat_B[4][22] +
                  mat_A[5][5] * mat_B[5][22] +
                  mat_A[5][6] * mat_B[6][22] +
                  mat_A[5][7] * mat_B[7][22] +
                  mat_A[5][8] * mat_B[8][22] +
                  mat_A[5][9] * mat_B[9][22] +
                  mat_A[5][10] * mat_B[10][22] +
                  mat_A[5][11] * mat_B[11][22] +
                  mat_A[5][12] * mat_B[12][22] +
                  mat_A[5][13] * mat_B[13][22] +
                  mat_A[5][14] * mat_B[14][22] +
                  mat_A[5][15] * mat_B[15][22] +
                  mat_A[5][16] * mat_B[16][22] +
                  mat_A[5][17] * mat_B[17][22] +
                  mat_A[5][18] * mat_B[18][22] +
                  mat_A[5][19] * mat_B[19][22] +
                  mat_A[5][20] * mat_B[20][22] +
                  mat_A[5][21] * mat_B[21][22] +
                  mat_A[5][22] * mat_B[22][22] +
                  mat_A[5][23] * mat_B[23][22] +
                  mat_A[5][24] * mat_B[24][22] +
                  mat_A[5][25] * mat_B[25][22] +
                  mat_A[5][26] * mat_B[26][22] +
                  mat_A[5][27] * mat_B[27][22] +
                  mat_A[5][28] * mat_B[28][22] +
                  mat_A[5][29] * mat_B[29][22] +
                  mat_A[5][30] * mat_B[30][22] +
                  mat_A[5][31] * mat_B[31][22];
    mat_C[5][23] <= 
                  mat_A[5][0] * mat_B[0][23] +
                  mat_A[5][1] * mat_B[1][23] +
                  mat_A[5][2] * mat_B[2][23] +
                  mat_A[5][3] * mat_B[3][23] +
                  mat_A[5][4] * mat_B[4][23] +
                  mat_A[5][5] * mat_B[5][23] +
                  mat_A[5][6] * mat_B[6][23] +
                  mat_A[5][7] * mat_B[7][23] +
                  mat_A[5][8] * mat_B[8][23] +
                  mat_A[5][9] * mat_B[9][23] +
                  mat_A[5][10] * mat_B[10][23] +
                  mat_A[5][11] * mat_B[11][23] +
                  mat_A[5][12] * mat_B[12][23] +
                  mat_A[5][13] * mat_B[13][23] +
                  mat_A[5][14] * mat_B[14][23] +
                  mat_A[5][15] * mat_B[15][23] +
                  mat_A[5][16] * mat_B[16][23] +
                  mat_A[5][17] * mat_B[17][23] +
                  mat_A[5][18] * mat_B[18][23] +
                  mat_A[5][19] * mat_B[19][23] +
                  mat_A[5][20] * mat_B[20][23] +
                  mat_A[5][21] * mat_B[21][23] +
                  mat_A[5][22] * mat_B[22][23] +
                  mat_A[5][23] * mat_B[23][23] +
                  mat_A[5][24] * mat_B[24][23] +
                  mat_A[5][25] * mat_B[25][23] +
                  mat_A[5][26] * mat_B[26][23] +
                  mat_A[5][27] * mat_B[27][23] +
                  mat_A[5][28] * mat_B[28][23] +
                  mat_A[5][29] * mat_B[29][23] +
                  mat_A[5][30] * mat_B[30][23] +
                  mat_A[5][31] * mat_B[31][23];
    mat_C[5][24] <= 
                  mat_A[5][0] * mat_B[0][24] +
                  mat_A[5][1] * mat_B[1][24] +
                  mat_A[5][2] * mat_B[2][24] +
                  mat_A[5][3] * mat_B[3][24] +
                  mat_A[5][4] * mat_B[4][24] +
                  mat_A[5][5] * mat_B[5][24] +
                  mat_A[5][6] * mat_B[6][24] +
                  mat_A[5][7] * mat_B[7][24] +
                  mat_A[5][8] * mat_B[8][24] +
                  mat_A[5][9] * mat_B[9][24] +
                  mat_A[5][10] * mat_B[10][24] +
                  mat_A[5][11] * mat_B[11][24] +
                  mat_A[5][12] * mat_B[12][24] +
                  mat_A[5][13] * mat_B[13][24] +
                  mat_A[5][14] * mat_B[14][24] +
                  mat_A[5][15] * mat_B[15][24] +
                  mat_A[5][16] * mat_B[16][24] +
                  mat_A[5][17] * mat_B[17][24] +
                  mat_A[5][18] * mat_B[18][24] +
                  mat_A[5][19] * mat_B[19][24] +
                  mat_A[5][20] * mat_B[20][24] +
                  mat_A[5][21] * mat_B[21][24] +
                  mat_A[5][22] * mat_B[22][24] +
                  mat_A[5][23] * mat_B[23][24] +
                  mat_A[5][24] * mat_B[24][24] +
                  mat_A[5][25] * mat_B[25][24] +
                  mat_A[5][26] * mat_B[26][24] +
                  mat_A[5][27] * mat_B[27][24] +
                  mat_A[5][28] * mat_B[28][24] +
                  mat_A[5][29] * mat_B[29][24] +
                  mat_A[5][30] * mat_B[30][24] +
                  mat_A[5][31] * mat_B[31][24];
    mat_C[5][25] <= 
                  mat_A[5][0] * mat_B[0][25] +
                  mat_A[5][1] * mat_B[1][25] +
                  mat_A[5][2] * mat_B[2][25] +
                  mat_A[5][3] * mat_B[3][25] +
                  mat_A[5][4] * mat_B[4][25] +
                  mat_A[5][5] * mat_B[5][25] +
                  mat_A[5][6] * mat_B[6][25] +
                  mat_A[5][7] * mat_B[7][25] +
                  mat_A[5][8] * mat_B[8][25] +
                  mat_A[5][9] * mat_B[9][25] +
                  mat_A[5][10] * mat_B[10][25] +
                  mat_A[5][11] * mat_B[11][25] +
                  mat_A[5][12] * mat_B[12][25] +
                  mat_A[5][13] * mat_B[13][25] +
                  mat_A[5][14] * mat_B[14][25] +
                  mat_A[5][15] * mat_B[15][25] +
                  mat_A[5][16] * mat_B[16][25] +
                  mat_A[5][17] * mat_B[17][25] +
                  mat_A[5][18] * mat_B[18][25] +
                  mat_A[5][19] * mat_B[19][25] +
                  mat_A[5][20] * mat_B[20][25] +
                  mat_A[5][21] * mat_B[21][25] +
                  mat_A[5][22] * mat_B[22][25] +
                  mat_A[5][23] * mat_B[23][25] +
                  mat_A[5][24] * mat_B[24][25] +
                  mat_A[5][25] * mat_B[25][25] +
                  mat_A[5][26] * mat_B[26][25] +
                  mat_A[5][27] * mat_B[27][25] +
                  mat_A[5][28] * mat_B[28][25] +
                  mat_A[5][29] * mat_B[29][25] +
                  mat_A[5][30] * mat_B[30][25] +
                  mat_A[5][31] * mat_B[31][25];
    mat_C[5][26] <= 
                  mat_A[5][0] * mat_B[0][26] +
                  mat_A[5][1] * mat_B[1][26] +
                  mat_A[5][2] * mat_B[2][26] +
                  mat_A[5][3] * mat_B[3][26] +
                  mat_A[5][4] * mat_B[4][26] +
                  mat_A[5][5] * mat_B[5][26] +
                  mat_A[5][6] * mat_B[6][26] +
                  mat_A[5][7] * mat_B[7][26] +
                  mat_A[5][8] * mat_B[8][26] +
                  mat_A[5][9] * mat_B[9][26] +
                  mat_A[5][10] * mat_B[10][26] +
                  mat_A[5][11] * mat_B[11][26] +
                  mat_A[5][12] * mat_B[12][26] +
                  mat_A[5][13] * mat_B[13][26] +
                  mat_A[5][14] * mat_B[14][26] +
                  mat_A[5][15] * mat_B[15][26] +
                  mat_A[5][16] * mat_B[16][26] +
                  mat_A[5][17] * mat_B[17][26] +
                  mat_A[5][18] * mat_B[18][26] +
                  mat_A[5][19] * mat_B[19][26] +
                  mat_A[5][20] * mat_B[20][26] +
                  mat_A[5][21] * mat_B[21][26] +
                  mat_A[5][22] * mat_B[22][26] +
                  mat_A[5][23] * mat_B[23][26] +
                  mat_A[5][24] * mat_B[24][26] +
                  mat_A[5][25] * mat_B[25][26] +
                  mat_A[5][26] * mat_B[26][26] +
                  mat_A[5][27] * mat_B[27][26] +
                  mat_A[5][28] * mat_B[28][26] +
                  mat_A[5][29] * mat_B[29][26] +
                  mat_A[5][30] * mat_B[30][26] +
                  mat_A[5][31] * mat_B[31][26];
    mat_C[5][27] <= 
                  mat_A[5][0] * mat_B[0][27] +
                  mat_A[5][1] * mat_B[1][27] +
                  mat_A[5][2] * mat_B[2][27] +
                  mat_A[5][3] * mat_B[3][27] +
                  mat_A[5][4] * mat_B[4][27] +
                  mat_A[5][5] * mat_B[5][27] +
                  mat_A[5][6] * mat_B[6][27] +
                  mat_A[5][7] * mat_B[7][27] +
                  mat_A[5][8] * mat_B[8][27] +
                  mat_A[5][9] * mat_B[9][27] +
                  mat_A[5][10] * mat_B[10][27] +
                  mat_A[5][11] * mat_B[11][27] +
                  mat_A[5][12] * mat_B[12][27] +
                  mat_A[5][13] * mat_B[13][27] +
                  mat_A[5][14] * mat_B[14][27] +
                  mat_A[5][15] * mat_B[15][27] +
                  mat_A[5][16] * mat_B[16][27] +
                  mat_A[5][17] * mat_B[17][27] +
                  mat_A[5][18] * mat_B[18][27] +
                  mat_A[5][19] * mat_B[19][27] +
                  mat_A[5][20] * mat_B[20][27] +
                  mat_A[5][21] * mat_B[21][27] +
                  mat_A[5][22] * mat_B[22][27] +
                  mat_A[5][23] * mat_B[23][27] +
                  mat_A[5][24] * mat_B[24][27] +
                  mat_A[5][25] * mat_B[25][27] +
                  mat_A[5][26] * mat_B[26][27] +
                  mat_A[5][27] * mat_B[27][27] +
                  mat_A[5][28] * mat_B[28][27] +
                  mat_A[5][29] * mat_B[29][27] +
                  mat_A[5][30] * mat_B[30][27] +
                  mat_A[5][31] * mat_B[31][27];
    mat_C[5][28] <= 
                  mat_A[5][0] * mat_B[0][28] +
                  mat_A[5][1] * mat_B[1][28] +
                  mat_A[5][2] * mat_B[2][28] +
                  mat_A[5][3] * mat_B[3][28] +
                  mat_A[5][4] * mat_B[4][28] +
                  mat_A[5][5] * mat_B[5][28] +
                  mat_A[5][6] * mat_B[6][28] +
                  mat_A[5][7] * mat_B[7][28] +
                  mat_A[5][8] * mat_B[8][28] +
                  mat_A[5][9] * mat_B[9][28] +
                  mat_A[5][10] * mat_B[10][28] +
                  mat_A[5][11] * mat_B[11][28] +
                  mat_A[5][12] * mat_B[12][28] +
                  mat_A[5][13] * mat_B[13][28] +
                  mat_A[5][14] * mat_B[14][28] +
                  mat_A[5][15] * mat_B[15][28] +
                  mat_A[5][16] * mat_B[16][28] +
                  mat_A[5][17] * mat_B[17][28] +
                  mat_A[5][18] * mat_B[18][28] +
                  mat_A[5][19] * mat_B[19][28] +
                  mat_A[5][20] * mat_B[20][28] +
                  mat_A[5][21] * mat_B[21][28] +
                  mat_A[5][22] * mat_B[22][28] +
                  mat_A[5][23] * mat_B[23][28] +
                  mat_A[5][24] * mat_B[24][28] +
                  mat_A[5][25] * mat_B[25][28] +
                  mat_A[5][26] * mat_B[26][28] +
                  mat_A[5][27] * mat_B[27][28] +
                  mat_A[5][28] * mat_B[28][28] +
                  mat_A[5][29] * mat_B[29][28] +
                  mat_A[5][30] * mat_B[30][28] +
                  mat_A[5][31] * mat_B[31][28];
    mat_C[5][29] <= 
                  mat_A[5][0] * mat_B[0][29] +
                  mat_A[5][1] * mat_B[1][29] +
                  mat_A[5][2] * mat_B[2][29] +
                  mat_A[5][3] * mat_B[3][29] +
                  mat_A[5][4] * mat_B[4][29] +
                  mat_A[5][5] * mat_B[5][29] +
                  mat_A[5][6] * mat_B[6][29] +
                  mat_A[5][7] * mat_B[7][29] +
                  mat_A[5][8] * mat_B[8][29] +
                  mat_A[5][9] * mat_B[9][29] +
                  mat_A[5][10] * mat_B[10][29] +
                  mat_A[5][11] * mat_B[11][29] +
                  mat_A[5][12] * mat_B[12][29] +
                  mat_A[5][13] * mat_B[13][29] +
                  mat_A[5][14] * mat_B[14][29] +
                  mat_A[5][15] * mat_B[15][29] +
                  mat_A[5][16] * mat_B[16][29] +
                  mat_A[5][17] * mat_B[17][29] +
                  mat_A[5][18] * mat_B[18][29] +
                  mat_A[5][19] * mat_B[19][29] +
                  mat_A[5][20] * mat_B[20][29] +
                  mat_A[5][21] * mat_B[21][29] +
                  mat_A[5][22] * mat_B[22][29] +
                  mat_A[5][23] * mat_B[23][29] +
                  mat_A[5][24] * mat_B[24][29] +
                  mat_A[5][25] * mat_B[25][29] +
                  mat_A[5][26] * mat_B[26][29] +
                  mat_A[5][27] * mat_B[27][29] +
                  mat_A[5][28] * mat_B[28][29] +
                  mat_A[5][29] * mat_B[29][29] +
                  mat_A[5][30] * mat_B[30][29] +
                  mat_A[5][31] * mat_B[31][29];
    mat_C[5][30] <= 
                  mat_A[5][0] * mat_B[0][30] +
                  mat_A[5][1] * mat_B[1][30] +
                  mat_A[5][2] * mat_B[2][30] +
                  mat_A[5][3] * mat_B[3][30] +
                  mat_A[5][4] * mat_B[4][30] +
                  mat_A[5][5] * mat_B[5][30] +
                  mat_A[5][6] * mat_B[6][30] +
                  mat_A[5][7] * mat_B[7][30] +
                  mat_A[5][8] * mat_B[8][30] +
                  mat_A[5][9] * mat_B[9][30] +
                  mat_A[5][10] * mat_B[10][30] +
                  mat_A[5][11] * mat_B[11][30] +
                  mat_A[5][12] * mat_B[12][30] +
                  mat_A[5][13] * mat_B[13][30] +
                  mat_A[5][14] * mat_B[14][30] +
                  mat_A[5][15] * mat_B[15][30] +
                  mat_A[5][16] * mat_B[16][30] +
                  mat_A[5][17] * mat_B[17][30] +
                  mat_A[5][18] * mat_B[18][30] +
                  mat_A[5][19] * mat_B[19][30] +
                  mat_A[5][20] * mat_B[20][30] +
                  mat_A[5][21] * mat_B[21][30] +
                  mat_A[5][22] * mat_B[22][30] +
                  mat_A[5][23] * mat_B[23][30] +
                  mat_A[5][24] * mat_B[24][30] +
                  mat_A[5][25] * mat_B[25][30] +
                  mat_A[5][26] * mat_B[26][30] +
                  mat_A[5][27] * mat_B[27][30] +
                  mat_A[5][28] * mat_B[28][30] +
                  mat_A[5][29] * mat_B[29][30] +
                  mat_A[5][30] * mat_B[30][30] +
                  mat_A[5][31] * mat_B[31][30];
    mat_C[5][31] <= 
                  mat_A[5][0] * mat_B[0][31] +
                  mat_A[5][1] * mat_B[1][31] +
                  mat_A[5][2] * mat_B[2][31] +
                  mat_A[5][3] * mat_B[3][31] +
                  mat_A[5][4] * mat_B[4][31] +
                  mat_A[5][5] * mat_B[5][31] +
                  mat_A[5][6] * mat_B[6][31] +
                  mat_A[5][7] * mat_B[7][31] +
                  mat_A[5][8] * mat_B[8][31] +
                  mat_A[5][9] * mat_B[9][31] +
                  mat_A[5][10] * mat_B[10][31] +
                  mat_A[5][11] * mat_B[11][31] +
                  mat_A[5][12] * mat_B[12][31] +
                  mat_A[5][13] * mat_B[13][31] +
                  mat_A[5][14] * mat_B[14][31] +
                  mat_A[5][15] * mat_B[15][31] +
                  mat_A[5][16] * mat_B[16][31] +
                  mat_A[5][17] * mat_B[17][31] +
                  mat_A[5][18] * mat_B[18][31] +
                  mat_A[5][19] * mat_B[19][31] +
                  mat_A[5][20] * mat_B[20][31] +
                  mat_A[5][21] * mat_B[21][31] +
                  mat_A[5][22] * mat_B[22][31] +
                  mat_A[5][23] * mat_B[23][31] +
                  mat_A[5][24] * mat_B[24][31] +
                  mat_A[5][25] * mat_B[25][31] +
                  mat_A[5][26] * mat_B[26][31] +
                  mat_A[5][27] * mat_B[27][31] +
                  mat_A[5][28] * mat_B[28][31] +
                  mat_A[5][29] * mat_B[29][31] +
                  mat_A[5][30] * mat_B[30][31] +
                  mat_A[5][31] * mat_B[31][31];
    mat_C[6][0] <= 
                  mat_A[6][0] * mat_B[0][0] +
                  mat_A[6][1] * mat_B[1][0] +
                  mat_A[6][2] * mat_B[2][0] +
                  mat_A[6][3] * mat_B[3][0] +
                  mat_A[6][4] * mat_B[4][0] +
                  mat_A[6][5] * mat_B[5][0] +
                  mat_A[6][6] * mat_B[6][0] +
                  mat_A[6][7] * mat_B[7][0] +
                  mat_A[6][8] * mat_B[8][0] +
                  mat_A[6][9] * mat_B[9][0] +
                  mat_A[6][10] * mat_B[10][0] +
                  mat_A[6][11] * mat_B[11][0] +
                  mat_A[6][12] * mat_B[12][0] +
                  mat_A[6][13] * mat_B[13][0] +
                  mat_A[6][14] * mat_B[14][0] +
                  mat_A[6][15] * mat_B[15][0] +
                  mat_A[6][16] * mat_B[16][0] +
                  mat_A[6][17] * mat_B[17][0] +
                  mat_A[6][18] * mat_B[18][0] +
                  mat_A[6][19] * mat_B[19][0] +
                  mat_A[6][20] * mat_B[20][0] +
                  mat_A[6][21] * mat_B[21][0] +
                  mat_A[6][22] * mat_B[22][0] +
                  mat_A[6][23] * mat_B[23][0] +
                  mat_A[6][24] * mat_B[24][0] +
                  mat_A[6][25] * mat_B[25][0] +
                  mat_A[6][26] * mat_B[26][0] +
                  mat_A[6][27] * mat_B[27][0] +
                  mat_A[6][28] * mat_B[28][0] +
                  mat_A[6][29] * mat_B[29][0] +
                  mat_A[6][30] * mat_B[30][0] +
                  mat_A[6][31] * mat_B[31][0];
    mat_C[6][1] <= 
                  mat_A[6][0] * mat_B[0][1] +
                  mat_A[6][1] * mat_B[1][1] +
                  mat_A[6][2] * mat_B[2][1] +
                  mat_A[6][3] * mat_B[3][1] +
                  mat_A[6][4] * mat_B[4][1] +
                  mat_A[6][5] * mat_B[5][1] +
                  mat_A[6][6] * mat_B[6][1] +
                  mat_A[6][7] * mat_B[7][1] +
                  mat_A[6][8] * mat_B[8][1] +
                  mat_A[6][9] * mat_B[9][1] +
                  mat_A[6][10] * mat_B[10][1] +
                  mat_A[6][11] * mat_B[11][1] +
                  mat_A[6][12] * mat_B[12][1] +
                  mat_A[6][13] * mat_B[13][1] +
                  mat_A[6][14] * mat_B[14][1] +
                  mat_A[6][15] * mat_B[15][1] +
                  mat_A[6][16] * mat_B[16][1] +
                  mat_A[6][17] * mat_B[17][1] +
                  mat_A[6][18] * mat_B[18][1] +
                  mat_A[6][19] * mat_B[19][1] +
                  mat_A[6][20] * mat_B[20][1] +
                  mat_A[6][21] * mat_B[21][1] +
                  mat_A[6][22] * mat_B[22][1] +
                  mat_A[6][23] * mat_B[23][1] +
                  mat_A[6][24] * mat_B[24][1] +
                  mat_A[6][25] * mat_B[25][1] +
                  mat_A[6][26] * mat_B[26][1] +
                  mat_A[6][27] * mat_B[27][1] +
                  mat_A[6][28] * mat_B[28][1] +
                  mat_A[6][29] * mat_B[29][1] +
                  mat_A[6][30] * mat_B[30][1] +
                  mat_A[6][31] * mat_B[31][1];
    mat_C[6][2] <= 
                  mat_A[6][0] * mat_B[0][2] +
                  mat_A[6][1] * mat_B[1][2] +
                  mat_A[6][2] * mat_B[2][2] +
                  mat_A[6][3] * mat_B[3][2] +
                  mat_A[6][4] * mat_B[4][2] +
                  mat_A[6][5] * mat_B[5][2] +
                  mat_A[6][6] * mat_B[6][2] +
                  mat_A[6][7] * mat_B[7][2] +
                  mat_A[6][8] * mat_B[8][2] +
                  mat_A[6][9] * mat_B[9][2] +
                  mat_A[6][10] * mat_B[10][2] +
                  mat_A[6][11] * mat_B[11][2] +
                  mat_A[6][12] * mat_B[12][2] +
                  mat_A[6][13] * mat_B[13][2] +
                  mat_A[6][14] * mat_B[14][2] +
                  mat_A[6][15] * mat_B[15][2] +
                  mat_A[6][16] * mat_B[16][2] +
                  mat_A[6][17] * mat_B[17][2] +
                  mat_A[6][18] * mat_B[18][2] +
                  mat_A[6][19] * mat_B[19][2] +
                  mat_A[6][20] * mat_B[20][2] +
                  mat_A[6][21] * mat_B[21][2] +
                  mat_A[6][22] * mat_B[22][2] +
                  mat_A[6][23] * mat_B[23][2] +
                  mat_A[6][24] * mat_B[24][2] +
                  mat_A[6][25] * mat_B[25][2] +
                  mat_A[6][26] * mat_B[26][2] +
                  mat_A[6][27] * mat_B[27][2] +
                  mat_A[6][28] * mat_B[28][2] +
                  mat_A[6][29] * mat_B[29][2] +
                  mat_A[6][30] * mat_B[30][2] +
                  mat_A[6][31] * mat_B[31][2];
    mat_C[6][3] <= 
                  mat_A[6][0] * mat_B[0][3] +
                  mat_A[6][1] * mat_B[1][3] +
                  mat_A[6][2] * mat_B[2][3] +
                  mat_A[6][3] * mat_B[3][3] +
                  mat_A[6][4] * mat_B[4][3] +
                  mat_A[6][5] * mat_B[5][3] +
                  mat_A[6][6] * mat_B[6][3] +
                  mat_A[6][7] * mat_B[7][3] +
                  mat_A[6][8] * mat_B[8][3] +
                  mat_A[6][9] * mat_B[9][3] +
                  mat_A[6][10] * mat_B[10][3] +
                  mat_A[6][11] * mat_B[11][3] +
                  mat_A[6][12] * mat_B[12][3] +
                  mat_A[6][13] * mat_B[13][3] +
                  mat_A[6][14] * mat_B[14][3] +
                  mat_A[6][15] * mat_B[15][3] +
                  mat_A[6][16] * mat_B[16][3] +
                  mat_A[6][17] * mat_B[17][3] +
                  mat_A[6][18] * mat_B[18][3] +
                  mat_A[6][19] * mat_B[19][3] +
                  mat_A[6][20] * mat_B[20][3] +
                  mat_A[6][21] * mat_B[21][3] +
                  mat_A[6][22] * mat_B[22][3] +
                  mat_A[6][23] * mat_B[23][3] +
                  mat_A[6][24] * mat_B[24][3] +
                  mat_A[6][25] * mat_B[25][3] +
                  mat_A[6][26] * mat_B[26][3] +
                  mat_A[6][27] * mat_B[27][3] +
                  mat_A[6][28] * mat_B[28][3] +
                  mat_A[6][29] * mat_B[29][3] +
                  mat_A[6][30] * mat_B[30][3] +
                  mat_A[6][31] * mat_B[31][3];
    mat_C[6][4] <= 
                  mat_A[6][0] * mat_B[0][4] +
                  mat_A[6][1] * mat_B[1][4] +
                  mat_A[6][2] * mat_B[2][4] +
                  mat_A[6][3] * mat_B[3][4] +
                  mat_A[6][4] * mat_B[4][4] +
                  mat_A[6][5] * mat_B[5][4] +
                  mat_A[6][6] * mat_B[6][4] +
                  mat_A[6][7] * mat_B[7][4] +
                  mat_A[6][8] * mat_B[8][4] +
                  mat_A[6][9] * mat_B[9][4] +
                  mat_A[6][10] * mat_B[10][4] +
                  mat_A[6][11] * mat_B[11][4] +
                  mat_A[6][12] * mat_B[12][4] +
                  mat_A[6][13] * mat_B[13][4] +
                  mat_A[6][14] * mat_B[14][4] +
                  mat_A[6][15] * mat_B[15][4] +
                  mat_A[6][16] * mat_B[16][4] +
                  mat_A[6][17] * mat_B[17][4] +
                  mat_A[6][18] * mat_B[18][4] +
                  mat_A[6][19] * mat_B[19][4] +
                  mat_A[6][20] * mat_B[20][4] +
                  mat_A[6][21] * mat_B[21][4] +
                  mat_A[6][22] * mat_B[22][4] +
                  mat_A[6][23] * mat_B[23][4] +
                  mat_A[6][24] * mat_B[24][4] +
                  mat_A[6][25] * mat_B[25][4] +
                  mat_A[6][26] * mat_B[26][4] +
                  mat_A[6][27] * mat_B[27][4] +
                  mat_A[6][28] * mat_B[28][4] +
                  mat_A[6][29] * mat_B[29][4] +
                  mat_A[6][30] * mat_B[30][4] +
                  mat_A[6][31] * mat_B[31][4];
    mat_C[6][5] <= 
                  mat_A[6][0] * mat_B[0][5] +
                  mat_A[6][1] * mat_B[1][5] +
                  mat_A[6][2] * mat_B[2][5] +
                  mat_A[6][3] * mat_B[3][5] +
                  mat_A[6][4] * mat_B[4][5] +
                  mat_A[6][5] * mat_B[5][5] +
                  mat_A[6][6] * mat_B[6][5] +
                  mat_A[6][7] * mat_B[7][5] +
                  mat_A[6][8] * mat_B[8][5] +
                  mat_A[6][9] * mat_B[9][5] +
                  mat_A[6][10] * mat_B[10][5] +
                  mat_A[6][11] * mat_B[11][5] +
                  mat_A[6][12] * mat_B[12][5] +
                  mat_A[6][13] * mat_B[13][5] +
                  mat_A[6][14] * mat_B[14][5] +
                  mat_A[6][15] * mat_B[15][5] +
                  mat_A[6][16] * mat_B[16][5] +
                  mat_A[6][17] * mat_B[17][5] +
                  mat_A[6][18] * mat_B[18][5] +
                  mat_A[6][19] * mat_B[19][5] +
                  mat_A[6][20] * mat_B[20][5] +
                  mat_A[6][21] * mat_B[21][5] +
                  mat_A[6][22] * mat_B[22][5] +
                  mat_A[6][23] * mat_B[23][5] +
                  mat_A[6][24] * mat_B[24][5] +
                  mat_A[6][25] * mat_B[25][5] +
                  mat_A[6][26] * mat_B[26][5] +
                  mat_A[6][27] * mat_B[27][5] +
                  mat_A[6][28] * mat_B[28][5] +
                  mat_A[6][29] * mat_B[29][5] +
                  mat_A[6][30] * mat_B[30][5] +
                  mat_A[6][31] * mat_B[31][5];
    mat_C[6][6] <= 
                  mat_A[6][0] * mat_B[0][6] +
                  mat_A[6][1] * mat_B[1][6] +
                  mat_A[6][2] * mat_B[2][6] +
                  mat_A[6][3] * mat_B[3][6] +
                  mat_A[6][4] * mat_B[4][6] +
                  mat_A[6][5] * mat_B[5][6] +
                  mat_A[6][6] * mat_B[6][6] +
                  mat_A[6][7] * mat_B[7][6] +
                  mat_A[6][8] * mat_B[8][6] +
                  mat_A[6][9] * mat_B[9][6] +
                  mat_A[6][10] * mat_B[10][6] +
                  mat_A[6][11] * mat_B[11][6] +
                  mat_A[6][12] * mat_B[12][6] +
                  mat_A[6][13] * mat_B[13][6] +
                  mat_A[6][14] * mat_B[14][6] +
                  mat_A[6][15] * mat_B[15][6] +
                  mat_A[6][16] * mat_B[16][6] +
                  mat_A[6][17] * mat_B[17][6] +
                  mat_A[6][18] * mat_B[18][6] +
                  mat_A[6][19] * mat_B[19][6] +
                  mat_A[6][20] * mat_B[20][6] +
                  mat_A[6][21] * mat_B[21][6] +
                  mat_A[6][22] * mat_B[22][6] +
                  mat_A[6][23] * mat_B[23][6] +
                  mat_A[6][24] * mat_B[24][6] +
                  mat_A[6][25] * mat_B[25][6] +
                  mat_A[6][26] * mat_B[26][6] +
                  mat_A[6][27] * mat_B[27][6] +
                  mat_A[6][28] * mat_B[28][6] +
                  mat_A[6][29] * mat_B[29][6] +
                  mat_A[6][30] * mat_B[30][6] +
                  mat_A[6][31] * mat_B[31][6];
    mat_C[6][7] <= 
                  mat_A[6][0] * mat_B[0][7] +
                  mat_A[6][1] * mat_B[1][7] +
                  mat_A[6][2] * mat_B[2][7] +
                  mat_A[6][3] * mat_B[3][7] +
                  mat_A[6][4] * mat_B[4][7] +
                  mat_A[6][5] * mat_B[5][7] +
                  mat_A[6][6] * mat_B[6][7] +
                  mat_A[6][7] * mat_B[7][7] +
                  mat_A[6][8] * mat_B[8][7] +
                  mat_A[6][9] * mat_B[9][7] +
                  mat_A[6][10] * mat_B[10][7] +
                  mat_A[6][11] * mat_B[11][7] +
                  mat_A[6][12] * mat_B[12][7] +
                  mat_A[6][13] * mat_B[13][7] +
                  mat_A[6][14] * mat_B[14][7] +
                  mat_A[6][15] * mat_B[15][7] +
                  mat_A[6][16] * mat_B[16][7] +
                  mat_A[6][17] * mat_B[17][7] +
                  mat_A[6][18] * mat_B[18][7] +
                  mat_A[6][19] * mat_B[19][7] +
                  mat_A[6][20] * mat_B[20][7] +
                  mat_A[6][21] * mat_B[21][7] +
                  mat_A[6][22] * mat_B[22][7] +
                  mat_A[6][23] * mat_B[23][7] +
                  mat_A[6][24] * mat_B[24][7] +
                  mat_A[6][25] * mat_B[25][7] +
                  mat_A[6][26] * mat_B[26][7] +
                  mat_A[6][27] * mat_B[27][7] +
                  mat_A[6][28] * mat_B[28][7] +
                  mat_A[6][29] * mat_B[29][7] +
                  mat_A[6][30] * mat_B[30][7] +
                  mat_A[6][31] * mat_B[31][7];
    mat_C[6][8] <= 
                  mat_A[6][0] * mat_B[0][8] +
                  mat_A[6][1] * mat_B[1][8] +
                  mat_A[6][2] * mat_B[2][8] +
                  mat_A[6][3] * mat_B[3][8] +
                  mat_A[6][4] * mat_B[4][8] +
                  mat_A[6][5] * mat_B[5][8] +
                  mat_A[6][6] * mat_B[6][8] +
                  mat_A[6][7] * mat_B[7][8] +
                  mat_A[6][8] * mat_B[8][8] +
                  mat_A[6][9] * mat_B[9][8] +
                  mat_A[6][10] * mat_B[10][8] +
                  mat_A[6][11] * mat_B[11][8] +
                  mat_A[6][12] * mat_B[12][8] +
                  mat_A[6][13] * mat_B[13][8] +
                  mat_A[6][14] * mat_B[14][8] +
                  mat_A[6][15] * mat_B[15][8] +
                  mat_A[6][16] * mat_B[16][8] +
                  mat_A[6][17] * mat_B[17][8] +
                  mat_A[6][18] * mat_B[18][8] +
                  mat_A[6][19] * mat_B[19][8] +
                  mat_A[6][20] * mat_B[20][8] +
                  mat_A[6][21] * mat_B[21][8] +
                  mat_A[6][22] * mat_B[22][8] +
                  mat_A[6][23] * mat_B[23][8] +
                  mat_A[6][24] * mat_B[24][8] +
                  mat_A[6][25] * mat_B[25][8] +
                  mat_A[6][26] * mat_B[26][8] +
                  mat_A[6][27] * mat_B[27][8] +
                  mat_A[6][28] * mat_B[28][8] +
                  mat_A[6][29] * mat_B[29][8] +
                  mat_A[6][30] * mat_B[30][8] +
                  mat_A[6][31] * mat_B[31][8];
    mat_C[6][9] <= 
                  mat_A[6][0] * mat_B[0][9] +
                  mat_A[6][1] * mat_B[1][9] +
                  mat_A[6][2] * mat_B[2][9] +
                  mat_A[6][3] * mat_B[3][9] +
                  mat_A[6][4] * mat_B[4][9] +
                  mat_A[6][5] * mat_B[5][9] +
                  mat_A[6][6] * mat_B[6][9] +
                  mat_A[6][7] * mat_B[7][9] +
                  mat_A[6][8] * mat_B[8][9] +
                  mat_A[6][9] * mat_B[9][9] +
                  mat_A[6][10] * mat_B[10][9] +
                  mat_A[6][11] * mat_B[11][9] +
                  mat_A[6][12] * mat_B[12][9] +
                  mat_A[6][13] * mat_B[13][9] +
                  mat_A[6][14] * mat_B[14][9] +
                  mat_A[6][15] * mat_B[15][9] +
                  mat_A[6][16] * mat_B[16][9] +
                  mat_A[6][17] * mat_B[17][9] +
                  mat_A[6][18] * mat_B[18][9] +
                  mat_A[6][19] * mat_B[19][9] +
                  mat_A[6][20] * mat_B[20][9] +
                  mat_A[6][21] * mat_B[21][9] +
                  mat_A[6][22] * mat_B[22][9] +
                  mat_A[6][23] * mat_B[23][9] +
                  mat_A[6][24] * mat_B[24][9] +
                  mat_A[6][25] * mat_B[25][9] +
                  mat_A[6][26] * mat_B[26][9] +
                  mat_A[6][27] * mat_B[27][9] +
                  mat_A[6][28] * mat_B[28][9] +
                  mat_A[6][29] * mat_B[29][9] +
                  mat_A[6][30] * mat_B[30][9] +
                  mat_A[6][31] * mat_B[31][9];
    mat_C[6][10] <= 
                  mat_A[6][0] * mat_B[0][10] +
                  mat_A[6][1] * mat_B[1][10] +
                  mat_A[6][2] * mat_B[2][10] +
                  mat_A[6][3] * mat_B[3][10] +
                  mat_A[6][4] * mat_B[4][10] +
                  mat_A[6][5] * mat_B[5][10] +
                  mat_A[6][6] * mat_B[6][10] +
                  mat_A[6][7] * mat_B[7][10] +
                  mat_A[6][8] * mat_B[8][10] +
                  mat_A[6][9] * mat_B[9][10] +
                  mat_A[6][10] * mat_B[10][10] +
                  mat_A[6][11] * mat_B[11][10] +
                  mat_A[6][12] * mat_B[12][10] +
                  mat_A[6][13] * mat_B[13][10] +
                  mat_A[6][14] * mat_B[14][10] +
                  mat_A[6][15] * mat_B[15][10] +
                  mat_A[6][16] * mat_B[16][10] +
                  mat_A[6][17] * mat_B[17][10] +
                  mat_A[6][18] * mat_B[18][10] +
                  mat_A[6][19] * mat_B[19][10] +
                  mat_A[6][20] * mat_B[20][10] +
                  mat_A[6][21] * mat_B[21][10] +
                  mat_A[6][22] * mat_B[22][10] +
                  mat_A[6][23] * mat_B[23][10] +
                  mat_A[6][24] * mat_B[24][10] +
                  mat_A[6][25] * mat_B[25][10] +
                  mat_A[6][26] * mat_B[26][10] +
                  mat_A[6][27] * mat_B[27][10] +
                  mat_A[6][28] * mat_B[28][10] +
                  mat_A[6][29] * mat_B[29][10] +
                  mat_A[6][30] * mat_B[30][10] +
                  mat_A[6][31] * mat_B[31][10];
    mat_C[6][11] <= 
                  mat_A[6][0] * mat_B[0][11] +
                  mat_A[6][1] * mat_B[1][11] +
                  mat_A[6][2] * mat_B[2][11] +
                  mat_A[6][3] * mat_B[3][11] +
                  mat_A[6][4] * mat_B[4][11] +
                  mat_A[6][5] * mat_B[5][11] +
                  mat_A[6][6] * mat_B[6][11] +
                  mat_A[6][7] * mat_B[7][11] +
                  mat_A[6][8] * mat_B[8][11] +
                  mat_A[6][9] * mat_B[9][11] +
                  mat_A[6][10] * mat_B[10][11] +
                  mat_A[6][11] * mat_B[11][11] +
                  mat_A[6][12] * mat_B[12][11] +
                  mat_A[6][13] * mat_B[13][11] +
                  mat_A[6][14] * mat_B[14][11] +
                  mat_A[6][15] * mat_B[15][11] +
                  mat_A[6][16] * mat_B[16][11] +
                  mat_A[6][17] * mat_B[17][11] +
                  mat_A[6][18] * mat_B[18][11] +
                  mat_A[6][19] * mat_B[19][11] +
                  mat_A[6][20] * mat_B[20][11] +
                  mat_A[6][21] * mat_B[21][11] +
                  mat_A[6][22] * mat_B[22][11] +
                  mat_A[6][23] * mat_B[23][11] +
                  mat_A[6][24] * mat_B[24][11] +
                  mat_A[6][25] * mat_B[25][11] +
                  mat_A[6][26] * mat_B[26][11] +
                  mat_A[6][27] * mat_B[27][11] +
                  mat_A[6][28] * mat_B[28][11] +
                  mat_A[6][29] * mat_B[29][11] +
                  mat_A[6][30] * mat_B[30][11] +
                  mat_A[6][31] * mat_B[31][11];
    mat_C[6][12] <= 
                  mat_A[6][0] * mat_B[0][12] +
                  mat_A[6][1] * mat_B[1][12] +
                  mat_A[6][2] * mat_B[2][12] +
                  mat_A[6][3] * mat_B[3][12] +
                  mat_A[6][4] * mat_B[4][12] +
                  mat_A[6][5] * mat_B[5][12] +
                  mat_A[6][6] * mat_B[6][12] +
                  mat_A[6][7] * mat_B[7][12] +
                  mat_A[6][8] * mat_B[8][12] +
                  mat_A[6][9] * mat_B[9][12] +
                  mat_A[6][10] * mat_B[10][12] +
                  mat_A[6][11] * mat_B[11][12] +
                  mat_A[6][12] * mat_B[12][12] +
                  mat_A[6][13] * mat_B[13][12] +
                  mat_A[6][14] * mat_B[14][12] +
                  mat_A[6][15] * mat_B[15][12] +
                  mat_A[6][16] * mat_B[16][12] +
                  mat_A[6][17] * mat_B[17][12] +
                  mat_A[6][18] * mat_B[18][12] +
                  mat_A[6][19] * mat_B[19][12] +
                  mat_A[6][20] * mat_B[20][12] +
                  mat_A[6][21] * mat_B[21][12] +
                  mat_A[6][22] * mat_B[22][12] +
                  mat_A[6][23] * mat_B[23][12] +
                  mat_A[6][24] * mat_B[24][12] +
                  mat_A[6][25] * mat_B[25][12] +
                  mat_A[6][26] * mat_B[26][12] +
                  mat_A[6][27] * mat_B[27][12] +
                  mat_A[6][28] * mat_B[28][12] +
                  mat_A[6][29] * mat_B[29][12] +
                  mat_A[6][30] * mat_B[30][12] +
                  mat_A[6][31] * mat_B[31][12];
    mat_C[6][13] <= 
                  mat_A[6][0] * mat_B[0][13] +
                  mat_A[6][1] * mat_B[1][13] +
                  mat_A[6][2] * mat_B[2][13] +
                  mat_A[6][3] * mat_B[3][13] +
                  mat_A[6][4] * mat_B[4][13] +
                  mat_A[6][5] * mat_B[5][13] +
                  mat_A[6][6] * mat_B[6][13] +
                  mat_A[6][7] * mat_B[7][13] +
                  mat_A[6][8] * mat_B[8][13] +
                  mat_A[6][9] * mat_B[9][13] +
                  mat_A[6][10] * mat_B[10][13] +
                  mat_A[6][11] * mat_B[11][13] +
                  mat_A[6][12] * mat_B[12][13] +
                  mat_A[6][13] * mat_B[13][13] +
                  mat_A[6][14] * mat_B[14][13] +
                  mat_A[6][15] * mat_B[15][13] +
                  mat_A[6][16] * mat_B[16][13] +
                  mat_A[6][17] * mat_B[17][13] +
                  mat_A[6][18] * mat_B[18][13] +
                  mat_A[6][19] * mat_B[19][13] +
                  mat_A[6][20] * mat_B[20][13] +
                  mat_A[6][21] * mat_B[21][13] +
                  mat_A[6][22] * mat_B[22][13] +
                  mat_A[6][23] * mat_B[23][13] +
                  mat_A[6][24] * mat_B[24][13] +
                  mat_A[6][25] * mat_B[25][13] +
                  mat_A[6][26] * mat_B[26][13] +
                  mat_A[6][27] * mat_B[27][13] +
                  mat_A[6][28] * mat_B[28][13] +
                  mat_A[6][29] * mat_B[29][13] +
                  mat_A[6][30] * mat_B[30][13] +
                  mat_A[6][31] * mat_B[31][13];
    mat_C[6][14] <= 
                  mat_A[6][0] * mat_B[0][14] +
                  mat_A[6][1] * mat_B[1][14] +
                  mat_A[6][2] * mat_B[2][14] +
                  mat_A[6][3] * mat_B[3][14] +
                  mat_A[6][4] * mat_B[4][14] +
                  mat_A[6][5] * mat_B[5][14] +
                  mat_A[6][6] * mat_B[6][14] +
                  mat_A[6][7] * mat_B[7][14] +
                  mat_A[6][8] * mat_B[8][14] +
                  mat_A[6][9] * mat_B[9][14] +
                  mat_A[6][10] * mat_B[10][14] +
                  mat_A[6][11] * mat_B[11][14] +
                  mat_A[6][12] * mat_B[12][14] +
                  mat_A[6][13] * mat_B[13][14] +
                  mat_A[6][14] * mat_B[14][14] +
                  mat_A[6][15] * mat_B[15][14] +
                  mat_A[6][16] * mat_B[16][14] +
                  mat_A[6][17] * mat_B[17][14] +
                  mat_A[6][18] * mat_B[18][14] +
                  mat_A[6][19] * mat_B[19][14] +
                  mat_A[6][20] * mat_B[20][14] +
                  mat_A[6][21] * mat_B[21][14] +
                  mat_A[6][22] * mat_B[22][14] +
                  mat_A[6][23] * mat_B[23][14] +
                  mat_A[6][24] * mat_B[24][14] +
                  mat_A[6][25] * mat_B[25][14] +
                  mat_A[6][26] * mat_B[26][14] +
                  mat_A[6][27] * mat_B[27][14] +
                  mat_A[6][28] * mat_B[28][14] +
                  mat_A[6][29] * mat_B[29][14] +
                  mat_A[6][30] * mat_B[30][14] +
                  mat_A[6][31] * mat_B[31][14];
    mat_C[6][15] <= 
                  mat_A[6][0] * mat_B[0][15] +
                  mat_A[6][1] * mat_B[1][15] +
                  mat_A[6][2] * mat_B[2][15] +
                  mat_A[6][3] * mat_B[3][15] +
                  mat_A[6][4] * mat_B[4][15] +
                  mat_A[6][5] * mat_B[5][15] +
                  mat_A[6][6] * mat_B[6][15] +
                  mat_A[6][7] * mat_B[7][15] +
                  mat_A[6][8] * mat_B[8][15] +
                  mat_A[6][9] * mat_B[9][15] +
                  mat_A[6][10] * mat_B[10][15] +
                  mat_A[6][11] * mat_B[11][15] +
                  mat_A[6][12] * mat_B[12][15] +
                  mat_A[6][13] * mat_B[13][15] +
                  mat_A[6][14] * mat_B[14][15] +
                  mat_A[6][15] * mat_B[15][15] +
                  mat_A[6][16] * mat_B[16][15] +
                  mat_A[6][17] * mat_B[17][15] +
                  mat_A[6][18] * mat_B[18][15] +
                  mat_A[6][19] * mat_B[19][15] +
                  mat_A[6][20] * mat_B[20][15] +
                  mat_A[6][21] * mat_B[21][15] +
                  mat_A[6][22] * mat_B[22][15] +
                  mat_A[6][23] * mat_B[23][15] +
                  mat_A[6][24] * mat_B[24][15] +
                  mat_A[6][25] * mat_B[25][15] +
                  mat_A[6][26] * mat_B[26][15] +
                  mat_A[6][27] * mat_B[27][15] +
                  mat_A[6][28] * mat_B[28][15] +
                  mat_A[6][29] * mat_B[29][15] +
                  mat_A[6][30] * mat_B[30][15] +
                  mat_A[6][31] * mat_B[31][15];
    mat_C[6][16] <= 
                  mat_A[6][0] * mat_B[0][16] +
                  mat_A[6][1] * mat_B[1][16] +
                  mat_A[6][2] * mat_B[2][16] +
                  mat_A[6][3] * mat_B[3][16] +
                  mat_A[6][4] * mat_B[4][16] +
                  mat_A[6][5] * mat_B[5][16] +
                  mat_A[6][6] * mat_B[6][16] +
                  mat_A[6][7] * mat_B[7][16] +
                  mat_A[6][8] * mat_B[8][16] +
                  mat_A[6][9] * mat_B[9][16] +
                  mat_A[6][10] * mat_B[10][16] +
                  mat_A[6][11] * mat_B[11][16] +
                  mat_A[6][12] * mat_B[12][16] +
                  mat_A[6][13] * mat_B[13][16] +
                  mat_A[6][14] * mat_B[14][16] +
                  mat_A[6][15] * mat_B[15][16] +
                  mat_A[6][16] * mat_B[16][16] +
                  mat_A[6][17] * mat_B[17][16] +
                  mat_A[6][18] * mat_B[18][16] +
                  mat_A[6][19] * mat_B[19][16] +
                  mat_A[6][20] * mat_B[20][16] +
                  mat_A[6][21] * mat_B[21][16] +
                  mat_A[6][22] * mat_B[22][16] +
                  mat_A[6][23] * mat_B[23][16] +
                  mat_A[6][24] * mat_B[24][16] +
                  mat_A[6][25] * mat_B[25][16] +
                  mat_A[6][26] * mat_B[26][16] +
                  mat_A[6][27] * mat_B[27][16] +
                  mat_A[6][28] * mat_B[28][16] +
                  mat_A[6][29] * mat_B[29][16] +
                  mat_A[6][30] * mat_B[30][16] +
                  mat_A[6][31] * mat_B[31][16];
    mat_C[6][17] <= 
                  mat_A[6][0] * mat_B[0][17] +
                  mat_A[6][1] * mat_B[1][17] +
                  mat_A[6][2] * mat_B[2][17] +
                  mat_A[6][3] * mat_B[3][17] +
                  mat_A[6][4] * mat_B[4][17] +
                  mat_A[6][5] * mat_B[5][17] +
                  mat_A[6][6] * mat_B[6][17] +
                  mat_A[6][7] * mat_B[7][17] +
                  mat_A[6][8] * mat_B[8][17] +
                  mat_A[6][9] * mat_B[9][17] +
                  mat_A[6][10] * mat_B[10][17] +
                  mat_A[6][11] * mat_B[11][17] +
                  mat_A[6][12] * mat_B[12][17] +
                  mat_A[6][13] * mat_B[13][17] +
                  mat_A[6][14] * mat_B[14][17] +
                  mat_A[6][15] * mat_B[15][17] +
                  mat_A[6][16] * mat_B[16][17] +
                  mat_A[6][17] * mat_B[17][17] +
                  mat_A[6][18] * mat_B[18][17] +
                  mat_A[6][19] * mat_B[19][17] +
                  mat_A[6][20] * mat_B[20][17] +
                  mat_A[6][21] * mat_B[21][17] +
                  mat_A[6][22] * mat_B[22][17] +
                  mat_A[6][23] * mat_B[23][17] +
                  mat_A[6][24] * mat_B[24][17] +
                  mat_A[6][25] * mat_B[25][17] +
                  mat_A[6][26] * mat_B[26][17] +
                  mat_A[6][27] * mat_B[27][17] +
                  mat_A[6][28] * mat_B[28][17] +
                  mat_A[6][29] * mat_B[29][17] +
                  mat_A[6][30] * mat_B[30][17] +
                  mat_A[6][31] * mat_B[31][17];
    mat_C[6][18] <= 
                  mat_A[6][0] * mat_B[0][18] +
                  mat_A[6][1] * mat_B[1][18] +
                  mat_A[6][2] * mat_B[2][18] +
                  mat_A[6][3] * mat_B[3][18] +
                  mat_A[6][4] * mat_B[4][18] +
                  mat_A[6][5] * mat_B[5][18] +
                  mat_A[6][6] * mat_B[6][18] +
                  mat_A[6][7] * mat_B[7][18] +
                  mat_A[6][8] * mat_B[8][18] +
                  mat_A[6][9] * mat_B[9][18] +
                  mat_A[6][10] * mat_B[10][18] +
                  mat_A[6][11] * mat_B[11][18] +
                  mat_A[6][12] * mat_B[12][18] +
                  mat_A[6][13] * mat_B[13][18] +
                  mat_A[6][14] * mat_B[14][18] +
                  mat_A[6][15] * mat_B[15][18] +
                  mat_A[6][16] * mat_B[16][18] +
                  mat_A[6][17] * mat_B[17][18] +
                  mat_A[6][18] * mat_B[18][18] +
                  mat_A[6][19] * mat_B[19][18] +
                  mat_A[6][20] * mat_B[20][18] +
                  mat_A[6][21] * mat_B[21][18] +
                  mat_A[6][22] * mat_B[22][18] +
                  mat_A[6][23] * mat_B[23][18] +
                  mat_A[6][24] * mat_B[24][18] +
                  mat_A[6][25] * mat_B[25][18] +
                  mat_A[6][26] * mat_B[26][18] +
                  mat_A[6][27] * mat_B[27][18] +
                  mat_A[6][28] * mat_B[28][18] +
                  mat_A[6][29] * mat_B[29][18] +
                  mat_A[6][30] * mat_B[30][18] +
                  mat_A[6][31] * mat_B[31][18];
    mat_C[6][19] <= 
                  mat_A[6][0] * mat_B[0][19] +
                  mat_A[6][1] * mat_B[1][19] +
                  mat_A[6][2] * mat_B[2][19] +
                  mat_A[6][3] * mat_B[3][19] +
                  mat_A[6][4] * mat_B[4][19] +
                  mat_A[6][5] * mat_B[5][19] +
                  mat_A[6][6] * mat_B[6][19] +
                  mat_A[6][7] * mat_B[7][19] +
                  mat_A[6][8] * mat_B[8][19] +
                  mat_A[6][9] * mat_B[9][19] +
                  mat_A[6][10] * mat_B[10][19] +
                  mat_A[6][11] * mat_B[11][19] +
                  mat_A[6][12] * mat_B[12][19] +
                  mat_A[6][13] * mat_B[13][19] +
                  mat_A[6][14] * mat_B[14][19] +
                  mat_A[6][15] * mat_B[15][19] +
                  mat_A[6][16] * mat_B[16][19] +
                  mat_A[6][17] * mat_B[17][19] +
                  mat_A[6][18] * mat_B[18][19] +
                  mat_A[6][19] * mat_B[19][19] +
                  mat_A[6][20] * mat_B[20][19] +
                  mat_A[6][21] * mat_B[21][19] +
                  mat_A[6][22] * mat_B[22][19] +
                  mat_A[6][23] * mat_B[23][19] +
                  mat_A[6][24] * mat_B[24][19] +
                  mat_A[6][25] * mat_B[25][19] +
                  mat_A[6][26] * mat_B[26][19] +
                  mat_A[6][27] * mat_B[27][19] +
                  mat_A[6][28] * mat_B[28][19] +
                  mat_A[6][29] * mat_B[29][19] +
                  mat_A[6][30] * mat_B[30][19] +
                  mat_A[6][31] * mat_B[31][19];
    mat_C[6][20] <= 
                  mat_A[6][0] * mat_B[0][20] +
                  mat_A[6][1] * mat_B[1][20] +
                  mat_A[6][2] * mat_B[2][20] +
                  mat_A[6][3] * mat_B[3][20] +
                  mat_A[6][4] * mat_B[4][20] +
                  mat_A[6][5] * mat_B[5][20] +
                  mat_A[6][6] * mat_B[6][20] +
                  mat_A[6][7] * mat_B[7][20] +
                  mat_A[6][8] * mat_B[8][20] +
                  mat_A[6][9] * mat_B[9][20] +
                  mat_A[6][10] * mat_B[10][20] +
                  mat_A[6][11] * mat_B[11][20] +
                  mat_A[6][12] * mat_B[12][20] +
                  mat_A[6][13] * mat_B[13][20] +
                  mat_A[6][14] * mat_B[14][20] +
                  mat_A[6][15] * mat_B[15][20] +
                  mat_A[6][16] * mat_B[16][20] +
                  mat_A[6][17] * mat_B[17][20] +
                  mat_A[6][18] * mat_B[18][20] +
                  mat_A[6][19] * mat_B[19][20] +
                  mat_A[6][20] * mat_B[20][20] +
                  mat_A[6][21] * mat_B[21][20] +
                  mat_A[6][22] * mat_B[22][20] +
                  mat_A[6][23] * mat_B[23][20] +
                  mat_A[6][24] * mat_B[24][20] +
                  mat_A[6][25] * mat_B[25][20] +
                  mat_A[6][26] * mat_B[26][20] +
                  mat_A[6][27] * mat_B[27][20] +
                  mat_A[6][28] * mat_B[28][20] +
                  mat_A[6][29] * mat_B[29][20] +
                  mat_A[6][30] * mat_B[30][20] +
                  mat_A[6][31] * mat_B[31][20];
    mat_C[6][21] <= 
                  mat_A[6][0] * mat_B[0][21] +
                  mat_A[6][1] * mat_B[1][21] +
                  mat_A[6][2] * mat_B[2][21] +
                  mat_A[6][3] * mat_B[3][21] +
                  mat_A[6][4] * mat_B[4][21] +
                  mat_A[6][5] * mat_B[5][21] +
                  mat_A[6][6] * mat_B[6][21] +
                  mat_A[6][7] * mat_B[7][21] +
                  mat_A[6][8] * mat_B[8][21] +
                  mat_A[6][9] * mat_B[9][21] +
                  mat_A[6][10] * mat_B[10][21] +
                  mat_A[6][11] * mat_B[11][21] +
                  mat_A[6][12] * mat_B[12][21] +
                  mat_A[6][13] * mat_B[13][21] +
                  mat_A[6][14] * mat_B[14][21] +
                  mat_A[6][15] * mat_B[15][21] +
                  mat_A[6][16] * mat_B[16][21] +
                  mat_A[6][17] * mat_B[17][21] +
                  mat_A[6][18] * mat_B[18][21] +
                  mat_A[6][19] * mat_B[19][21] +
                  mat_A[6][20] * mat_B[20][21] +
                  mat_A[6][21] * mat_B[21][21] +
                  mat_A[6][22] * mat_B[22][21] +
                  mat_A[6][23] * mat_B[23][21] +
                  mat_A[6][24] * mat_B[24][21] +
                  mat_A[6][25] * mat_B[25][21] +
                  mat_A[6][26] * mat_B[26][21] +
                  mat_A[6][27] * mat_B[27][21] +
                  mat_A[6][28] * mat_B[28][21] +
                  mat_A[6][29] * mat_B[29][21] +
                  mat_A[6][30] * mat_B[30][21] +
                  mat_A[6][31] * mat_B[31][21];
    mat_C[6][22] <= 
                  mat_A[6][0] * mat_B[0][22] +
                  mat_A[6][1] * mat_B[1][22] +
                  mat_A[6][2] * mat_B[2][22] +
                  mat_A[6][3] * mat_B[3][22] +
                  mat_A[6][4] * mat_B[4][22] +
                  mat_A[6][5] * mat_B[5][22] +
                  mat_A[6][6] * mat_B[6][22] +
                  mat_A[6][7] * mat_B[7][22] +
                  mat_A[6][8] * mat_B[8][22] +
                  mat_A[6][9] * mat_B[9][22] +
                  mat_A[6][10] * mat_B[10][22] +
                  mat_A[6][11] * mat_B[11][22] +
                  mat_A[6][12] * mat_B[12][22] +
                  mat_A[6][13] * mat_B[13][22] +
                  mat_A[6][14] * mat_B[14][22] +
                  mat_A[6][15] * mat_B[15][22] +
                  mat_A[6][16] * mat_B[16][22] +
                  mat_A[6][17] * mat_B[17][22] +
                  mat_A[6][18] * mat_B[18][22] +
                  mat_A[6][19] * mat_B[19][22] +
                  mat_A[6][20] * mat_B[20][22] +
                  mat_A[6][21] * mat_B[21][22] +
                  mat_A[6][22] * mat_B[22][22] +
                  mat_A[6][23] * mat_B[23][22] +
                  mat_A[6][24] * mat_B[24][22] +
                  mat_A[6][25] * mat_B[25][22] +
                  mat_A[6][26] * mat_B[26][22] +
                  mat_A[6][27] * mat_B[27][22] +
                  mat_A[6][28] * mat_B[28][22] +
                  mat_A[6][29] * mat_B[29][22] +
                  mat_A[6][30] * mat_B[30][22] +
                  mat_A[6][31] * mat_B[31][22];
    mat_C[6][23] <= 
                  mat_A[6][0] * mat_B[0][23] +
                  mat_A[6][1] * mat_B[1][23] +
                  mat_A[6][2] * mat_B[2][23] +
                  mat_A[6][3] * mat_B[3][23] +
                  mat_A[6][4] * mat_B[4][23] +
                  mat_A[6][5] * mat_B[5][23] +
                  mat_A[6][6] * mat_B[6][23] +
                  mat_A[6][7] * mat_B[7][23] +
                  mat_A[6][8] * mat_B[8][23] +
                  mat_A[6][9] * mat_B[9][23] +
                  mat_A[6][10] * mat_B[10][23] +
                  mat_A[6][11] * mat_B[11][23] +
                  mat_A[6][12] * mat_B[12][23] +
                  mat_A[6][13] * mat_B[13][23] +
                  mat_A[6][14] * mat_B[14][23] +
                  mat_A[6][15] * mat_B[15][23] +
                  mat_A[6][16] * mat_B[16][23] +
                  mat_A[6][17] * mat_B[17][23] +
                  mat_A[6][18] * mat_B[18][23] +
                  mat_A[6][19] * mat_B[19][23] +
                  mat_A[6][20] * mat_B[20][23] +
                  mat_A[6][21] * mat_B[21][23] +
                  mat_A[6][22] * mat_B[22][23] +
                  mat_A[6][23] * mat_B[23][23] +
                  mat_A[6][24] * mat_B[24][23] +
                  mat_A[6][25] * mat_B[25][23] +
                  mat_A[6][26] * mat_B[26][23] +
                  mat_A[6][27] * mat_B[27][23] +
                  mat_A[6][28] * mat_B[28][23] +
                  mat_A[6][29] * mat_B[29][23] +
                  mat_A[6][30] * mat_B[30][23] +
                  mat_A[6][31] * mat_B[31][23];
    mat_C[6][24] <= 
                  mat_A[6][0] * mat_B[0][24] +
                  mat_A[6][1] * mat_B[1][24] +
                  mat_A[6][2] * mat_B[2][24] +
                  mat_A[6][3] * mat_B[3][24] +
                  mat_A[6][4] * mat_B[4][24] +
                  mat_A[6][5] * mat_B[5][24] +
                  mat_A[6][6] * mat_B[6][24] +
                  mat_A[6][7] * mat_B[7][24] +
                  mat_A[6][8] * mat_B[8][24] +
                  mat_A[6][9] * mat_B[9][24] +
                  mat_A[6][10] * mat_B[10][24] +
                  mat_A[6][11] * mat_B[11][24] +
                  mat_A[6][12] * mat_B[12][24] +
                  mat_A[6][13] * mat_B[13][24] +
                  mat_A[6][14] * mat_B[14][24] +
                  mat_A[6][15] * mat_B[15][24] +
                  mat_A[6][16] * mat_B[16][24] +
                  mat_A[6][17] * mat_B[17][24] +
                  mat_A[6][18] * mat_B[18][24] +
                  mat_A[6][19] * mat_B[19][24] +
                  mat_A[6][20] * mat_B[20][24] +
                  mat_A[6][21] * mat_B[21][24] +
                  mat_A[6][22] * mat_B[22][24] +
                  mat_A[6][23] * mat_B[23][24] +
                  mat_A[6][24] * mat_B[24][24] +
                  mat_A[6][25] * mat_B[25][24] +
                  mat_A[6][26] * mat_B[26][24] +
                  mat_A[6][27] * mat_B[27][24] +
                  mat_A[6][28] * mat_B[28][24] +
                  mat_A[6][29] * mat_B[29][24] +
                  mat_A[6][30] * mat_B[30][24] +
                  mat_A[6][31] * mat_B[31][24];
    mat_C[6][25] <= 
                  mat_A[6][0] * mat_B[0][25] +
                  mat_A[6][1] * mat_B[1][25] +
                  mat_A[6][2] * mat_B[2][25] +
                  mat_A[6][3] * mat_B[3][25] +
                  mat_A[6][4] * mat_B[4][25] +
                  mat_A[6][5] * mat_B[5][25] +
                  mat_A[6][6] * mat_B[6][25] +
                  mat_A[6][7] * mat_B[7][25] +
                  mat_A[6][8] * mat_B[8][25] +
                  mat_A[6][9] * mat_B[9][25] +
                  mat_A[6][10] * mat_B[10][25] +
                  mat_A[6][11] * mat_B[11][25] +
                  mat_A[6][12] * mat_B[12][25] +
                  mat_A[6][13] * mat_B[13][25] +
                  mat_A[6][14] * mat_B[14][25] +
                  mat_A[6][15] * mat_B[15][25] +
                  mat_A[6][16] * mat_B[16][25] +
                  mat_A[6][17] * mat_B[17][25] +
                  mat_A[6][18] * mat_B[18][25] +
                  mat_A[6][19] * mat_B[19][25] +
                  mat_A[6][20] * mat_B[20][25] +
                  mat_A[6][21] * mat_B[21][25] +
                  mat_A[6][22] * mat_B[22][25] +
                  mat_A[6][23] * mat_B[23][25] +
                  mat_A[6][24] * mat_B[24][25] +
                  mat_A[6][25] * mat_B[25][25] +
                  mat_A[6][26] * mat_B[26][25] +
                  mat_A[6][27] * mat_B[27][25] +
                  mat_A[6][28] * mat_B[28][25] +
                  mat_A[6][29] * mat_B[29][25] +
                  mat_A[6][30] * mat_B[30][25] +
                  mat_A[6][31] * mat_B[31][25];
    mat_C[6][26] <= 
                  mat_A[6][0] * mat_B[0][26] +
                  mat_A[6][1] * mat_B[1][26] +
                  mat_A[6][2] * mat_B[2][26] +
                  mat_A[6][3] * mat_B[3][26] +
                  mat_A[6][4] * mat_B[4][26] +
                  mat_A[6][5] * mat_B[5][26] +
                  mat_A[6][6] * mat_B[6][26] +
                  mat_A[6][7] * mat_B[7][26] +
                  mat_A[6][8] * mat_B[8][26] +
                  mat_A[6][9] * mat_B[9][26] +
                  mat_A[6][10] * mat_B[10][26] +
                  mat_A[6][11] * mat_B[11][26] +
                  mat_A[6][12] * mat_B[12][26] +
                  mat_A[6][13] * mat_B[13][26] +
                  mat_A[6][14] * mat_B[14][26] +
                  mat_A[6][15] * mat_B[15][26] +
                  mat_A[6][16] * mat_B[16][26] +
                  mat_A[6][17] * mat_B[17][26] +
                  mat_A[6][18] * mat_B[18][26] +
                  mat_A[6][19] * mat_B[19][26] +
                  mat_A[6][20] * mat_B[20][26] +
                  mat_A[6][21] * mat_B[21][26] +
                  mat_A[6][22] * mat_B[22][26] +
                  mat_A[6][23] * mat_B[23][26] +
                  mat_A[6][24] * mat_B[24][26] +
                  mat_A[6][25] * mat_B[25][26] +
                  mat_A[6][26] * mat_B[26][26] +
                  mat_A[6][27] * mat_B[27][26] +
                  mat_A[6][28] * mat_B[28][26] +
                  mat_A[6][29] * mat_B[29][26] +
                  mat_A[6][30] * mat_B[30][26] +
                  mat_A[6][31] * mat_B[31][26];
    mat_C[6][27] <= 
                  mat_A[6][0] * mat_B[0][27] +
                  mat_A[6][1] * mat_B[1][27] +
                  mat_A[6][2] * mat_B[2][27] +
                  mat_A[6][3] * mat_B[3][27] +
                  mat_A[6][4] * mat_B[4][27] +
                  mat_A[6][5] * mat_B[5][27] +
                  mat_A[6][6] * mat_B[6][27] +
                  mat_A[6][7] * mat_B[7][27] +
                  mat_A[6][8] * mat_B[8][27] +
                  mat_A[6][9] * mat_B[9][27] +
                  mat_A[6][10] * mat_B[10][27] +
                  mat_A[6][11] * mat_B[11][27] +
                  mat_A[6][12] * mat_B[12][27] +
                  mat_A[6][13] * mat_B[13][27] +
                  mat_A[6][14] * mat_B[14][27] +
                  mat_A[6][15] * mat_B[15][27] +
                  mat_A[6][16] * mat_B[16][27] +
                  mat_A[6][17] * mat_B[17][27] +
                  mat_A[6][18] * mat_B[18][27] +
                  mat_A[6][19] * mat_B[19][27] +
                  mat_A[6][20] * mat_B[20][27] +
                  mat_A[6][21] * mat_B[21][27] +
                  mat_A[6][22] * mat_B[22][27] +
                  mat_A[6][23] * mat_B[23][27] +
                  mat_A[6][24] * mat_B[24][27] +
                  mat_A[6][25] * mat_B[25][27] +
                  mat_A[6][26] * mat_B[26][27] +
                  mat_A[6][27] * mat_B[27][27] +
                  mat_A[6][28] * mat_B[28][27] +
                  mat_A[6][29] * mat_B[29][27] +
                  mat_A[6][30] * mat_B[30][27] +
                  mat_A[6][31] * mat_B[31][27];
    mat_C[6][28] <= 
                  mat_A[6][0] * mat_B[0][28] +
                  mat_A[6][1] * mat_B[1][28] +
                  mat_A[6][2] * mat_B[2][28] +
                  mat_A[6][3] * mat_B[3][28] +
                  mat_A[6][4] * mat_B[4][28] +
                  mat_A[6][5] * mat_B[5][28] +
                  mat_A[6][6] * mat_B[6][28] +
                  mat_A[6][7] * mat_B[7][28] +
                  mat_A[6][8] * mat_B[8][28] +
                  mat_A[6][9] * mat_B[9][28] +
                  mat_A[6][10] * mat_B[10][28] +
                  mat_A[6][11] * mat_B[11][28] +
                  mat_A[6][12] * mat_B[12][28] +
                  mat_A[6][13] * mat_B[13][28] +
                  mat_A[6][14] * mat_B[14][28] +
                  mat_A[6][15] * mat_B[15][28] +
                  mat_A[6][16] * mat_B[16][28] +
                  mat_A[6][17] * mat_B[17][28] +
                  mat_A[6][18] * mat_B[18][28] +
                  mat_A[6][19] * mat_B[19][28] +
                  mat_A[6][20] * mat_B[20][28] +
                  mat_A[6][21] * mat_B[21][28] +
                  mat_A[6][22] * mat_B[22][28] +
                  mat_A[6][23] * mat_B[23][28] +
                  mat_A[6][24] * mat_B[24][28] +
                  mat_A[6][25] * mat_B[25][28] +
                  mat_A[6][26] * mat_B[26][28] +
                  mat_A[6][27] * mat_B[27][28] +
                  mat_A[6][28] * mat_B[28][28] +
                  mat_A[6][29] * mat_B[29][28] +
                  mat_A[6][30] * mat_B[30][28] +
                  mat_A[6][31] * mat_B[31][28];
    mat_C[6][29] <= 
                  mat_A[6][0] * mat_B[0][29] +
                  mat_A[6][1] * mat_B[1][29] +
                  mat_A[6][2] * mat_B[2][29] +
                  mat_A[6][3] * mat_B[3][29] +
                  mat_A[6][4] * mat_B[4][29] +
                  mat_A[6][5] * mat_B[5][29] +
                  mat_A[6][6] * mat_B[6][29] +
                  mat_A[6][7] * mat_B[7][29] +
                  mat_A[6][8] * mat_B[8][29] +
                  mat_A[6][9] * mat_B[9][29] +
                  mat_A[6][10] * mat_B[10][29] +
                  mat_A[6][11] * mat_B[11][29] +
                  mat_A[6][12] * mat_B[12][29] +
                  mat_A[6][13] * mat_B[13][29] +
                  mat_A[6][14] * mat_B[14][29] +
                  mat_A[6][15] * mat_B[15][29] +
                  mat_A[6][16] * mat_B[16][29] +
                  mat_A[6][17] * mat_B[17][29] +
                  mat_A[6][18] * mat_B[18][29] +
                  mat_A[6][19] * mat_B[19][29] +
                  mat_A[6][20] * mat_B[20][29] +
                  mat_A[6][21] * mat_B[21][29] +
                  mat_A[6][22] * mat_B[22][29] +
                  mat_A[6][23] * mat_B[23][29] +
                  mat_A[6][24] * mat_B[24][29] +
                  mat_A[6][25] * mat_B[25][29] +
                  mat_A[6][26] * mat_B[26][29] +
                  mat_A[6][27] * mat_B[27][29] +
                  mat_A[6][28] * mat_B[28][29] +
                  mat_A[6][29] * mat_B[29][29] +
                  mat_A[6][30] * mat_B[30][29] +
                  mat_A[6][31] * mat_B[31][29];
    mat_C[6][30] <= 
                  mat_A[6][0] * mat_B[0][30] +
                  mat_A[6][1] * mat_B[1][30] +
                  mat_A[6][2] * mat_B[2][30] +
                  mat_A[6][3] * mat_B[3][30] +
                  mat_A[6][4] * mat_B[4][30] +
                  mat_A[6][5] * mat_B[5][30] +
                  mat_A[6][6] * mat_B[6][30] +
                  mat_A[6][7] * mat_B[7][30] +
                  mat_A[6][8] * mat_B[8][30] +
                  mat_A[6][9] * mat_B[9][30] +
                  mat_A[6][10] * mat_B[10][30] +
                  mat_A[6][11] * mat_B[11][30] +
                  mat_A[6][12] * mat_B[12][30] +
                  mat_A[6][13] * mat_B[13][30] +
                  mat_A[6][14] * mat_B[14][30] +
                  mat_A[6][15] * mat_B[15][30] +
                  mat_A[6][16] * mat_B[16][30] +
                  mat_A[6][17] * mat_B[17][30] +
                  mat_A[6][18] * mat_B[18][30] +
                  mat_A[6][19] * mat_B[19][30] +
                  mat_A[6][20] * mat_B[20][30] +
                  mat_A[6][21] * mat_B[21][30] +
                  mat_A[6][22] * mat_B[22][30] +
                  mat_A[6][23] * mat_B[23][30] +
                  mat_A[6][24] * mat_B[24][30] +
                  mat_A[6][25] * mat_B[25][30] +
                  mat_A[6][26] * mat_B[26][30] +
                  mat_A[6][27] * mat_B[27][30] +
                  mat_A[6][28] * mat_B[28][30] +
                  mat_A[6][29] * mat_B[29][30] +
                  mat_A[6][30] * mat_B[30][30] +
                  mat_A[6][31] * mat_B[31][30];
    mat_C[6][31] <= 
                  mat_A[6][0] * mat_B[0][31] +
                  mat_A[6][1] * mat_B[1][31] +
                  mat_A[6][2] * mat_B[2][31] +
                  mat_A[6][3] * mat_B[3][31] +
                  mat_A[6][4] * mat_B[4][31] +
                  mat_A[6][5] * mat_B[5][31] +
                  mat_A[6][6] * mat_B[6][31] +
                  mat_A[6][7] * mat_B[7][31] +
                  mat_A[6][8] * mat_B[8][31] +
                  mat_A[6][9] * mat_B[9][31] +
                  mat_A[6][10] * mat_B[10][31] +
                  mat_A[6][11] * mat_B[11][31] +
                  mat_A[6][12] * mat_B[12][31] +
                  mat_A[6][13] * mat_B[13][31] +
                  mat_A[6][14] * mat_B[14][31] +
                  mat_A[6][15] * mat_B[15][31] +
                  mat_A[6][16] * mat_B[16][31] +
                  mat_A[6][17] * mat_B[17][31] +
                  mat_A[6][18] * mat_B[18][31] +
                  mat_A[6][19] * mat_B[19][31] +
                  mat_A[6][20] * mat_B[20][31] +
                  mat_A[6][21] * mat_B[21][31] +
                  mat_A[6][22] * mat_B[22][31] +
                  mat_A[6][23] * mat_B[23][31] +
                  mat_A[6][24] * mat_B[24][31] +
                  mat_A[6][25] * mat_B[25][31] +
                  mat_A[6][26] * mat_B[26][31] +
                  mat_A[6][27] * mat_B[27][31] +
                  mat_A[6][28] * mat_B[28][31] +
                  mat_A[6][29] * mat_B[29][31] +
                  mat_A[6][30] * mat_B[30][31] +
                  mat_A[6][31] * mat_B[31][31];
    mat_C[7][0] <= 
                  mat_A[7][0] * mat_B[0][0] +
                  mat_A[7][1] * mat_B[1][0] +
                  mat_A[7][2] * mat_B[2][0] +
                  mat_A[7][3] * mat_B[3][0] +
                  mat_A[7][4] * mat_B[4][0] +
                  mat_A[7][5] * mat_B[5][0] +
                  mat_A[7][6] * mat_B[6][0] +
                  mat_A[7][7] * mat_B[7][0] +
                  mat_A[7][8] * mat_B[8][0] +
                  mat_A[7][9] * mat_B[9][0] +
                  mat_A[7][10] * mat_B[10][0] +
                  mat_A[7][11] * mat_B[11][0] +
                  mat_A[7][12] * mat_B[12][0] +
                  mat_A[7][13] * mat_B[13][0] +
                  mat_A[7][14] * mat_B[14][0] +
                  mat_A[7][15] * mat_B[15][0] +
                  mat_A[7][16] * mat_B[16][0] +
                  mat_A[7][17] * mat_B[17][0] +
                  mat_A[7][18] * mat_B[18][0] +
                  mat_A[7][19] * mat_B[19][0] +
                  mat_A[7][20] * mat_B[20][0] +
                  mat_A[7][21] * mat_B[21][0] +
                  mat_A[7][22] * mat_B[22][0] +
                  mat_A[7][23] * mat_B[23][0] +
                  mat_A[7][24] * mat_B[24][0] +
                  mat_A[7][25] * mat_B[25][0] +
                  mat_A[7][26] * mat_B[26][0] +
                  mat_A[7][27] * mat_B[27][0] +
                  mat_A[7][28] * mat_B[28][0] +
                  mat_A[7][29] * mat_B[29][0] +
                  mat_A[7][30] * mat_B[30][0] +
                  mat_A[7][31] * mat_B[31][0];
    mat_C[7][1] <= 
                  mat_A[7][0] * mat_B[0][1] +
                  mat_A[7][1] * mat_B[1][1] +
                  mat_A[7][2] * mat_B[2][1] +
                  mat_A[7][3] * mat_B[3][1] +
                  mat_A[7][4] * mat_B[4][1] +
                  mat_A[7][5] * mat_B[5][1] +
                  mat_A[7][6] * mat_B[6][1] +
                  mat_A[7][7] * mat_B[7][1] +
                  mat_A[7][8] * mat_B[8][1] +
                  mat_A[7][9] * mat_B[9][1] +
                  mat_A[7][10] * mat_B[10][1] +
                  mat_A[7][11] * mat_B[11][1] +
                  mat_A[7][12] * mat_B[12][1] +
                  mat_A[7][13] * mat_B[13][1] +
                  mat_A[7][14] * mat_B[14][1] +
                  mat_A[7][15] * mat_B[15][1] +
                  mat_A[7][16] * mat_B[16][1] +
                  mat_A[7][17] * mat_B[17][1] +
                  mat_A[7][18] * mat_B[18][1] +
                  mat_A[7][19] * mat_B[19][1] +
                  mat_A[7][20] * mat_B[20][1] +
                  mat_A[7][21] * mat_B[21][1] +
                  mat_A[7][22] * mat_B[22][1] +
                  mat_A[7][23] * mat_B[23][1] +
                  mat_A[7][24] * mat_B[24][1] +
                  mat_A[7][25] * mat_B[25][1] +
                  mat_A[7][26] * mat_B[26][1] +
                  mat_A[7][27] * mat_B[27][1] +
                  mat_A[7][28] * mat_B[28][1] +
                  mat_A[7][29] * mat_B[29][1] +
                  mat_A[7][30] * mat_B[30][1] +
                  mat_A[7][31] * mat_B[31][1];
    mat_C[7][2] <= 
                  mat_A[7][0] * mat_B[0][2] +
                  mat_A[7][1] * mat_B[1][2] +
                  mat_A[7][2] * mat_B[2][2] +
                  mat_A[7][3] * mat_B[3][2] +
                  mat_A[7][4] * mat_B[4][2] +
                  mat_A[7][5] * mat_B[5][2] +
                  mat_A[7][6] * mat_B[6][2] +
                  mat_A[7][7] * mat_B[7][2] +
                  mat_A[7][8] * mat_B[8][2] +
                  mat_A[7][9] * mat_B[9][2] +
                  mat_A[7][10] * mat_B[10][2] +
                  mat_A[7][11] * mat_B[11][2] +
                  mat_A[7][12] * mat_B[12][2] +
                  mat_A[7][13] * mat_B[13][2] +
                  mat_A[7][14] * mat_B[14][2] +
                  mat_A[7][15] * mat_B[15][2] +
                  mat_A[7][16] * mat_B[16][2] +
                  mat_A[7][17] * mat_B[17][2] +
                  mat_A[7][18] * mat_B[18][2] +
                  mat_A[7][19] * mat_B[19][2] +
                  mat_A[7][20] * mat_B[20][2] +
                  mat_A[7][21] * mat_B[21][2] +
                  mat_A[7][22] * mat_B[22][2] +
                  mat_A[7][23] * mat_B[23][2] +
                  mat_A[7][24] * mat_B[24][2] +
                  mat_A[7][25] * mat_B[25][2] +
                  mat_A[7][26] * mat_B[26][2] +
                  mat_A[7][27] * mat_B[27][2] +
                  mat_A[7][28] * mat_B[28][2] +
                  mat_A[7][29] * mat_B[29][2] +
                  mat_A[7][30] * mat_B[30][2] +
                  mat_A[7][31] * mat_B[31][2];
    mat_C[7][3] <= 
                  mat_A[7][0] * mat_B[0][3] +
                  mat_A[7][1] * mat_B[1][3] +
                  mat_A[7][2] * mat_B[2][3] +
                  mat_A[7][3] * mat_B[3][3] +
                  mat_A[7][4] * mat_B[4][3] +
                  mat_A[7][5] * mat_B[5][3] +
                  mat_A[7][6] * mat_B[6][3] +
                  mat_A[7][7] * mat_B[7][3] +
                  mat_A[7][8] * mat_B[8][3] +
                  mat_A[7][9] * mat_B[9][3] +
                  mat_A[7][10] * mat_B[10][3] +
                  mat_A[7][11] * mat_B[11][3] +
                  mat_A[7][12] * mat_B[12][3] +
                  mat_A[7][13] * mat_B[13][3] +
                  mat_A[7][14] * mat_B[14][3] +
                  mat_A[7][15] * mat_B[15][3] +
                  mat_A[7][16] * mat_B[16][3] +
                  mat_A[7][17] * mat_B[17][3] +
                  mat_A[7][18] * mat_B[18][3] +
                  mat_A[7][19] * mat_B[19][3] +
                  mat_A[7][20] * mat_B[20][3] +
                  mat_A[7][21] * mat_B[21][3] +
                  mat_A[7][22] * mat_B[22][3] +
                  mat_A[7][23] * mat_B[23][3] +
                  mat_A[7][24] * mat_B[24][3] +
                  mat_A[7][25] * mat_B[25][3] +
                  mat_A[7][26] * mat_B[26][3] +
                  mat_A[7][27] * mat_B[27][3] +
                  mat_A[7][28] * mat_B[28][3] +
                  mat_A[7][29] * mat_B[29][3] +
                  mat_A[7][30] * mat_B[30][3] +
                  mat_A[7][31] * mat_B[31][3];
    mat_C[7][4] <= 
                  mat_A[7][0] * mat_B[0][4] +
                  mat_A[7][1] * mat_B[1][4] +
                  mat_A[7][2] * mat_B[2][4] +
                  mat_A[7][3] * mat_B[3][4] +
                  mat_A[7][4] * mat_B[4][4] +
                  mat_A[7][5] * mat_B[5][4] +
                  mat_A[7][6] * mat_B[6][4] +
                  mat_A[7][7] * mat_B[7][4] +
                  mat_A[7][8] * mat_B[8][4] +
                  mat_A[7][9] * mat_B[9][4] +
                  mat_A[7][10] * mat_B[10][4] +
                  mat_A[7][11] * mat_B[11][4] +
                  mat_A[7][12] * mat_B[12][4] +
                  mat_A[7][13] * mat_B[13][4] +
                  mat_A[7][14] * mat_B[14][4] +
                  mat_A[7][15] * mat_B[15][4] +
                  mat_A[7][16] * mat_B[16][4] +
                  mat_A[7][17] * mat_B[17][4] +
                  mat_A[7][18] * mat_B[18][4] +
                  mat_A[7][19] * mat_B[19][4] +
                  mat_A[7][20] * mat_B[20][4] +
                  mat_A[7][21] * mat_B[21][4] +
                  mat_A[7][22] * mat_B[22][4] +
                  mat_A[7][23] * mat_B[23][4] +
                  mat_A[7][24] * mat_B[24][4] +
                  mat_A[7][25] * mat_B[25][4] +
                  mat_A[7][26] * mat_B[26][4] +
                  mat_A[7][27] * mat_B[27][4] +
                  mat_A[7][28] * mat_B[28][4] +
                  mat_A[7][29] * mat_B[29][4] +
                  mat_A[7][30] * mat_B[30][4] +
                  mat_A[7][31] * mat_B[31][4];
    mat_C[7][5] <= 
                  mat_A[7][0] * mat_B[0][5] +
                  mat_A[7][1] * mat_B[1][5] +
                  mat_A[7][2] * mat_B[2][5] +
                  mat_A[7][3] * mat_B[3][5] +
                  mat_A[7][4] * mat_B[4][5] +
                  mat_A[7][5] * mat_B[5][5] +
                  mat_A[7][6] * mat_B[6][5] +
                  mat_A[7][7] * mat_B[7][5] +
                  mat_A[7][8] * mat_B[8][5] +
                  mat_A[7][9] * mat_B[9][5] +
                  mat_A[7][10] * mat_B[10][5] +
                  mat_A[7][11] * mat_B[11][5] +
                  mat_A[7][12] * mat_B[12][5] +
                  mat_A[7][13] * mat_B[13][5] +
                  mat_A[7][14] * mat_B[14][5] +
                  mat_A[7][15] * mat_B[15][5] +
                  mat_A[7][16] * mat_B[16][5] +
                  mat_A[7][17] * mat_B[17][5] +
                  mat_A[7][18] * mat_B[18][5] +
                  mat_A[7][19] * mat_B[19][5] +
                  mat_A[7][20] * mat_B[20][5] +
                  mat_A[7][21] * mat_B[21][5] +
                  mat_A[7][22] * mat_B[22][5] +
                  mat_A[7][23] * mat_B[23][5] +
                  mat_A[7][24] * mat_B[24][5] +
                  mat_A[7][25] * mat_B[25][5] +
                  mat_A[7][26] * mat_B[26][5] +
                  mat_A[7][27] * mat_B[27][5] +
                  mat_A[7][28] * mat_B[28][5] +
                  mat_A[7][29] * mat_B[29][5] +
                  mat_A[7][30] * mat_B[30][5] +
                  mat_A[7][31] * mat_B[31][5];
    mat_C[7][6] <= 
                  mat_A[7][0] * mat_B[0][6] +
                  mat_A[7][1] * mat_B[1][6] +
                  mat_A[7][2] * mat_B[2][6] +
                  mat_A[7][3] * mat_B[3][6] +
                  mat_A[7][4] * mat_B[4][6] +
                  mat_A[7][5] * mat_B[5][6] +
                  mat_A[7][6] * mat_B[6][6] +
                  mat_A[7][7] * mat_B[7][6] +
                  mat_A[7][8] * mat_B[8][6] +
                  mat_A[7][9] * mat_B[9][6] +
                  mat_A[7][10] * mat_B[10][6] +
                  mat_A[7][11] * mat_B[11][6] +
                  mat_A[7][12] * mat_B[12][6] +
                  mat_A[7][13] * mat_B[13][6] +
                  mat_A[7][14] * mat_B[14][6] +
                  mat_A[7][15] * mat_B[15][6] +
                  mat_A[7][16] * mat_B[16][6] +
                  mat_A[7][17] * mat_B[17][6] +
                  mat_A[7][18] * mat_B[18][6] +
                  mat_A[7][19] * mat_B[19][6] +
                  mat_A[7][20] * mat_B[20][6] +
                  mat_A[7][21] * mat_B[21][6] +
                  mat_A[7][22] * mat_B[22][6] +
                  mat_A[7][23] * mat_B[23][6] +
                  mat_A[7][24] * mat_B[24][6] +
                  mat_A[7][25] * mat_B[25][6] +
                  mat_A[7][26] * mat_B[26][6] +
                  mat_A[7][27] * mat_B[27][6] +
                  mat_A[7][28] * mat_B[28][6] +
                  mat_A[7][29] * mat_B[29][6] +
                  mat_A[7][30] * mat_B[30][6] +
                  mat_A[7][31] * mat_B[31][6];
    mat_C[7][7] <= 
                  mat_A[7][0] * mat_B[0][7] +
                  mat_A[7][1] * mat_B[1][7] +
                  mat_A[7][2] * mat_B[2][7] +
                  mat_A[7][3] * mat_B[3][7] +
                  mat_A[7][4] * mat_B[4][7] +
                  mat_A[7][5] * mat_B[5][7] +
                  mat_A[7][6] * mat_B[6][7] +
                  mat_A[7][7] * mat_B[7][7] +
                  mat_A[7][8] * mat_B[8][7] +
                  mat_A[7][9] * mat_B[9][7] +
                  mat_A[7][10] * mat_B[10][7] +
                  mat_A[7][11] * mat_B[11][7] +
                  mat_A[7][12] * mat_B[12][7] +
                  mat_A[7][13] * mat_B[13][7] +
                  mat_A[7][14] * mat_B[14][7] +
                  mat_A[7][15] * mat_B[15][7] +
                  mat_A[7][16] * mat_B[16][7] +
                  mat_A[7][17] * mat_B[17][7] +
                  mat_A[7][18] * mat_B[18][7] +
                  mat_A[7][19] * mat_B[19][7] +
                  mat_A[7][20] * mat_B[20][7] +
                  mat_A[7][21] * mat_B[21][7] +
                  mat_A[7][22] * mat_B[22][7] +
                  mat_A[7][23] * mat_B[23][7] +
                  mat_A[7][24] * mat_B[24][7] +
                  mat_A[7][25] * mat_B[25][7] +
                  mat_A[7][26] * mat_B[26][7] +
                  mat_A[7][27] * mat_B[27][7] +
                  mat_A[7][28] * mat_B[28][7] +
                  mat_A[7][29] * mat_B[29][7] +
                  mat_A[7][30] * mat_B[30][7] +
                  mat_A[7][31] * mat_B[31][7];
    mat_C[7][8] <= 
                  mat_A[7][0] * mat_B[0][8] +
                  mat_A[7][1] * mat_B[1][8] +
                  mat_A[7][2] * mat_B[2][8] +
                  mat_A[7][3] * mat_B[3][8] +
                  mat_A[7][4] * mat_B[4][8] +
                  mat_A[7][5] * mat_B[5][8] +
                  mat_A[7][6] * mat_B[6][8] +
                  mat_A[7][7] * mat_B[7][8] +
                  mat_A[7][8] * mat_B[8][8] +
                  mat_A[7][9] * mat_B[9][8] +
                  mat_A[7][10] * mat_B[10][8] +
                  mat_A[7][11] * mat_B[11][8] +
                  mat_A[7][12] * mat_B[12][8] +
                  mat_A[7][13] * mat_B[13][8] +
                  mat_A[7][14] * mat_B[14][8] +
                  mat_A[7][15] * mat_B[15][8] +
                  mat_A[7][16] * mat_B[16][8] +
                  mat_A[7][17] * mat_B[17][8] +
                  mat_A[7][18] * mat_B[18][8] +
                  mat_A[7][19] * mat_B[19][8] +
                  mat_A[7][20] * mat_B[20][8] +
                  mat_A[7][21] * mat_B[21][8] +
                  mat_A[7][22] * mat_B[22][8] +
                  mat_A[7][23] * mat_B[23][8] +
                  mat_A[7][24] * mat_B[24][8] +
                  mat_A[7][25] * mat_B[25][8] +
                  mat_A[7][26] * mat_B[26][8] +
                  mat_A[7][27] * mat_B[27][8] +
                  mat_A[7][28] * mat_B[28][8] +
                  mat_A[7][29] * mat_B[29][8] +
                  mat_A[7][30] * mat_B[30][8] +
                  mat_A[7][31] * mat_B[31][8];
    mat_C[7][9] <= 
                  mat_A[7][0] * mat_B[0][9] +
                  mat_A[7][1] * mat_B[1][9] +
                  mat_A[7][2] * mat_B[2][9] +
                  mat_A[7][3] * mat_B[3][9] +
                  mat_A[7][4] * mat_B[4][9] +
                  mat_A[7][5] * mat_B[5][9] +
                  mat_A[7][6] * mat_B[6][9] +
                  mat_A[7][7] * mat_B[7][9] +
                  mat_A[7][8] * mat_B[8][9] +
                  mat_A[7][9] * mat_B[9][9] +
                  mat_A[7][10] * mat_B[10][9] +
                  mat_A[7][11] * mat_B[11][9] +
                  mat_A[7][12] * mat_B[12][9] +
                  mat_A[7][13] * mat_B[13][9] +
                  mat_A[7][14] * mat_B[14][9] +
                  mat_A[7][15] * mat_B[15][9] +
                  mat_A[7][16] * mat_B[16][9] +
                  mat_A[7][17] * mat_B[17][9] +
                  mat_A[7][18] * mat_B[18][9] +
                  mat_A[7][19] * mat_B[19][9] +
                  mat_A[7][20] * mat_B[20][9] +
                  mat_A[7][21] * mat_B[21][9] +
                  mat_A[7][22] * mat_B[22][9] +
                  mat_A[7][23] * mat_B[23][9] +
                  mat_A[7][24] * mat_B[24][9] +
                  mat_A[7][25] * mat_B[25][9] +
                  mat_A[7][26] * mat_B[26][9] +
                  mat_A[7][27] * mat_B[27][9] +
                  mat_A[7][28] * mat_B[28][9] +
                  mat_A[7][29] * mat_B[29][9] +
                  mat_A[7][30] * mat_B[30][9] +
                  mat_A[7][31] * mat_B[31][9];
    mat_C[7][10] <= 
                  mat_A[7][0] * mat_B[0][10] +
                  mat_A[7][1] * mat_B[1][10] +
                  mat_A[7][2] * mat_B[2][10] +
                  mat_A[7][3] * mat_B[3][10] +
                  mat_A[7][4] * mat_B[4][10] +
                  mat_A[7][5] * mat_B[5][10] +
                  mat_A[7][6] * mat_B[6][10] +
                  mat_A[7][7] * mat_B[7][10] +
                  mat_A[7][8] * mat_B[8][10] +
                  mat_A[7][9] * mat_B[9][10] +
                  mat_A[7][10] * mat_B[10][10] +
                  mat_A[7][11] * mat_B[11][10] +
                  mat_A[7][12] * mat_B[12][10] +
                  mat_A[7][13] * mat_B[13][10] +
                  mat_A[7][14] * mat_B[14][10] +
                  mat_A[7][15] * mat_B[15][10] +
                  mat_A[7][16] * mat_B[16][10] +
                  mat_A[7][17] * mat_B[17][10] +
                  mat_A[7][18] * mat_B[18][10] +
                  mat_A[7][19] * mat_B[19][10] +
                  mat_A[7][20] * mat_B[20][10] +
                  mat_A[7][21] * mat_B[21][10] +
                  mat_A[7][22] * mat_B[22][10] +
                  mat_A[7][23] * mat_B[23][10] +
                  mat_A[7][24] * mat_B[24][10] +
                  mat_A[7][25] * mat_B[25][10] +
                  mat_A[7][26] * mat_B[26][10] +
                  mat_A[7][27] * mat_B[27][10] +
                  mat_A[7][28] * mat_B[28][10] +
                  mat_A[7][29] * mat_B[29][10] +
                  mat_A[7][30] * mat_B[30][10] +
                  mat_A[7][31] * mat_B[31][10];
    mat_C[7][11] <= 
                  mat_A[7][0] * mat_B[0][11] +
                  mat_A[7][1] * mat_B[1][11] +
                  mat_A[7][2] * mat_B[2][11] +
                  mat_A[7][3] * mat_B[3][11] +
                  mat_A[7][4] * mat_B[4][11] +
                  mat_A[7][5] * mat_B[5][11] +
                  mat_A[7][6] * mat_B[6][11] +
                  mat_A[7][7] * mat_B[7][11] +
                  mat_A[7][8] * mat_B[8][11] +
                  mat_A[7][9] * mat_B[9][11] +
                  mat_A[7][10] * mat_B[10][11] +
                  mat_A[7][11] * mat_B[11][11] +
                  mat_A[7][12] * mat_B[12][11] +
                  mat_A[7][13] * mat_B[13][11] +
                  mat_A[7][14] * mat_B[14][11] +
                  mat_A[7][15] * mat_B[15][11] +
                  mat_A[7][16] * mat_B[16][11] +
                  mat_A[7][17] * mat_B[17][11] +
                  mat_A[7][18] * mat_B[18][11] +
                  mat_A[7][19] * mat_B[19][11] +
                  mat_A[7][20] * mat_B[20][11] +
                  mat_A[7][21] * mat_B[21][11] +
                  mat_A[7][22] * mat_B[22][11] +
                  mat_A[7][23] * mat_B[23][11] +
                  mat_A[7][24] * mat_B[24][11] +
                  mat_A[7][25] * mat_B[25][11] +
                  mat_A[7][26] * mat_B[26][11] +
                  mat_A[7][27] * mat_B[27][11] +
                  mat_A[7][28] * mat_B[28][11] +
                  mat_A[7][29] * mat_B[29][11] +
                  mat_A[7][30] * mat_B[30][11] +
                  mat_A[7][31] * mat_B[31][11];
    mat_C[7][12] <= 
                  mat_A[7][0] * mat_B[0][12] +
                  mat_A[7][1] * mat_B[1][12] +
                  mat_A[7][2] * mat_B[2][12] +
                  mat_A[7][3] * mat_B[3][12] +
                  mat_A[7][4] * mat_B[4][12] +
                  mat_A[7][5] * mat_B[5][12] +
                  mat_A[7][6] * mat_B[6][12] +
                  mat_A[7][7] * mat_B[7][12] +
                  mat_A[7][8] * mat_B[8][12] +
                  mat_A[7][9] * mat_B[9][12] +
                  mat_A[7][10] * mat_B[10][12] +
                  mat_A[7][11] * mat_B[11][12] +
                  mat_A[7][12] * mat_B[12][12] +
                  mat_A[7][13] * mat_B[13][12] +
                  mat_A[7][14] * mat_B[14][12] +
                  mat_A[7][15] * mat_B[15][12] +
                  mat_A[7][16] * mat_B[16][12] +
                  mat_A[7][17] * mat_B[17][12] +
                  mat_A[7][18] * mat_B[18][12] +
                  mat_A[7][19] * mat_B[19][12] +
                  mat_A[7][20] * mat_B[20][12] +
                  mat_A[7][21] * mat_B[21][12] +
                  mat_A[7][22] * mat_B[22][12] +
                  mat_A[7][23] * mat_B[23][12] +
                  mat_A[7][24] * mat_B[24][12] +
                  mat_A[7][25] * mat_B[25][12] +
                  mat_A[7][26] * mat_B[26][12] +
                  mat_A[7][27] * mat_B[27][12] +
                  mat_A[7][28] * mat_B[28][12] +
                  mat_A[7][29] * mat_B[29][12] +
                  mat_A[7][30] * mat_B[30][12] +
                  mat_A[7][31] * mat_B[31][12];
    mat_C[7][13] <= 
                  mat_A[7][0] * mat_B[0][13] +
                  mat_A[7][1] * mat_B[1][13] +
                  mat_A[7][2] * mat_B[2][13] +
                  mat_A[7][3] * mat_B[3][13] +
                  mat_A[7][4] * mat_B[4][13] +
                  mat_A[7][5] * mat_B[5][13] +
                  mat_A[7][6] * mat_B[6][13] +
                  mat_A[7][7] * mat_B[7][13] +
                  mat_A[7][8] * mat_B[8][13] +
                  mat_A[7][9] * mat_B[9][13] +
                  mat_A[7][10] * mat_B[10][13] +
                  mat_A[7][11] * mat_B[11][13] +
                  mat_A[7][12] * mat_B[12][13] +
                  mat_A[7][13] * mat_B[13][13] +
                  mat_A[7][14] * mat_B[14][13] +
                  mat_A[7][15] * mat_B[15][13] +
                  mat_A[7][16] * mat_B[16][13] +
                  mat_A[7][17] * mat_B[17][13] +
                  mat_A[7][18] * mat_B[18][13] +
                  mat_A[7][19] * mat_B[19][13] +
                  mat_A[7][20] * mat_B[20][13] +
                  mat_A[7][21] * mat_B[21][13] +
                  mat_A[7][22] * mat_B[22][13] +
                  mat_A[7][23] * mat_B[23][13] +
                  mat_A[7][24] * mat_B[24][13] +
                  mat_A[7][25] * mat_B[25][13] +
                  mat_A[7][26] * mat_B[26][13] +
                  mat_A[7][27] * mat_B[27][13] +
                  mat_A[7][28] * mat_B[28][13] +
                  mat_A[7][29] * mat_B[29][13] +
                  mat_A[7][30] * mat_B[30][13] +
                  mat_A[7][31] * mat_B[31][13];
    mat_C[7][14] <= 
                  mat_A[7][0] * mat_B[0][14] +
                  mat_A[7][1] * mat_B[1][14] +
                  mat_A[7][2] * mat_B[2][14] +
                  mat_A[7][3] * mat_B[3][14] +
                  mat_A[7][4] * mat_B[4][14] +
                  mat_A[7][5] * mat_B[5][14] +
                  mat_A[7][6] * mat_B[6][14] +
                  mat_A[7][7] * mat_B[7][14] +
                  mat_A[7][8] * mat_B[8][14] +
                  mat_A[7][9] * mat_B[9][14] +
                  mat_A[7][10] * mat_B[10][14] +
                  mat_A[7][11] * mat_B[11][14] +
                  mat_A[7][12] * mat_B[12][14] +
                  mat_A[7][13] * mat_B[13][14] +
                  mat_A[7][14] * mat_B[14][14] +
                  mat_A[7][15] * mat_B[15][14] +
                  mat_A[7][16] * mat_B[16][14] +
                  mat_A[7][17] * mat_B[17][14] +
                  mat_A[7][18] * mat_B[18][14] +
                  mat_A[7][19] * mat_B[19][14] +
                  mat_A[7][20] * mat_B[20][14] +
                  mat_A[7][21] * mat_B[21][14] +
                  mat_A[7][22] * mat_B[22][14] +
                  mat_A[7][23] * mat_B[23][14] +
                  mat_A[7][24] * mat_B[24][14] +
                  mat_A[7][25] * mat_B[25][14] +
                  mat_A[7][26] * mat_B[26][14] +
                  mat_A[7][27] * mat_B[27][14] +
                  mat_A[7][28] * mat_B[28][14] +
                  mat_A[7][29] * mat_B[29][14] +
                  mat_A[7][30] * mat_B[30][14] +
                  mat_A[7][31] * mat_B[31][14];
    mat_C[7][15] <= 
                  mat_A[7][0] * mat_B[0][15] +
                  mat_A[7][1] * mat_B[1][15] +
                  mat_A[7][2] * mat_B[2][15] +
                  mat_A[7][3] * mat_B[3][15] +
                  mat_A[7][4] * mat_B[4][15] +
                  mat_A[7][5] * mat_B[5][15] +
                  mat_A[7][6] * mat_B[6][15] +
                  mat_A[7][7] * mat_B[7][15] +
                  mat_A[7][8] * mat_B[8][15] +
                  mat_A[7][9] * mat_B[9][15] +
                  mat_A[7][10] * mat_B[10][15] +
                  mat_A[7][11] * mat_B[11][15] +
                  mat_A[7][12] * mat_B[12][15] +
                  mat_A[7][13] * mat_B[13][15] +
                  mat_A[7][14] * mat_B[14][15] +
                  mat_A[7][15] * mat_B[15][15] +
                  mat_A[7][16] * mat_B[16][15] +
                  mat_A[7][17] * mat_B[17][15] +
                  mat_A[7][18] * mat_B[18][15] +
                  mat_A[7][19] * mat_B[19][15] +
                  mat_A[7][20] * mat_B[20][15] +
                  mat_A[7][21] * mat_B[21][15] +
                  mat_A[7][22] * mat_B[22][15] +
                  mat_A[7][23] * mat_B[23][15] +
                  mat_A[7][24] * mat_B[24][15] +
                  mat_A[7][25] * mat_B[25][15] +
                  mat_A[7][26] * mat_B[26][15] +
                  mat_A[7][27] * mat_B[27][15] +
                  mat_A[7][28] * mat_B[28][15] +
                  mat_A[7][29] * mat_B[29][15] +
                  mat_A[7][30] * mat_B[30][15] +
                  mat_A[7][31] * mat_B[31][15];
    mat_C[7][16] <= 
                  mat_A[7][0] * mat_B[0][16] +
                  mat_A[7][1] * mat_B[1][16] +
                  mat_A[7][2] * mat_B[2][16] +
                  mat_A[7][3] * mat_B[3][16] +
                  mat_A[7][4] * mat_B[4][16] +
                  mat_A[7][5] * mat_B[5][16] +
                  mat_A[7][6] * mat_B[6][16] +
                  mat_A[7][7] * mat_B[7][16] +
                  mat_A[7][8] * mat_B[8][16] +
                  mat_A[7][9] * mat_B[9][16] +
                  mat_A[7][10] * mat_B[10][16] +
                  mat_A[7][11] * mat_B[11][16] +
                  mat_A[7][12] * mat_B[12][16] +
                  mat_A[7][13] * mat_B[13][16] +
                  mat_A[7][14] * mat_B[14][16] +
                  mat_A[7][15] * mat_B[15][16] +
                  mat_A[7][16] * mat_B[16][16] +
                  mat_A[7][17] * mat_B[17][16] +
                  mat_A[7][18] * mat_B[18][16] +
                  mat_A[7][19] * mat_B[19][16] +
                  mat_A[7][20] * mat_B[20][16] +
                  mat_A[7][21] * mat_B[21][16] +
                  mat_A[7][22] * mat_B[22][16] +
                  mat_A[7][23] * mat_B[23][16] +
                  mat_A[7][24] * mat_B[24][16] +
                  mat_A[7][25] * mat_B[25][16] +
                  mat_A[7][26] * mat_B[26][16] +
                  mat_A[7][27] * mat_B[27][16] +
                  mat_A[7][28] * mat_B[28][16] +
                  mat_A[7][29] * mat_B[29][16] +
                  mat_A[7][30] * mat_B[30][16] +
                  mat_A[7][31] * mat_B[31][16];
    mat_C[7][17] <= 
                  mat_A[7][0] * mat_B[0][17] +
                  mat_A[7][1] * mat_B[1][17] +
                  mat_A[7][2] * mat_B[2][17] +
                  mat_A[7][3] * mat_B[3][17] +
                  mat_A[7][4] * mat_B[4][17] +
                  mat_A[7][5] * mat_B[5][17] +
                  mat_A[7][6] * mat_B[6][17] +
                  mat_A[7][7] * mat_B[7][17] +
                  mat_A[7][8] * mat_B[8][17] +
                  mat_A[7][9] * mat_B[9][17] +
                  mat_A[7][10] * mat_B[10][17] +
                  mat_A[7][11] * mat_B[11][17] +
                  mat_A[7][12] * mat_B[12][17] +
                  mat_A[7][13] * mat_B[13][17] +
                  mat_A[7][14] * mat_B[14][17] +
                  mat_A[7][15] * mat_B[15][17] +
                  mat_A[7][16] * mat_B[16][17] +
                  mat_A[7][17] * mat_B[17][17] +
                  mat_A[7][18] * mat_B[18][17] +
                  mat_A[7][19] * mat_B[19][17] +
                  mat_A[7][20] * mat_B[20][17] +
                  mat_A[7][21] * mat_B[21][17] +
                  mat_A[7][22] * mat_B[22][17] +
                  mat_A[7][23] * mat_B[23][17] +
                  mat_A[7][24] * mat_B[24][17] +
                  mat_A[7][25] * mat_B[25][17] +
                  mat_A[7][26] * mat_B[26][17] +
                  mat_A[7][27] * mat_B[27][17] +
                  mat_A[7][28] * mat_B[28][17] +
                  mat_A[7][29] * mat_B[29][17] +
                  mat_A[7][30] * mat_B[30][17] +
                  mat_A[7][31] * mat_B[31][17];
    mat_C[7][18] <= 
                  mat_A[7][0] * mat_B[0][18] +
                  mat_A[7][1] * mat_B[1][18] +
                  mat_A[7][2] * mat_B[2][18] +
                  mat_A[7][3] * mat_B[3][18] +
                  mat_A[7][4] * mat_B[4][18] +
                  mat_A[7][5] * mat_B[5][18] +
                  mat_A[7][6] * mat_B[6][18] +
                  mat_A[7][7] * mat_B[7][18] +
                  mat_A[7][8] * mat_B[8][18] +
                  mat_A[7][9] * mat_B[9][18] +
                  mat_A[7][10] * mat_B[10][18] +
                  mat_A[7][11] * mat_B[11][18] +
                  mat_A[7][12] * mat_B[12][18] +
                  mat_A[7][13] * mat_B[13][18] +
                  mat_A[7][14] * mat_B[14][18] +
                  mat_A[7][15] * mat_B[15][18] +
                  mat_A[7][16] * mat_B[16][18] +
                  mat_A[7][17] * mat_B[17][18] +
                  mat_A[7][18] * mat_B[18][18] +
                  mat_A[7][19] * mat_B[19][18] +
                  mat_A[7][20] * mat_B[20][18] +
                  mat_A[7][21] * mat_B[21][18] +
                  mat_A[7][22] * mat_B[22][18] +
                  mat_A[7][23] * mat_B[23][18] +
                  mat_A[7][24] * mat_B[24][18] +
                  mat_A[7][25] * mat_B[25][18] +
                  mat_A[7][26] * mat_B[26][18] +
                  mat_A[7][27] * mat_B[27][18] +
                  mat_A[7][28] * mat_B[28][18] +
                  mat_A[7][29] * mat_B[29][18] +
                  mat_A[7][30] * mat_B[30][18] +
                  mat_A[7][31] * mat_B[31][18];
    mat_C[7][19] <= 
                  mat_A[7][0] * mat_B[0][19] +
                  mat_A[7][1] * mat_B[1][19] +
                  mat_A[7][2] * mat_B[2][19] +
                  mat_A[7][3] * mat_B[3][19] +
                  mat_A[7][4] * mat_B[4][19] +
                  mat_A[7][5] * mat_B[5][19] +
                  mat_A[7][6] * mat_B[6][19] +
                  mat_A[7][7] * mat_B[7][19] +
                  mat_A[7][8] * mat_B[8][19] +
                  mat_A[7][9] * mat_B[9][19] +
                  mat_A[7][10] * mat_B[10][19] +
                  mat_A[7][11] * mat_B[11][19] +
                  mat_A[7][12] * mat_B[12][19] +
                  mat_A[7][13] * mat_B[13][19] +
                  mat_A[7][14] * mat_B[14][19] +
                  mat_A[7][15] * mat_B[15][19] +
                  mat_A[7][16] * mat_B[16][19] +
                  mat_A[7][17] * mat_B[17][19] +
                  mat_A[7][18] * mat_B[18][19] +
                  mat_A[7][19] * mat_B[19][19] +
                  mat_A[7][20] * mat_B[20][19] +
                  mat_A[7][21] * mat_B[21][19] +
                  mat_A[7][22] * mat_B[22][19] +
                  mat_A[7][23] * mat_B[23][19] +
                  mat_A[7][24] * mat_B[24][19] +
                  mat_A[7][25] * mat_B[25][19] +
                  mat_A[7][26] * mat_B[26][19] +
                  mat_A[7][27] * mat_B[27][19] +
                  mat_A[7][28] * mat_B[28][19] +
                  mat_A[7][29] * mat_B[29][19] +
                  mat_A[7][30] * mat_B[30][19] +
                  mat_A[7][31] * mat_B[31][19];
    mat_C[7][20] <= 
                  mat_A[7][0] * mat_B[0][20] +
                  mat_A[7][1] * mat_B[1][20] +
                  mat_A[7][2] * mat_B[2][20] +
                  mat_A[7][3] * mat_B[3][20] +
                  mat_A[7][4] * mat_B[4][20] +
                  mat_A[7][5] * mat_B[5][20] +
                  mat_A[7][6] * mat_B[6][20] +
                  mat_A[7][7] * mat_B[7][20] +
                  mat_A[7][8] * mat_B[8][20] +
                  mat_A[7][9] * mat_B[9][20] +
                  mat_A[7][10] * mat_B[10][20] +
                  mat_A[7][11] * mat_B[11][20] +
                  mat_A[7][12] * mat_B[12][20] +
                  mat_A[7][13] * mat_B[13][20] +
                  mat_A[7][14] * mat_B[14][20] +
                  mat_A[7][15] * mat_B[15][20] +
                  mat_A[7][16] * mat_B[16][20] +
                  mat_A[7][17] * mat_B[17][20] +
                  mat_A[7][18] * mat_B[18][20] +
                  mat_A[7][19] * mat_B[19][20] +
                  mat_A[7][20] * mat_B[20][20] +
                  mat_A[7][21] * mat_B[21][20] +
                  mat_A[7][22] * mat_B[22][20] +
                  mat_A[7][23] * mat_B[23][20] +
                  mat_A[7][24] * mat_B[24][20] +
                  mat_A[7][25] * mat_B[25][20] +
                  mat_A[7][26] * mat_B[26][20] +
                  mat_A[7][27] * mat_B[27][20] +
                  mat_A[7][28] * mat_B[28][20] +
                  mat_A[7][29] * mat_B[29][20] +
                  mat_A[7][30] * mat_B[30][20] +
                  mat_A[7][31] * mat_B[31][20];
    mat_C[7][21] <= 
                  mat_A[7][0] * mat_B[0][21] +
                  mat_A[7][1] * mat_B[1][21] +
                  mat_A[7][2] * mat_B[2][21] +
                  mat_A[7][3] * mat_B[3][21] +
                  mat_A[7][4] * mat_B[4][21] +
                  mat_A[7][5] * mat_B[5][21] +
                  mat_A[7][6] * mat_B[6][21] +
                  mat_A[7][7] * mat_B[7][21] +
                  mat_A[7][8] * mat_B[8][21] +
                  mat_A[7][9] * mat_B[9][21] +
                  mat_A[7][10] * mat_B[10][21] +
                  mat_A[7][11] * mat_B[11][21] +
                  mat_A[7][12] * mat_B[12][21] +
                  mat_A[7][13] * mat_B[13][21] +
                  mat_A[7][14] * mat_B[14][21] +
                  mat_A[7][15] * mat_B[15][21] +
                  mat_A[7][16] * mat_B[16][21] +
                  mat_A[7][17] * mat_B[17][21] +
                  mat_A[7][18] * mat_B[18][21] +
                  mat_A[7][19] * mat_B[19][21] +
                  mat_A[7][20] * mat_B[20][21] +
                  mat_A[7][21] * mat_B[21][21] +
                  mat_A[7][22] * mat_B[22][21] +
                  mat_A[7][23] * mat_B[23][21] +
                  mat_A[7][24] * mat_B[24][21] +
                  mat_A[7][25] * mat_B[25][21] +
                  mat_A[7][26] * mat_B[26][21] +
                  mat_A[7][27] * mat_B[27][21] +
                  mat_A[7][28] * mat_B[28][21] +
                  mat_A[7][29] * mat_B[29][21] +
                  mat_A[7][30] * mat_B[30][21] +
                  mat_A[7][31] * mat_B[31][21];
    mat_C[7][22] <= 
                  mat_A[7][0] * mat_B[0][22] +
                  mat_A[7][1] * mat_B[1][22] +
                  mat_A[7][2] * mat_B[2][22] +
                  mat_A[7][3] * mat_B[3][22] +
                  mat_A[7][4] * mat_B[4][22] +
                  mat_A[7][5] * mat_B[5][22] +
                  mat_A[7][6] * mat_B[6][22] +
                  mat_A[7][7] * mat_B[7][22] +
                  mat_A[7][8] * mat_B[8][22] +
                  mat_A[7][9] * mat_B[9][22] +
                  mat_A[7][10] * mat_B[10][22] +
                  mat_A[7][11] * mat_B[11][22] +
                  mat_A[7][12] * mat_B[12][22] +
                  mat_A[7][13] * mat_B[13][22] +
                  mat_A[7][14] * mat_B[14][22] +
                  mat_A[7][15] * mat_B[15][22] +
                  mat_A[7][16] * mat_B[16][22] +
                  mat_A[7][17] * mat_B[17][22] +
                  mat_A[7][18] * mat_B[18][22] +
                  mat_A[7][19] * mat_B[19][22] +
                  mat_A[7][20] * mat_B[20][22] +
                  mat_A[7][21] * mat_B[21][22] +
                  mat_A[7][22] * mat_B[22][22] +
                  mat_A[7][23] * mat_B[23][22] +
                  mat_A[7][24] * mat_B[24][22] +
                  mat_A[7][25] * mat_B[25][22] +
                  mat_A[7][26] * mat_B[26][22] +
                  mat_A[7][27] * mat_B[27][22] +
                  mat_A[7][28] * mat_B[28][22] +
                  mat_A[7][29] * mat_B[29][22] +
                  mat_A[7][30] * mat_B[30][22] +
                  mat_A[7][31] * mat_B[31][22];
    mat_C[7][23] <= 
                  mat_A[7][0] * mat_B[0][23] +
                  mat_A[7][1] * mat_B[1][23] +
                  mat_A[7][2] * mat_B[2][23] +
                  mat_A[7][3] * mat_B[3][23] +
                  mat_A[7][4] * mat_B[4][23] +
                  mat_A[7][5] * mat_B[5][23] +
                  mat_A[7][6] * mat_B[6][23] +
                  mat_A[7][7] * mat_B[7][23] +
                  mat_A[7][8] * mat_B[8][23] +
                  mat_A[7][9] * mat_B[9][23] +
                  mat_A[7][10] * mat_B[10][23] +
                  mat_A[7][11] * mat_B[11][23] +
                  mat_A[7][12] * mat_B[12][23] +
                  mat_A[7][13] * mat_B[13][23] +
                  mat_A[7][14] * mat_B[14][23] +
                  mat_A[7][15] * mat_B[15][23] +
                  mat_A[7][16] * mat_B[16][23] +
                  mat_A[7][17] * mat_B[17][23] +
                  mat_A[7][18] * mat_B[18][23] +
                  mat_A[7][19] * mat_B[19][23] +
                  mat_A[7][20] * mat_B[20][23] +
                  mat_A[7][21] * mat_B[21][23] +
                  mat_A[7][22] * mat_B[22][23] +
                  mat_A[7][23] * mat_B[23][23] +
                  mat_A[7][24] * mat_B[24][23] +
                  mat_A[7][25] * mat_B[25][23] +
                  mat_A[7][26] * mat_B[26][23] +
                  mat_A[7][27] * mat_B[27][23] +
                  mat_A[7][28] * mat_B[28][23] +
                  mat_A[7][29] * mat_B[29][23] +
                  mat_A[7][30] * mat_B[30][23] +
                  mat_A[7][31] * mat_B[31][23];
    mat_C[7][24] <= 
                  mat_A[7][0] * mat_B[0][24] +
                  mat_A[7][1] * mat_B[1][24] +
                  mat_A[7][2] * mat_B[2][24] +
                  mat_A[7][3] * mat_B[3][24] +
                  mat_A[7][4] * mat_B[4][24] +
                  mat_A[7][5] * mat_B[5][24] +
                  mat_A[7][6] * mat_B[6][24] +
                  mat_A[7][7] * mat_B[7][24] +
                  mat_A[7][8] * mat_B[8][24] +
                  mat_A[7][9] * mat_B[9][24] +
                  mat_A[7][10] * mat_B[10][24] +
                  mat_A[7][11] * mat_B[11][24] +
                  mat_A[7][12] * mat_B[12][24] +
                  mat_A[7][13] * mat_B[13][24] +
                  mat_A[7][14] * mat_B[14][24] +
                  mat_A[7][15] * mat_B[15][24] +
                  mat_A[7][16] * mat_B[16][24] +
                  mat_A[7][17] * mat_B[17][24] +
                  mat_A[7][18] * mat_B[18][24] +
                  mat_A[7][19] * mat_B[19][24] +
                  mat_A[7][20] * mat_B[20][24] +
                  mat_A[7][21] * mat_B[21][24] +
                  mat_A[7][22] * mat_B[22][24] +
                  mat_A[7][23] * mat_B[23][24] +
                  mat_A[7][24] * mat_B[24][24] +
                  mat_A[7][25] * mat_B[25][24] +
                  mat_A[7][26] * mat_B[26][24] +
                  mat_A[7][27] * mat_B[27][24] +
                  mat_A[7][28] * mat_B[28][24] +
                  mat_A[7][29] * mat_B[29][24] +
                  mat_A[7][30] * mat_B[30][24] +
                  mat_A[7][31] * mat_B[31][24];
    mat_C[7][25] <= 
                  mat_A[7][0] * mat_B[0][25] +
                  mat_A[7][1] * mat_B[1][25] +
                  mat_A[7][2] * mat_B[2][25] +
                  mat_A[7][3] * mat_B[3][25] +
                  mat_A[7][4] * mat_B[4][25] +
                  mat_A[7][5] * mat_B[5][25] +
                  mat_A[7][6] * mat_B[6][25] +
                  mat_A[7][7] * mat_B[7][25] +
                  mat_A[7][8] * mat_B[8][25] +
                  mat_A[7][9] * mat_B[9][25] +
                  mat_A[7][10] * mat_B[10][25] +
                  mat_A[7][11] * mat_B[11][25] +
                  mat_A[7][12] * mat_B[12][25] +
                  mat_A[7][13] * mat_B[13][25] +
                  mat_A[7][14] * mat_B[14][25] +
                  mat_A[7][15] * mat_B[15][25] +
                  mat_A[7][16] * mat_B[16][25] +
                  mat_A[7][17] * mat_B[17][25] +
                  mat_A[7][18] * mat_B[18][25] +
                  mat_A[7][19] * mat_B[19][25] +
                  mat_A[7][20] * mat_B[20][25] +
                  mat_A[7][21] * mat_B[21][25] +
                  mat_A[7][22] * mat_B[22][25] +
                  mat_A[7][23] * mat_B[23][25] +
                  mat_A[7][24] * mat_B[24][25] +
                  mat_A[7][25] * mat_B[25][25] +
                  mat_A[7][26] * mat_B[26][25] +
                  mat_A[7][27] * mat_B[27][25] +
                  mat_A[7][28] * mat_B[28][25] +
                  mat_A[7][29] * mat_B[29][25] +
                  mat_A[7][30] * mat_B[30][25] +
                  mat_A[7][31] * mat_B[31][25];
    mat_C[7][26] <= 
                  mat_A[7][0] * mat_B[0][26] +
                  mat_A[7][1] * mat_B[1][26] +
                  mat_A[7][2] * mat_B[2][26] +
                  mat_A[7][3] * mat_B[3][26] +
                  mat_A[7][4] * mat_B[4][26] +
                  mat_A[7][5] * mat_B[5][26] +
                  mat_A[7][6] * mat_B[6][26] +
                  mat_A[7][7] * mat_B[7][26] +
                  mat_A[7][8] * mat_B[8][26] +
                  mat_A[7][9] * mat_B[9][26] +
                  mat_A[7][10] * mat_B[10][26] +
                  mat_A[7][11] * mat_B[11][26] +
                  mat_A[7][12] * mat_B[12][26] +
                  mat_A[7][13] * mat_B[13][26] +
                  mat_A[7][14] * mat_B[14][26] +
                  mat_A[7][15] * mat_B[15][26] +
                  mat_A[7][16] * mat_B[16][26] +
                  mat_A[7][17] * mat_B[17][26] +
                  mat_A[7][18] * mat_B[18][26] +
                  mat_A[7][19] * mat_B[19][26] +
                  mat_A[7][20] * mat_B[20][26] +
                  mat_A[7][21] * mat_B[21][26] +
                  mat_A[7][22] * mat_B[22][26] +
                  mat_A[7][23] * mat_B[23][26] +
                  mat_A[7][24] * mat_B[24][26] +
                  mat_A[7][25] * mat_B[25][26] +
                  mat_A[7][26] * mat_B[26][26] +
                  mat_A[7][27] * mat_B[27][26] +
                  mat_A[7][28] * mat_B[28][26] +
                  mat_A[7][29] * mat_B[29][26] +
                  mat_A[7][30] * mat_B[30][26] +
                  mat_A[7][31] * mat_B[31][26];
    mat_C[7][27] <= 
                  mat_A[7][0] * mat_B[0][27] +
                  mat_A[7][1] * mat_B[1][27] +
                  mat_A[7][2] * mat_B[2][27] +
                  mat_A[7][3] * mat_B[3][27] +
                  mat_A[7][4] * mat_B[4][27] +
                  mat_A[7][5] * mat_B[5][27] +
                  mat_A[7][6] * mat_B[6][27] +
                  mat_A[7][7] * mat_B[7][27] +
                  mat_A[7][8] * mat_B[8][27] +
                  mat_A[7][9] * mat_B[9][27] +
                  mat_A[7][10] * mat_B[10][27] +
                  mat_A[7][11] * mat_B[11][27] +
                  mat_A[7][12] * mat_B[12][27] +
                  mat_A[7][13] * mat_B[13][27] +
                  mat_A[7][14] * mat_B[14][27] +
                  mat_A[7][15] * mat_B[15][27] +
                  mat_A[7][16] * mat_B[16][27] +
                  mat_A[7][17] * mat_B[17][27] +
                  mat_A[7][18] * mat_B[18][27] +
                  mat_A[7][19] * mat_B[19][27] +
                  mat_A[7][20] * mat_B[20][27] +
                  mat_A[7][21] * mat_B[21][27] +
                  mat_A[7][22] * mat_B[22][27] +
                  mat_A[7][23] * mat_B[23][27] +
                  mat_A[7][24] * mat_B[24][27] +
                  mat_A[7][25] * mat_B[25][27] +
                  mat_A[7][26] * mat_B[26][27] +
                  mat_A[7][27] * mat_B[27][27] +
                  mat_A[7][28] * mat_B[28][27] +
                  mat_A[7][29] * mat_B[29][27] +
                  mat_A[7][30] * mat_B[30][27] +
                  mat_A[7][31] * mat_B[31][27];
    mat_C[7][28] <= 
                  mat_A[7][0] * mat_B[0][28] +
                  mat_A[7][1] * mat_B[1][28] +
                  mat_A[7][2] * mat_B[2][28] +
                  mat_A[7][3] * mat_B[3][28] +
                  mat_A[7][4] * mat_B[4][28] +
                  mat_A[7][5] * mat_B[5][28] +
                  mat_A[7][6] * mat_B[6][28] +
                  mat_A[7][7] * mat_B[7][28] +
                  mat_A[7][8] * mat_B[8][28] +
                  mat_A[7][9] * mat_B[9][28] +
                  mat_A[7][10] * mat_B[10][28] +
                  mat_A[7][11] * mat_B[11][28] +
                  mat_A[7][12] * mat_B[12][28] +
                  mat_A[7][13] * mat_B[13][28] +
                  mat_A[7][14] * mat_B[14][28] +
                  mat_A[7][15] * mat_B[15][28] +
                  mat_A[7][16] * mat_B[16][28] +
                  mat_A[7][17] * mat_B[17][28] +
                  mat_A[7][18] * mat_B[18][28] +
                  mat_A[7][19] * mat_B[19][28] +
                  mat_A[7][20] * mat_B[20][28] +
                  mat_A[7][21] * mat_B[21][28] +
                  mat_A[7][22] * mat_B[22][28] +
                  mat_A[7][23] * mat_B[23][28] +
                  mat_A[7][24] * mat_B[24][28] +
                  mat_A[7][25] * mat_B[25][28] +
                  mat_A[7][26] * mat_B[26][28] +
                  mat_A[7][27] * mat_B[27][28] +
                  mat_A[7][28] * mat_B[28][28] +
                  mat_A[7][29] * mat_B[29][28] +
                  mat_A[7][30] * mat_B[30][28] +
                  mat_A[7][31] * mat_B[31][28];
    mat_C[7][29] <= 
                  mat_A[7][0] * mat_B[0][29] +
                  mat_A[7][1] * mat_B[1][29] +
                  mat_A[7][2] * mat_B[2][29] +
                  mat_A[7][3] * mat_B[3][29] +
                  mat_A[7][4] * mat_B[4][29] +
                  mat_A[7][5] * mat_B[5][29] +
                  mat_A[7][6] * mat_B[6][29] +
                  mat_A[7][7] * mat_B[7][29] +
                  mat_A[7][8] * mat_B[8][29] +
                  mat_A[7][9] * mat_B[9][29] +
                  mat_A[7][10] * mat_B[10][29] +
                  mat_A[7][11] * mat_B[11][29] +
                  mat_A[7][12] * mat_B[12][29] +
                  mat_A[7][13] * mat_B[13][29] +
                  mat_A[7][14] * mat_B[14][29] +
                  mat_A[7][15] * mat_B[15][29] +
                  mat_A[7][16] * mat_B[16][29] +
                  mat_A[7][17] * mat_B[17][29] +
                  mat_A[7][18] * mat_B[18][29] +
                  mat_A[7][19] * mat_B[19][29] +
                  mat_A[7][20] * mat_B[20][29] +
                  mat_A[7][21] * mat_B[21][29] +
                  mat_A[7][22] * mat_B[22][29] +
                  mat_A[7][23] * mat_B[23][29] +
                  mat_A[7][24] * mat_B[24][29] +
                  mat_A[7][25] * mat_B[25][29] +
                  mat_A[7][26] * mat_B[26][29] +
                  mat_A[7][27] * mat_B[27][29] +
                  mat_A[7][28] * mat_B[28][29] +
                  mat_A[7][29] * mat_B[29][29] +
                  mat_A[7][30] * mat_B[30][29] +
                  mat_A[7][31] * mat_B[31][29];
    mat_C[7][30] <= 
                  mat_A[7][0] * mat_B[0][30] +
                  mat_A[7][1] * mat_B[1][30] +
                  mat_A[7][2] * mat_B[2][30] +
                  mat_A[7][3] * mat_B[3][30] +
                  mat_A[7][4] * mat_B[4][30] +
                  mat_A[7][5] * mat_B[5][30] +
                  mat_A[7][6] * mat_B[6][30] +
                  mat_A[7][7] * mat_B[7][30] +
                  mat_A[7][8] * mat_B[8][30] +
                  mat_A[7][9] * mat_B[9][30] +
                  mat_A[7][10] * mat_B[10][30] +
                  mat_A[7][11] * mat_B[11][30] +
                  mat_A[7][12] * mat_B[12][30] +
                  mat_A[7][13] * mat_B[13][30] +
                  mat_A[7][14] * mat_B[14][30] +
                  mat_A[7][15] * mat_B[15][30] +
                  mat_A[7][16] * mat_B[16][30] +
                  mat_A[7][17] * mat_B[17][30] +
                  mat_A[7][18] * mat_B[18][30] +
                  mat_A[7][19] * mat_B[19][30] +
                  mat_A[7][20] * mat_B[20][30] +
                  mat_A[7][21] * mat_B[21][30] +
                  mat_A[7][22] * mat_B[22][30] +
                  mat_A[7][23] * mat_B[23][30] +
                  mat_A[7][24] * mat_B[24][30] +
                  mat_A[7][25] * mat_B[25][30] +
                  mat_A[7][26] * mat_B[26][30] +
                  mat_A[7][27] * mat_B[27][30] +
                  mat_A[7][28] * mat_B[28][30] +
                  mat_A[7][29] * mat_B[29][30] +
                  mat_A[7][30] * mat_B[30][30] +
                  mat_A[7][31] * mat_B[31][30];
    mat_C[7][31] <= 
                  mat_A[7][0] * mat_B[0][31] +
                  mat_A[7][1] * mat_B[1][31] +
                  mat_A[7][2] * mat_B[2][31] +
                  mat_A[7][3] * mat_B[3][31] +
                  mat_A[7][4] * mat_B[4][31] +
                  mat_A[7][5] * mat_B[5][31] +
                  mat_A[7][6] * mat_B[6][31] +
                  mat_A[7][7] * mat_B[7][31] +
                  mat_A[7][8] * mat_B[8][31] +
                  mat_A[7][9] * mat_B[9][31] +
                  mat_A[7][10] * mat_B[10][31] +
                  mat_A[7][11] * mat_B[11][31] +
                  mat_A[7][12] * mat_B[12][31] +
                  mat_A[7][13] * mat_B[13][31] +
                  mat_A[7][14] * mat_B[14][31] +
                  mat_A[7][15] * mat_B[15][31] +
                  mat_A[7][16] * mat_B[16][31] +
                  mat_A[7][17] * mat_B[17][31] +
                  mat_A[7][18] * mat_B[18][31] +
                  mat_A[7][19] * mat_B[19][31] +
                  mat_A[7][20] * mat_B[20][31] +
                  mat_A[7][21] * mat_B[21][31] +
                  mat_A[7][22] * mat_B[22][31] +
                  mat_A[7][23] * mat_B[23][31] +
                  mat_A[7][24] * mat_B[24][31] +
                  mat_A[7][25] * mat_B[25][31] +
                  mat_A[7][26] * mat_B[26][31] +
                  mat_A[7][27] * mat_B[27][31] +
                  mat_A[7][28] * mat_B[28][31] +
                  mat_A[7][29] * mat_B[29][31] +
                  mat_A[7][30] * mat_B[30][31] +
                  mat_A[7][31] * mat_B[31][31];
    mat_C[8][0] <= 
                  mat_A[8][0] * mat_B[0][0] +
                  mat_A[8][1] * mat_B[1][0] +
                  mat_A[8][2] * mat_B[2][0] +
                  mat_A[8][3] * mat_B[3][0] +
                  mat_A[8][4] * mat_B[4][0] +
                  mat_A[8][5] * mat_B[5][0] +
                  mat_A[8][6] * mat_B[6][0] +
                  mat_A[8][7] * mat_B[7][0] +
                  mat_A[8][8] * mat_B[8][0] +
                  mat_A[8][9] * mat_B[9][0] +
                  mat_A[8][10] * mat_B[10][0] +
                  mat_A[8][11] * mat_B[11][0] +
                  mat_A[8][12] * mat_B[12][0] +
                  mat_A[8][13] * mat_B[13][0] +
                  mat_A[8][14] * mat_B[14][0] +
                  mat_A[8][15] * mat_B[15][0] +
                  mat_A[8][16] * mat_B[16][0] +
                  mat_A[8][17] * mat_B[17][0] +
                  mat_A[8][18] * mat_B[18][0] +
                  mat_A[8][19] * mat_B[19][0] +
                  mat_A[8][20] * mat_B[20][0] +
                  mat_A[8][21] * mat_B[21][0] +
                  mat_A[8][22] * mat_B[22][0] +
                  mat_A[8][23] * mat_B[23][0] +
                  mat_A[8][24] * mat_B[24][0] +
                  mat_A[8][25] * mat_B[25][0] +
                  mat_A[8][26] * mat_B[26][0] +
                  mat_A[8][27] * mat_B[27][0] +
                  mat_A[8][28] * mat_B[28][0] +
                  mat_A[8][29] * mat_B[29][0] +
                  mat_A[8][30] * mat_B[30][0] +
                  mat_A[8][31] * mat_B[31][0];
    mat_C[8][1] <= 
                  mat_A[8][0] * mat_B[0][1] +
                  mat_A[8][1] * mat_B[1][1] +
                  mat_A[8][2] * mat_B[2][1] +
                  mat_A[8][3] * mat_B[3][1] +
                  mat_A[8][4] * mat_B[4][1] +
                  mat_A[8][5] * mat_B[5][1] +
                  mat_A[8][6] * mat_B[6][1] +
                  mat_A[8][7] * mat_B[7][1] +
                  mat_A[8][8] * mat_B[8][1] +
                  mat_A[8][9] * mat_B[9][1] +
                  mat_A[8][10] * mat_B[10][1] +
                  mat_A[8][11] * mat_B[11][1] +
                  mat_A[8][12] * mat_B[12][1] +
                  mat_A[8][13] * mat_B[13][1] +
                  mat_A[8][14] * mat_B[14][1] +
                  mat_A[8][15] * mat_B[15][1] +
                  mat_A[8][16] * mat_B[16][1] +
                  mat_A[8][17] * mat_B[17][1] +
                  mat_A[8][18] * mat_B[18][1] +
                  mat_A[8][19] * mat_B[19][1] +
                  mat_A[8][20] * mat_B[20][1] +
                  mat_A[8][21] * mat_B[21][1] +
                  mat_A[8][22] * mat_B[22][1] +
                  mat_A[8][23] * mat_B[23][1] +
                  mat_A[8][24] * mat_B[24][1] +
                  mat_A[8][25] * mat_B[25][1] +
                  mat_A[8][26] * mat_B[26][1] +
                  mat_A[8][27] * mat_B[27][1] +
                  mat_A[8][28] * mat_B[28][1] +
                  mat_A[8][29] * mat_B[29][1] +
                  mat_A[8][30] * mat_B[30][1] +
                  mat_A[8][31] * mat_B[31][1];
    mat_C[8][2] <= 
                  mat_A[8][0] * mat_B[0][2] +
                  mat_A[8][1] * mat_B[1][2] +
                  mat_A[8][2] * mat_B[2][2] +
                  mat_A[8][3] * mat_B[3][2] +
                  mat_A[8][4] * mat_B[4][2] +
                  mat_A[8][5] * mat_B[5][2] +
                  mat_A[8][6] * mat_B[6][2] +
                  mat_A[8][7] * mat_B[7][2] +
                  mat_A[8][8] * mat_B[8][2] +
                  mat_A[8][9] * mat_B[9][2] +
                  mat_A[8][10] * mat_B[10][2] +
                  mat_A[8][11] * mat_B[11][2] +
                  mat_A[8][12] * mat_B[12][2] +
                  mat_A[8][13] * mat_B[13][2] +
                  mat_A[8][14] * mat_B[14][2] +
                  mat_A[8][15] * mat_B[15][2] +
                  mat_A[8][16] * mat_B[16][2] +
                  mat_A[8][17] * mat_B[17][2] +
                  mat_A[8][18] * mat_B[18][2] +
                  mat_A[8][19] * mat_B[19][2] +
                  mat_A[8][20] * mat_B[20][2] +
                  mat_A[8][21] * mat_B[21][2] +
                  mat_A[8][22] * mat_B[22][2] +
                  mat_A[8][23] * mat_B[23][2] +
                  mat_A[8][24] * mat_B[24][2] +
                  mat_A[8][25] * mat_B[25][2] +
                  mat_A[8][26] * mat_B[26][2] +
                  mat_A[8][27] * mat_B[27][2] +
                  mat_A[8][28] * mat_B[28][2] +
                  mat_A[8][29] * mat_B[29][2] +
                  mat_A[8][30] * mat_B[30][2] +
                  mat_A[8][31] * mat_B[31][2];
    mat_C[8][3] <= 
                  mat_A[8][0] * mat_B[0][3] +
                  mat_A[8][1] * mat_B[1][3] +
                  mat_A[8][2] * mat_B[2][3] +
                  mat_A[8][3] * mat_B[3][3] +
                  mat_A[8][4] * mat_B[4][3] +
                  mat_A[8][5] * mat_B[5][3] +
                  mat_A[8][6] * mat_B[6][3] +
                  mat_A[8][7] * mat_B[7][3] +
                  mat_A[8][8] * mat_B[8][3] +
                  mat_A[8][9] * mat_B[9][3] +
                  mat_A[8][10] * mat_B[10][3] +
                  mat_A[8][11] * mat_B[11][3] +
                  mat_A[8][12] * mat_B[12][3] +
                  mat_A[8][13] * mat_B[13][3] +
                  mat_A[8][14] * mat_B[14][3] +
                  mat_A[8][15] * mat_B[15][3] +
                  mat_A[8][16] * mat_B[16][3] +
                  mat_A[8][17] * mat_B[17][3] +
                  mat_A[8][18] * mat_B[18][3] +
                  mat_A[8][19] * mat_B[19][3] +
                  mat_A[8][20] * mat_B[20][3] +
                  mat_A[8][21] * mat_B[21][3] +
                  mat_A[8][22] * mat_B[22][3] +
                  mat_A[8][23] * mat_B[23][3] +
                  mat_A[8][24] * mat_B[24][3] +
                  mat_A[8][25] * mat_B[25][3] +
                  mat_A[8][26] * mat_B[26][3] +
                  mat_A[8][27] * mat_B[27][3] +
                  mat_A[8][28] * mat_B[28][3] +
                  mat_A[8][29] * mat_B[29][3] +
                  mat_A[8][30] * mat_B[30][3] +
                  mat_A[8][31] * mat_B[31][3];
    mat_C[8][4] <= 
                  mat_A[8][0] * mat_B[0][4] +
                  mat_A[8][1] * mat_B[1][4] +
                  mat_A[8][2] * mat_B[2][4] +
                  mat_A[8][3] * mat_B[3][4] +
                  mat_A[8][4] * mat_B[4][4] +
                  mat_A[8][5] * mat_B[5][4] +
                  mat_A[8][6] * mat_B[6][4] +
                  mat_A[8][7] * mat_B[7][4] +
                  mat_A[8][8] * mat_B[8][4] +
                  mat_A[8][9] * mat_B[9][4] +
                  mat_A[8][10] * mat_B[10][4] +
                  mat_A[8][11] * mat_B[11][4] +
                  mat_A[8][12] * mat_B[12][4] +
                  mat_A[8][13] * mat_B[13][4] +
                  mat_A[8][14] * mat_B[14][4] +
                  mat_A[8][15] * mat_B[15][4] +
                  mat_A[8][16] * mat_B[16][4] +
                  mat_A[8][17] * mat_B[17][4] +
                  mat_A[8][18] * mat_B[18][4] +
                  mat_A[8][19] * mat_B[19][4] +
                  mat_A[8][20] * mat_B[20][4] +
                  mat_A[8][21] * mat_B[21][4] +
                  mat_A[8][22] * mat_B[22][4] +
                  mat_A[8][23] * mat_B[23][4] +
                  mat_A[8][24] * mat_B[24][4] +
                  mat_A[8][25] * mat_B[25][4] +
                  mat_A[8][26] * mat_B[26][4] +
                  mat_A[8][27] * mat_B[27][4] +
                  mat_A[8][28] * mat_B[28][4] +
                  mat_A[8][29] * mat_B[29][4] +
                  mat_A[8][30] * mat_B[30][4] +
                  mat_A[8][31] * mat_B[31][4];
    mat_C[8][5] <= 
                  mat_A[8][0] * mat_B[0][5] +
                  mat_A[8][1] * mat_B[1][5] +
                  mat_A[8][2] * mat_B[2][5] +
                  mat_A[8][3] * mat_B[3][5] +
                  mat_A[8][4] * mat_B[4][5] +
                  mat_A[8][5] * mat_B[5][5] +
                  mat_A[8][6] * mat_B[6][5] +
                  mat_A[8][7] * mat_B[7][5] +
                  mat_A[8][8] * mat_B[8][5] +
                  mat_A[8][9] * mat_B[9][5] +
                  mat_A[8][10] * mat_B[10][5] +
                  mat_A[8][11] * mat_B[11][5] +
                  mat_A[8][12] * mat_B[12][5] +
                  mat_A[8][13] * mat_B[13][5] +
                  mat_A[8][14] * mat_B[14][5] +
                  mat_A[8][15] * mat_B[15][5] +
                  mat_A[8][16] * mat_B[16][5] +
                  mat_A[8][17] * mat_B[17][5] +
                  mat_A[8][18] * mat_B[18][5] +
                  mat_A[8][19] * mat_B[19][5] +
                  mat_A[8][20] * mat_B[20][5] +
                  mat_A[8][21] * mat_B[21][5] +
                  mat_A[8][22] * mat_B[22][5] +
                  mat_A[8][23] * mat_B[23][5] +
                  mat_A[8][24] * mat_B[24][5] +
                  mat_A[8][25] * mat_B[25][5] +
                  mat_A[8][26] * mat_B[26][5] +
                  mat_A[8][27] * mat_B[27][5] +
                  mat_A[8][28] * mat_B[28][5] +
                  mat_A[8][29] * mat_B[29][5] +
                  mat_A[8][30] * mat_B[30][5] +
                  mat_A[8][31] * mat_B[31][5];
    mat_C[8][6] <= 
                  mat_A[8][0] * mat_B[0][6] +
                  mat_A[8][1] * mat_B[1][6] +
                  mat_A[8][2] * mat_B[2][6] +
                  mat_A[8][3] * mat_B[3][6] +
                  mat_A[8][4] * mat_B[4][6] +
                  mat_A[8][5] * mat_B[5][6] +
                  mat_A[8][6] * mat_B[6][6] +
                  mat_A[8][7] * mat_B[7][6] +
                  mat_A[8][8] * mat_B[8][6] +
                  mat_A[8][9] * mat_B[9][6] +
                  mat_A[8][10] * mat_B[10][6] +
                  mat_A[8][11] * mat_B[11][6] +
                  mat_A[8][12] * mat_B[12][6] +
                  mat_A[8][13] * mat_B[13][6] +
                  mat_A[8][14] * mat_B[14][6] +
                  mat_A[8][15] * mat_B[15][6] +
                  mat_A[8][16] * mat_B[16][6] +
                  mat_A[8][17] * mat_B[17][6] +
                  mat_A[8][18] * mat_B[18][6] +
                  mat_A[8][19] * mat_B[19][6] +
                  mat_A[8][20] * mat_B[20][6] +
                  mat_A[8][21] * mat_B[21][6] +
                  mat_A[8][22] * mat_B[22][6] +
                  mat_A[8][23] * mat_B[23][6] +
                  mat_A[8][24] * mat_B[24][6] +
                  mat_A[8][25] * mat_B[25][6] +
                  mat_A[8][26] * mat_B[26][6] +
                  mat_A[8][27] * mat_B[27][6] +
                  mat_A[8][28] * mat_B[28][6] +
                  mat_A[8][29] * mat_B[29][6] +
                  mat_A[8][30] * mat_B[30][6] +
                  mat_A[8][31] * mat_B[31][6];
    mat_C[8][7] <= 
                  mat_A[8][0] * mat_B[0][7] +
                  mat_A[8][1] * mat_B[1][7] +
                  mat_A[8][2] * mat_B[2][7] +
                  mat_A[8][3] * mat_B[3][7] +
                  mat_A[8][4] * mat_B[4][7] +
                  mat_A[8][5] * mat_B[5][7] +
                  mat_A[8][6] * mat_B[6][7] +
                  mat_A[8][7] * mat_B[7][7] +
                  mat_A[8][8] * mat_B[8][7] +
                  mat_A[8][9] * mat_B[9][7] +
                  mat_A[8][10] * mat_B[10][7] +
                  mat_A[8][11] * mat_B[11][7] +
                  mat_A[8][12] * mat_B[12][7] +
                  mat_A[8][13] * mat_B[13][7] +
                  mat_A[8][14] * mat_B[14][7] +
                  mat_A[8][15] * mat_B[15][7] +
                  mat_A[8][16] * mat_B[16][7] +
                  mat_A[8][17] * mat_B[17][7] +
                  mat_A[8][18] * mat_B[18][7] +
                  mat_A[8][19] * mat_B[19][7] +
                  mat_A[8][20] * mat_B[20][7] +
                  mat_A[8][21] * mat_B[21][7] +
                  mat_A[8][22] * mat_B[22][7] +
                  mat_A[8][23] * mat_B[23][7] +
                  mat_A[8][24] * mat_B[24][7] +
                  mat_A[8][25] * mat_B[25][7] +
                  mat_A[8][26] * mat_B[26][7] +
                  mat_A[8][27] * mat_B[27][7] +
                  mat_A[8][28] * mat_B[28][7] +
                  mat_A[8][29] * mat_B[29][7] +
                  mat_A[8][30] * mat_B[30][7] +
                  mat_A[8][31] * mat_B[31][7];
    mat_C[8][8] <= 
                  mat_A[8][0] * mat_B[0][8] +
                  mat_A[8][1] * mat_B[1][8] +
                  mat_A[8][2] * mat_B[2][8] +
                  mat_A[8][3] * mat_B[3][8] +
                  mat_A[8][4] * mat_B[4][8] +
                  mat_A[8][5] * mat_B[5][8] +
                  mat_A[8][6] * mat_B[6][8] +
                  mat_A[8][7] * mat_B[7][8] +
                  mat_A[8][8] * mat_B[8][8] +
                  mat_A[8][9] * mat_B[9][8] +
                  mat_A[8][10] * mat_B[10][8] +
                  mat_A[8][11] * mat_B[11][8] +
                  mat_A[8][12] * mat_B[12][8] +
                  mat_A[8][13] * mat_B[13][8] +
                  mat_A[8][14] * mat_B[14][8] +
                  mat_A[8][15] * mat_B[15][8] +
                  mat_A[8][16] * mat_B[16][8] +
                  mat_A[8][17] * mat_B[17][8] +
                  mat_A[8][18] * mat_B[18][8] +
                  mat_A[8][19] * mat_B[19][8] +
                  mat_A[8][20] * mat_B[20][8] +
                  mat_A[8][21] * mat_B[21][8] +
                  mat_A[8][22] * mat_B[22][8] +
                  mat_A[8][23] * mat_B[23][8] +
                  mat_A[8][24] * mat_B[24][8] +
                  mat_A[8][25] * mat_B[25][8] +
                  mat_A[8][26] * mat_B[26][8] +
                  mat_A[8][27] * mat_B[27][8] +
                  mat_A[8][28] * mat_B[28][8] +
                  mat_A[8][29] * mat_B[29][8] +
                  mat_A[8][30] * mat_B[30][8] +
                  mat_A[8][31] * mat_B[31][8];
    mat_C[8][9] <= 
                  mat_A[8][0] * mat_B[0][9] +
                  mat_A[8][1] * mat_B[1][9] +
                  mat_A[8][2] * mat_B[2][9] +
                  mat_A[8][3] * mat_B[3][9] +
                  mat_A[8][4] * mat_B[4][9] +
                  mat_A[8][5] * mat_B[5][9] +
                  mat_A[8][6] * mat_B[6][9] +
                  mat_A[8][7] * mat_B[7][9] +
                  mat_A[8][8] * mat_B[8][9] +
                  mat_A[8][9] * mat_B[9][9] +
                  mat_A[8][10] * mat_B[10][9] +
                  mat_A[8][11] * mat_B[11][9] +
                  mat_A[8][12] * mat_B[12][9] +
                  mat_A[8][13] * mat_B[13][9] +
                  mat_A[8][14] * mat_B[14][9] +
                  mat_A[8][15] * mat_B[15][9] +
                  mat_A[8][16] * mat_B[16][9] +
                  mat_A[8][17] * mat_B[17][9] +
                  mat_A[8][18] * mat_B[18][9] +
                  mat_A[8][19] * mat_B[19][9] +
                  mat_A[8][20] * mat_B[20][9] +
                  mat_A[8][21] * mat_B[21][9] +
                  mat_A[8][22] * mat_B[22][9] +
                  mat_A[8][23] * mat_B[23][9] +
                  mat_A[8][24] * mat_B[24][9] +
                  mat_A[8][25] * mat_B[25][9] +
                  mat_A[8][26] * mat_B[26][9] +
                  mat_A[8][27] * mat_B[27][9] +
                  mat_A[8][28] * mat_B[28][9] +
                  mat_A[8][29] * mat_B[29][9] +
                  mat_A[8][30] * mat_B[30][9] +
                  mat_A[8][31] * mat_B[31][9];
    mat_C[8][10] <= 
                  mat_A[8][0] * mat_B[0][10] +
                  mat_A[8][1] * mat_B[1][10] +
                  mat_A[8][2] * mat_B[2][10] +
                  mat_A[8][3] * mat_B[3][10] +
                  mat_A[8][4] * mat_B[4][10] +
                  mat_A[8][5] * mat_B[5][10] +
                  mat_A[8][6] * mat_B[6][10] +
                  mat_A[8][7] * mat_B[7][10] +
                  mat_A[8][8] * mat_B[8][10] +
                  mat_A[8][9] * mat_B[9][10] +
                  mat_A[8][10] * mat_B[10][10] +
                  mat_A[8][11] * mat_B[11][10] +
                  mat_A[8][12] * mat_B[12][10] +
                  mat_A[8][13] * mat_B[13][10] +
                  mat_A[8][14] * mat_B[14][10] +
                  mat_A[8][15] * mat_B[15][10] +
                  mat_A[8][16] * mat_B[16][10] +
                  mat_A[8][17] * mat_B[17][10] +
                  mat_A[8][18] * mat_B[18][10] +
                  mat_A[8][19] * mat_B[19][10] +
                  mat_A[8][20] * mat_B[20][10] +
                  mat_A[8][21] * mat_B[21][10] +
                  mat_A[8][22] * mat_B[22][10] +
                  mat_A[8][23] * mat_B[23][10] +
                  mat_A[8][24] * mat_B[24][10] +
                  mat_A[8][25] * mat_B[25][10] +
                  mat_A[8][26] * mat_B[26][10] +
                  mat_A[8][27] * mat_B[27][10] +
                  mat_A[8][28] * mat_B[28][10] +
                  mat_A[8][29] * mat_B[29][10] +
                  mat_A[8][30] * mat_B[30][10] +
                  mat_A[8][31] * mat_B[31][10];
    mat_C[8][11] <= 
                  mat_A[8][0] * mat_B[0][11] +
                  mat_A[8][1] * mat_B[1][11] +
                  mat_A[8][2] * mat_B[2][11] +
                  mat_A[8][3] * mat_B[3][11] +
                  mat_A[8][4] * mat_B[4][11] +
                  mat_A[8][5] * mat_B[5][11] +
                  mat_A[8][6] * mat_B[6][11] +
                  mat_A[8][7] * mat_B[7][11] +
                  mat_A[8][8] * mat_B[8][11] +
                  mat_A[8][9] * mat_B[9][11] +
                  mat_A[8][10] * mat_B[10][11] +
                  mat_A[8][11] * mat_B[11][11] +
                  mat_A[8][12] * mat_B[12][11] +
                  mat_A[8][13] * mat_B[13][11] +
                  mat_A[8][14] * mat_B[14][11] +
                  mat_A[8][15] * mat_B[15][11] +
                  mat_A[8][16] * mat_B[16][11] +
                  mat_A[8][17] * mat_B[17][11] +
                  mat_A[8][18] * mat_B[18][11] +
                  mat_A[8][19] * mat_B[19][11] +
                  mat_A[8][20] * mat_B[20][11] +
                  mat_A[8][21] * mat_B[21][11] +
                  mat_A[8][22] * mat_B[22][11] +
                  mat_A[8][23] * mat_B[23][11] +
                  mat_A[8][24] * mat_B[24][11] +
                  mat_A[8][25] * mat_B[25][11] +
                  mat_A[8][26] * mat_B[26][11] +
                  mat_A[8][27] * mat_B[27][11] +
                  mat_A[8][28] * mat_B[28][11] +
                  mat_A[8][29] * mat_B[29][11] +
                  mat_A[8][30] * mat_B[30][11] +
                  mat_A[8][31] * mat_B[31][11];
    mat_C[8][12] <= 
                  mat_A[8][0] * mat_B[0][12] +
                  mat_A[8][1] * mat_B[1][12] +
                  mat_A[8][2] * mat_B[2][12] +
                  mat_A[8][3] * mat_B[3][12] +
                  mat_A[8][4] * mat_B[4][12] +
                  mat_A[8][5] * mat_B[5][12] +
                  mat_A[8][6] * mat_B[6][12] +
                  mat_A[8][7] * mat_B[7][12] +
                  mat_A[8][8] * mat_B[8][12] +
                  mat_A[8][9] * mat_B[9][12] +
                  mat_A[8][10] * mat_B[10][12] +
                  mat_A[8][11] * mat_B[11][12] +
                  mat_A[8][12] * mat_B[12][12] +
                  mat_A[8][13] * mat_B[13][12] +
                  mat_A[8][14] * mat_B[14][12] +
                  mat_A[8][15] * mat_B[15][12] +
                  mat_A[8][16] * mat_B[16][12] +
                  mat_A[8][17] * mat_B[17][12] +
                  mat_A[8][18] * mat_B[18][12] +
                  mat_A[8][19] * mat_B[19][12] +
                  mat_A[8][20] * mat_B[20][12] +
                  mat_A[8][21] * mat_B[21][12] +
                  mat_A[8][22] * mat_B[22][12] +
                  mat_A[8][23] * mat_B[23][12] +
                  mat_A[8][24] * mat_B[24][12] +
                  mat_A[8][25] * mat_B[25][12] +
                  mat_A[8][26] * mat_B[26][12] +
                  mat_A[8][27] * mat_B[27][12] +
                  mat_A[8][28] * mat_B[28][12] +
                  mat_A[8][29] * mat_B[29][12] +
                  mat_A[8][30] * mat_B[30][12] +
                  mat_A[8][31] * mat_B[31][12];
    mat_C[8][13] <= 
                  mat_A[8][0] * mat_B[0][13] +
                  mat_A[8][1] * mat_B[1][13] +
                  mat_A[8][2] * mat_B[2][13] +
                  mat_A[8][3] * mat_B[3][13] +
                  mat_A[8][4] * mat_B[4][13] +
                  mat_A[8][5] * mat_B[5][13] +
                  mat_A[8][6] * mat_B[6][13] +
                  mat_A[8][7] * mat_B[7][13] +
                  mat_A[8][8] * mat_B[8][13] +
                  mat_A[8][9] * mat_B[9][13] +
                  mat_A[8][10] * mat_B[10][13] +
                  mat_A[8][11] * mat_B[11][13] +
                  mat_A[8][12] * mat_B[12][13] +
                  mat_A[8][13] * mat_B[13][13] +
                  mat_A[8][14] * mat_B[14][13] +
                  mat_A[8][15] * mat_B[15][13] +
                  mat_A[8][16] * mat_B[16][13] +
                  mat_A[8][17] * mat_B[17][13] +
                  mat_A[8][18] * mat_B[18][13] +
                  mat_A[8][19] * mat_B[19][13] +
                  mat_A[8][20] * mat_B[20][13] +
                  mat_A[8][21] * mat_B[21][13] +
                  mat_A[8][22] * mat_B[22][13] +
                  mat_A[8][23] * mat_B[23][13] +
                  mat_A[8][24] * mat_B[24][13] +
                  mat_A[8][25] * mat_B[25][13] +
                  mat_A[8][26] * mat_B[26][13] +
                  mat_A[8][27] * mat_B[27][13] +
                  mat_A[8][28] * mat_B[28][13] +
                  mat_A[8][29] * mat_B[29][13] +
                  mat_A[8][30] * mat_B[30][13] +
                  mat_A[8][31] * mat_B[31][13];
    mat_C[8][14] <= 
                  mat_A[8][0] * mat_B[0][14] +
                  mat_A[8][1] * mat_B[1][14] +
                  mat_A[8][2] * mat_B[2][14] +
                  mat_A[8][3] * mat_B[3][14] +
                  mat_A[8][4] * mat_B[4][14] +
                  mat_A[8][5] * mat_B[5][14] +
                  mat_A[8][6] * mat_B[6][14] +
                  mat_A[8][7] * mat_B[7][14] +
                  mat_A[8][8] * mat_B[8][14] +
                  mat_A[8][9] * mat_B[9][14] +
                  mat_A[8][10] * mat_B[10][14] +
                  mat_A[8][11] * mat_B[11][14] +
                  mat_A[8][12] * mat_B[12][14] +
                  mat_A[8][13] * mat_B[13][14] +
                  mat_A[8][14] * mat_B[14][14] +
                  mat_A[8][15] * mat_B[15][14] +
                  mat_A[8][16] * mat_B[16][14] +
                  mat_A[8][17] * mat_B[17][14] +
                  mat_A[8][18] * mat_B[18][14] +
                  mat_A[8][19] * mat_B[19][14] +
                  mat_A[8][20] * mat_B[20][14] +
                  mat_A[8][21] * mat_B[21][14] +
                  mat_A[8][22] * mat_B[22][14] +
                  mat_A[8][23] * mat_B[23][14] +
                  mat_A[8][24] * mat_B[24][14] +
                  mat_A[8][25] * mat_B[25][14] +
                  mat_A[8][26] * mat_B[26][14] +
                  mat_A[8][27] * mat_B[27][14] +
                  mat_A[8][28] * mat_B[28][14] +
                  mat_A[8][29] * mat_B[29][14] +
                  mat_A[8][30] * mat_B[30][14] +
                  mat_A[8][31] * mat_B[31][14];
    mat_C[8][15] <= 
                  mat_A[8][0] * mat_B[0][15] +
                  mat_A[8][1] * mat_B[1][15] +
                  mat_A[8][2] * mat_B[2][15] +
                  mat_A[8][3] * mat_B[3][15] +
                  mat_A[8][4] * mat_B[4][15] +
                  mat_A[8][5] * mat_B[5][15] +
                  mat_A[8][6] * mat_B[6][15] +
                  mat_A[8][7] * mat_B[7][15] +
                  mat_A[8][8] * mat_B[8][15] +
                  mat_A[8][9] * mat_B[9][15] +
                  mat_A[8][10] * mat_B[10][15] +
                  mat_A[8][11] * mat_B[11][15] +
                  mat_A[8][12] * mat_B[12][15] +
                  mat_A[8][13] * mat_B[13][15] +
                  mat_A[8][14] * mat_B[14][15] +
                  mat_A[8][15] * mat_B[15][15] +
                  mat_A[8][16] * mat_B[16][15] +
                  mat_A[8][17] * mat_B[17][15] +
                  mat_A[8][18] * mat_B[18][15] +
                  mat_A[8][19] * mat_B[19][15] +
                  mat_A[8][20] * mat_B[20][15] +
                  mat_A[8][21] * mat_B[21][15] +
                  mat_A[8][22] * mat_B[22][15] +
                  mat_A[8][23] * mat_B[23][15] +
                  mat_A[8][24] * mat_B[24][15] +
                  mat_A[8][25] * mat_B[25][15] +
                  mat_A[8][26] * mat_B[26][15] +
                  mat_A[8][27] * mat_B[27][15] +
                  mat_A[8][28] * mat_B[28][15] +
                  mat_A[8][29] * mat_B[29][15] +
                  mat_A[8][30] * mat_B[30][15] +
                  mat_A[8][31] * mat_B[31][15];
    mat_C[8][16] <= 
                  mat_A[8][0] * mat_B[0][16] +
                  mat_A[8][1] * mat_B[1][16] +
                  mat_A[8][2] * mat_B[2][16] +
                  mat_A[8][3] * mat_B[3][16] +
                  mat_A[8][4] * mat_B[4][16] +
                  mat_A[8][5] * mat_B[5][16] +
                  mat_A[8][6] * mat_B[6][16] +
                  mat_A[8][7] * mat_B[7][16] +
                  mat_A[8][8] * mat_B[8][16] +
                  mat_A[8][9] * mat_B[9][16] +
                  mat_A[8][10] * mat_B[10][16] +
                  mat_A[8][11] * mat_B[11][16] +
                  mat_A[8][12] * mat_B[12][16] +
                  mat_A[8][13] * mat_B[13][16] +
                  mat_A[8][14] * mat_B[14][16] +
                  mat_A[8][15] * mat_B[15][16] +
                  mat_A[8][16] * mat_B[16][16] +
                  mat_A[8][17] * mat_B[17][16] +
                  mat_A[8][18] * mat_B[18][16] +
                  mat_A[8][19] * mat_B[19][16] +
                  mat_A[8][20] * mat_B[20][16] +
                  mat_A[8][21] * mat_B[21][16] +
                  mat_A[8][22] * mat_B[22][16] +
                  mat_A[8][23] * mat_B[23][16] +
                  mat_A[8][24] * mat_B[24][16] +
                  mat_A[8][25] * mat_B[25][16] +
                  mat_A[8][26] * mat_B[26][16] +
                  mat_A[8][27] * mat_B[27][16] +
                  mat_A[8][28] * mat_B[28][16] +
                  mat_A[8][29] * mat_B[29][16] +
                  mat_A[8][30] * mat_B[30][16] +
                  mat_A[8][31] * mat_B[31][16];
    mat_C[8][17] <= 
                  mat_A[8][0] * mat_B[0][17] +
                  mat_A[8][1] * mat_B[1][17] +
                  mat_A[8][2] * mat_B[2][17] +
                  mat_A[8][3] * mat_B[3][17] +
                  mat_A[8][4] * mat_B[4][17] +
                  mat_A[8][5] * mat_B[5][17] +
                  mat_A[8][6] * mat_B[6][17] +
                  mat_A[8][7] * mat_B[7][17] +
                  mat_A[8][8] * mat_B[8][17] +
                  mat_A[8][9] * mat_B[9][17] +
                  mat_A[8][10] * mat_B[10][17] +
                  mat_A[8][11] * mat_B[11][17] +
                  mat_A[8][12] * mat_B[12][17] +
                  mat_A[8][13] * mat_B[13][17] +
                  mat_A[8][14] * mat_B[14][17] +
                  mat_A[8][15] * mat_B[15][17] +
                  mat_A[8][16] * mat_B[16][17] +
                  mat_A[8][17] * mat_B[17][17] +
                  mat_A[8][18] * mat_B[18][17] +
                  mat_A[8][19] * mat_B[19][17] +
                  mat_A[8][20] * mat_B[20][17] +
                  mat_A[8][21] * mat_B[21][17] +
                  mat_A[8][22] * mat_B[22][17] +
                  mat_A[8][23] * mat_B[23][17] +
                  mat_A[8][24] * mat_B[24][17] +
                  mat_A[8][25] * mat_B[25][17] +
                  mat_A[8][26] * mat_B[26][17] +
                  mat_A[8][27] * mat_B[27][17] +
                  mat_A[8][28] * mat_B[28][17] +
                  mat_A[8][29] * mat_B[29][17] +
                  mat_A[8][30] * mat_B[30][17] +
                  mat_A[8][31] * mat_B[31][17];
    mat_C[8][18] <= 
                  mat_A[8][0] * mat_B[0][18] +
                  mat_A[8][1] * mat_B[1][18] +
                  mat_A[8][2] * mat_B[2][18] +
                  mat_A[8][3] * mat_B[3][18] +
                  mat_A[8][4] * mat_B[4][18] +
                  mat_A[8][5] * mat_B[5][18] +
                  mat_A[8][6] * mat_B[6][18] +
                  mat_A[8][7] * mat_B[7][18] +
                  mat_A[8][8] * mat_B[8][18] +
                  mat_A[8][9] * mat_B[9][18] +
                  mat_A[8][10] * mat_B[10][18] +
                  mat_A[8][11] * mat_B[11][18] +
                  mat_A[8][12] * mat_B[12][18] +
                  mat_A[8][13] * mat_B[13][18] +
                  mat_A[8][14] * mat_B[14][18] +
                  mat_A[8][15] * mat_B[15][18] +
                  mat_A[8][16] * mat_B[16][18] +
                  mat_A[8][17] * mat_B[17][18] +
                  mat_A[8][18] * mat_B[18][18] +
                  mat_A[8][19] * mat_B[19][18] +
                  mat_A[8][20] * mat_B[20][18] +
                  mat_A[8][21] * mat_B[21][18] +
                  mat_A[8][22] * mat_B[22][18] +
                  mat_A[8][23] * mat_B[23][18] +
                  mat_A[8][24] * mat_B[24][18] +
                  mat_A[8][25] * mat_B[25][18] +
                  mat_A[8][26] * mat_B[26][18] +
                  mat_A[8][27] * mat_B[27][18] +
                  mat_A[8][28] * mat_B[28][18] +
                  mat_A[8][29] * mat_B[29][18] +
                  mat_A[8][30] * mat_B[30][18] +
                  mat_A[8][31] * mat_B[31][18];
    mat_C[8][19] <= 
                  mat_A[8][0] * mat_B[0][19] +
                  mat_A[8][1] * mat_B[1][19] +
                  mat_A[8][2] * mat_B[2][19] +
                  mat_A[8][3] * mat_B[3][19] +
                  mat_A[8][4] * mat_B[4][19] +
                  mat_A[8][5] * mat_B[5][19] +
                  mat_A[8][6] * mat_B[6][19] +
                  mat_A[8][7] * mat_B[7][19] +
                  mat_A[8][8] * mat_B[8][19] +
                  mat_A[8][9] * mat_B[9][19] +
                  mat_A[8][10] * mat_B[10][19] +
                  mat_A[8][11] * mat_B[11][19] +
                  mat_A[8][12] * mat_B[12][19] +
                  mat_A[8][13] * mat_B[13][19] +
                  mat_A[8][14] * mat_B[14][19] +
                  mat_A[8][15] * mat_B[15][19] +
                  mat_A[8][16] * mat_B[16][19] +
                  mat_A[8][17] * mat_B[17][19] +
                  mat_A[8][18] * mat_B[18][19] +
                  mat_A[8][19] * mat_B[19][19] +
                  mat_A[8][20] * mat_B[20][19] +
                  mat_A[8][21] * mat_B[21][19] +
                  mat_A[8][22] * mat_B[22][19] +
                  mat_A[8][23] * mat_B[23][19] +
                  mat_A[8][24] * mat_B[24][19] +
                  mat_A[8][25] * mat_B[25][19] +
                  mat_A[8][26] * mat_B[26][19] +
                  mat_A[8][27] * mat_B[27][19] +
                  mat_A[8][28] * mat_B[28][19] +
                  mat_A[8][29] * mat_B[29][19] +
                  mat_A[8][30] * mat_B[30][19] +
                  mat_A[8][31] * mat_B[31][19];
    mat_C[8][20] <= 
                  mat_A[8][0] * mat_B[0][20] +
                  mat_A[8][1] * mat_B[1][20] +
                  mat_A[8][2] * mat_B[2][20] +
                  mat_A[8][3] * mat_B[3][20] +
                  mat_A[8][4] * mat_B[4][20] +
                  mat_A[8][5] * mat_B[5][20] +
                  mat_A[8][6] * mat_B[6][20] +
                  mat_A[8][7] * mat_B[7][20] +
                  mat_A[8][8] * mat_B[8][20] +
                  mat_A[8][9] * mat_B[9][20] +
                  mat_A[8][10] * mat_B[10][20] +
                  mat_A[8][11] * mat_B[11][20] +
                  mat_A[8][12] * mat_B[12][20] +
                  mat_A[8][13] * mat_B[13][20] +
                  mat_A[8][14] * mat_B[14][20] +
                  mat_A[8][15] * mat_B[15][20] +
                  mat_A[8][16] * mat_B[16][20] +
                  mat_A[8][17] * mat_B[17][20] +
                  mat_A[8][18] * mat_B[18][20] +
                  mat_A[8][19] * mat_B[19][20] +
                  mat_A[8][20] * mat_B[20][20] +
                  mat_A[8][21] * mat_B[21][20] +
                  mat_A[8][22] * mat_B[22][20] +
                  mat_A[8][23] * mat_B[23][20] +
                  mat_A[8][24] * mat_B[24][20] +
                  mat_A[8][25] * mat_B[25][20] +
                  mat_A[8][26] * mat_B[26][20] +
                  mat_A[8][27] * mat_B[27][20] +
                  mat_A[8][28] * mat_B[28][20] +
                  mat_A[8][29] * mat_B[29][20] +
                  mat_A[8][30] * mat_B[30][20] +
                  mat_A[8][31] * mat_B[31][20];
    mat_C[8][21] <= 
                  mat_A[8][0] * mat_B[0][21] +
                  mat_A[8][1] * mat_B[1][21] +
                  mat_A[8][2] * mat_B[2][21] +
                  mat_A[8][3] * mat_B[3][21] +
                  mat_A[8][4] * mat_B[4][21] +
                  mat_A[8][5] * mat_B[5][21] +
                  mat_A[8][6] * mat_B[6][21] +
                  mat_A[8][7] * mat_B[7][21] +
                  mat_A[8][8] * mat_B[8][21] +
                  mat_A[8][9] * mat_B[9][21] +
                  mat_A[8][10] * mat_B[10][21] +
                  mat_A[8][11] * mat_B[11][21] +
                  mat_A[8][12] * mat_B[12][21] +
                  mat_A[8][13] * mat_B[13][21] +
                  mat_A[8][14] * mat_B[14][21] +
                  mat_A[8][15] * mat_B[15][21] +
                  mat_A[8][16] * mat_B[16][21] +
                  mat_A[8][17] * mat_B[17][21] +
                  mat_A[8][18] * mat_B[18][21] +
                  mat_A[8][19] * mat_B[19][21] +
                  mat_A[8][20] * mat_B[20][21] +
                  mat_A[8][21] * mat_B[21][21] +
                  mat_A[8][22] * mat_B[22][21] +
                  mat_A[8][23] * mat_B[23][21] +
                  mat_A[8][24] * mat_B[24][21] +
                  mat_A[8][25] * mat_B[25][21] +
                  mat_A[8][26] * mat_B[26][21] +
                  mat_A[8][27] * mat_B[27][21] +
                  mat_A[8][28] * mat_B[28][21] +
                  mat_A[8][29] * mat_B[29][21] +
                  mat_A[8][30] * mat_B[30][21] +
                  mat_A[8][31] * mat_B[31][21];
    mat_C[8][22] <= 
                  mat_A[8][0] * mat_B[0][22] +
                  mat_A[8][1] * mat_B[1][22] +
                  mat_A[8][2] * mat_B[2][22] +
                  mat_A[8][3] * mat_B[3][22] +
                  mat_A[8][4] * mat_B[4][22] +
                  mat_A[8][5] * mat_B[5][22] +
                  mat_A[8][6] * mat_B[6][22] +
                  mat_A[8][7] * mat_B[7][22] +
                  mat_A[8][8] * mat_B[8][22] +
                  mat_A[8][9] * mat_B[9][22] +
                  mat_A[8][10] * mat_B[10][22] +
                  mat_A[8][11] * mat_B[11][22] +
                  mat_A[8][12] * mat_B[12][22] +
                  mat_A[8][13] * mat_B[13][22] +
                  mat_A[8][14] * mat_B[14][22] +
                  mat_A[8][15] * mat_B[15][22] +
                  mat_A[8][16] * mat_B[16][22] +
                  mat_A[8][17] * mat_B[17][22] +
                  mat_A[8][18] * mat_B[18][22] +
                  mat_A[8][19] * mat_B[19][22] +
                  mat_A[8][20] * mat_B[20][22] +
                  mat_A[8][21] * mat_B[21][22] +
                  mat_A[8][22] * mat_B[22][22] +
                  mat_A[8][23] * mat_B[23][22] +
                  mat_A[8][24] * mat_B[24][22] +
                  mat_A[8][25] * mat_B[25][22] +
                  mat_A[8][26] * mat_B[26][22] +
                  mat_A[8][27] * mat_B[27][22] +
                  mat_A[8][28] * mat_B[28][22] +
                  mat_A[8][29] * mat_B[29][22] +
                  mat_A[8][30] * mat_B[30][22] +
                  mat_A[8][31] * mat_B[31][22];
    mat_C[8][23] <= 
                  mat_A[8][0] * mat_B[0][23] +
                  mat_A[8][1] * mat_B[1][23] +
                  mat_A[8][2] * mat_B[2][23] +
                  mat_A[8][3] * mat_B[3][23] +
                  mat_A[8][4] * mat_B[4][23] +
                  mat_A[8][5] * mat_B[5][23] +
                  mat_A[8][6] * mat_B[6][23] +
                  mat_A[8][7] * mat_B[7][23] +
                  mat_A[8][8] * mat_B[8][23] +
                  mat_A[8][9] * mat_B[9][23] +
                  mat_A[8][10] * mat_B[10][23] +
                  mat_A[8][11] * mat_B[11][23] +
                  mat_A[8][12] * mat_B[12][23] +
                  mat_A[8][13] * mat_B[13][23] +
                  mat_A[8][14] * mat_B[14][23] +
                  mat_A[8][15] * mat_B[15][23] +
                  mat_A[8][16] * mat_B[16][23] +
                  mat_A[8][17] * mat_B[17][23] +
                  mat_A[8][18] * mat_B[18][23] +
                  mat_A[8][19] * mat_B[19][23] +
                  mat_A[8][20] * mat_B[20][23] +
                  mat_A[8][21] * mat_B[21][23] +
                  mat_A[8][22] * mat_B[22][23] +
                  mat_A[8][23] * mat_B[23][23] +
                  mat_A[8][24] * mat_B[24][23] +
                  mat_A[8][25] * mat_B[25][23] +
                  mat_A[8][26] * mat_B[26][23] +
                  mat_A[8][27] * mat_B[27][23] +
                  mat_A[8][28] * mat_B[28][23] +
                  mat_A[8][29] * mat_B[29][23] +
                  mat_A[8][30] * mat_B[30][23] +
                  mat_A[8][31] * mat_B[31][23];
    mat_C[8][24] <= 
                  mat_A[8][0] * mat_B[0][24] +
                  mat_A[8][1] * mat_B[1][24] +
                  mat_A[8][2] * mat_B[2][24] +
                  mat_A[8][3] * mat_B[3][24] +
                  mat_A[8][4] * mat_B[4][24] +
                  mat_A[8][5] * mat_B[5][24] +
                  mat_A[8][6] * mat_B[6][24] +
                  mat_A[8][7] * mat_B[7][24] +
                  mat_A[8][8] * mat_B[8][24] +
                  mat_A[8][9] * mat_B[9][24] +
                  mat_A[8][10] * mat_B[10][24] +
                  mat_A[8][11] * mat_B[11][24] +
                  mat_A[8][12] * mat_B[12][24] +
                  mat_A[8][13] * mat_B[13][24] +
                  mat_A[8][14] * mat_B[14][24] +
                  mat_A[8][15] * mat_B[15][24] +
                  mat_A[8][16] * mat_B[16][24] +
                  mat_A[8][17] * mat_B[17][24] +
                  mat_A[8][18] * mat_B[18][24] +
                  mat_A[8][19] * mat_B[19][24] +
                  mat_A[8][20] * mat_B[20][24] +
                  mat_A[8][21] * mat_B[21][24] +
                  mat_A[8][22] * mat_B[22][24] +
                  mat_A[8][23] * mat_B[23][24] +
                  mat_A[8][24] * mat_B[24][24] +
                  mat_A[8][25] * mat_B[25][24] +
                  mat_A[8][26] * mat_B[26][24] +
                  mat_A[8][27] * mat_B[27][24] +
                  mat_A[8][28] * mat_B[28][24] +
                  mat_A[8][29] * mat_B[29][24] +
                  mat_A[8][30] * mat_B[30][24] +
                  mat_A[8][31] * mat_B[31][24];
    mat_C[8][25] <= 
                  mat_A[8][0] * mat_B[0][25] +
                  mat_A[8][1] * mat_B[1][25] +
                  mat_A[8][2] * mat_B[2][25] +
                  mat_A[8][3] * mat_B[3][25] +
                  mat_A[8][4] * mat_B[4][25] +
                  mat_A[8][5] * mat_B[5][25] +
                  mat_A[8][6] * mat_B[6][25] +
                  mat_A[8][7] * mat_B[7][25] +
                  mat_A[8][8] * mat_B[8][25] +
                  mat_A[8][9] * mat_B[9][25] +
                  mat_A[8][10] * mat_B[10][25] +
                  mat_A[8][11] * mat_B[11][25] +
                  mat_A[8][12] * mat_B[12][25] +
                  mat_A[8][13] * mat_B[13][25] +
                  mat_A[8][14] * mat_B[14][25] +
                  mat_A[8][15] * mat_B[15][25] +
                  mat_A[8][16] * mat_B[16][25] +
                  mat_A[8][17] * mat_B[17][25] +
                  mat_A[8][18] * mat_B[18][25] +
                  mat_A[8][19] * mat_B[19][25] +
                  mat_A[8][20] * mat_B[20][25] +
                  mat_A[8][21] * mat_B[21][25] +
                  mat_A[8][22] * mat_B[22][25] +
                  mat_A[8][23] * mat_B[23][25] +
                  mat_A[8][24] * mat_B[24][25] +
                  mat_A[8][25] * mat_B[25][25] +
                  mat_A[8][26] * mat_B[26][25] +
                  mat_A[8][27] * mat_B[27][25] +
                  mat_A[8][28] * mat_B[28][25] +
                  mat_A[8][29] * mat_B[29][25] +
                  mat_A[8][30] * mat_B[30][25] +
                  mat_A[8][31] * mat_B[31][25];
    mat_C[8][26] <= 
                  mat_A[8][0] * mat_B[0][26] +
                  mat_A[8][1] * mat_B[1][26] +
                  mat_A[8][2] * mat_B[2][26] +
                  mat_A[8][3] * mat_B[3][26] +
                  mat_A[8][4] * mat_B[4][26] +
                  mat_A[8][5] * mat_B[5][26] +
                  mat_A[8][6] * mat_B[6][26] +
                  mat_A[8][7] * mat_B[7][26] +
                  mat_A[8][8] * mat_B[8][26] +
                  mat_A[8][9] * mat_B[9][26] +
                  mat_A[8][10] * mat_B[10][26] +
                  mat_A[8][11] * mat_B[11][26] +
                  mat_A[8][12] * mat_B[12][26] +
                  mat_A[8][13] * mat_B[13][26] +
                  mat_A[8][14] * mat_B[14][26] +
                  mat_A[8][15] * mat_B[15][26] +
                  mat_A[8][16] * mat_B[16][26] +
                  mat_A[8][17] * mat_B[17][26] +
                  mat_A[8][18] * mat_B[18][26] +
                  mat_A[8][19] * mat_B[19][26] +
                  mat_A[8][20] * mat_B[20][26] +
                  mat_A[8][21] * mat_B[21][26] +
                  mat_A[8][22] * mat_B[22][26] +
                  mat_A[8][23] * mat_B[23][26] +
                  mat_A[8][24] * mat_B[24][26] +
                  mat_A[8][25] * mat_B[25][26] +
                  mat_A[8][26] * mat_B[26][26] +
                  mat_A[8][27] * mat_B[27][26] +
                  mat_A[8][28] * mat_B[28][26] +
                  mat_A[8][29] * mat_B[29][26] +
                  mat_A[8][30] * mat_B[30][26] +
                  mat_A[8][31] * mat_B[31][26];
    mat_C[8][27] <= 
                  mat_A[8][0] * mat_B[0][27] +
                  mat_A[8][1] * mat_B[1][27] +
                  mat_A[8][2] * mat_B[2][27] +
                  mat_A[8][3] * mat_B[3][27] +
                  mat_A[8][4] * mat_B[4][27] +
                  mat_A[8][5] * mat_B[5][27] +
                  mat_A[8][6] * mat_B[6][27] +
                  mat_A[8][7] * mat_B[7][27] +
                  mat_A[8][8] * mat_B[8][27] +
                  mat_A[8][9] * mat_B[9][27] +
                  mat_A[8][10] * mat_B[10][27] +
                  mat_A[8][11] * mat_B[11][27] +
                  mat_A[8][12] * mat_B[12][27] +
                  mat_A[8][13] * mat_B[13][27] +
                  mat_A[8][14] * mat_B[14][27] +
                  mat_A[8][15] * mat_B[15][27] +
                  mat_A[8][16] * mat_B[16][27] +
                  mat_A[8][17] * mat_B[17][27] +
                  mat_A[8][18] * mat_B[18][27] +
                  mat_A[8][19] * mat_B[19][27] +
                  mat_A[8][20] * mat_B[20][27] +
                  mat_A[8][21] * mat_B[21][27] +
                  mat_A[8][22] * mat_B[22][27] +
                  mat_A[8][23] * mat_B[23][27] +
                  mat_A[8][24] * mat_B[24][27] +
                  mat_A[8][25] * mat_B[25][27] +
                  mat_A[8][26] * mat_B[26][27] +
                  mat_A[8][27] * mat_B[27][27] +
                  mat_A[8][28] * mat_B[28][27] +
                  mat_A[8][29] * mat_B[29][27] +
                  mat_A[8][30] * mat_B[30][27] +
                  mat_A[8][31] * mat_B[31][27];
    mat_C[8][28] <= 
                  mat_A[8][0] * mat_B[0][28] +
                  mat_A[8][1] * mat_B[1][28] +
                  mat_A[8][2] * mat_B[2][28] +
                  mat_A[8][3] * mat_B[3][28] +
                  mat_A[8][4] * mat_B[4][28] +
                  mat_A[8][5] * mat_B[5][28] +
                  mat_A[8][6] * mat_B[6][28] +
                  mat_A[8][7] * mat_B[7][28] +
                  mat_A[8][8] * mat_B[8][28] +
                  mat_A[8][9] * mat_B[9][28] +
                  mat_A[8][10] * mat_B[10][28] +
                  mat_A[8][11] * mat_B[11][28] +
                  mat_A[8][12] * mat_B[12][28] +
                  mat_A[8][13] * mat_B[13][28] +
                  mat_A[8][14] * mat_B[14][28] +
                  mat_A[8][15] * mat_B[15][28] +
                  mat_A[8][16] * mat_B[16][28] +
                  mat_A[8][17] * mat_B[17][28] +
                  mat_A[8][18] * mat_B[18][28] +
                  mat_A[8][19] * mat_B[19][28] +
                  mat_A[8][20] * mat_B[20][28] +
                  mat_A[8][21] * mat_B[21][28] +
                  mat_A[8][22] * mat_B[22][28] +
                  mat_A[8][23] * mat_B[23][28] +
                  mat_A[8][24] * mat_B[24][28] +
                  mat_A[8][25] * mat_B[25][28] +
                  mat_A[8][26] * mat_B[26][28] +
                  mat_A[8][27] * mat_B[27][28] +
                  mat_A[8][28] * mat_B[28][28] +
                  mat_A[8][29] * mat_B[29][28] +
                  mat_A[8][30] * mat_B[30][28] +
                  mat_A[8][31] * mat_B[31][28];
    mat_C[8][29] <= 
                  mat_A[8][0] * mat_B[0][29] +
                  mat_A[8][1] * mat_B[1][29] +
                  mat_A[8][2] * mat_B[2][29] +
                  mat_A[8][3] * mat_B[3][29] +
                  mat_A[8][4] * mat_B[4][29] +
                  mat_A[8][5] * mat_B[5][29] +
                  mat_A[8][6] * mat_B[6][29] +
                  mat_A[8][7] * mat_B[7][29] +
                  mat_A[8][8] * mat_B[8][29] +
                  mat_A[8][9] * mat_B[9][29] +
                  mat_A[8][10] * mat_B[10][29] +
                  mat_A[8][11] * mat_B[11][29] +
                  mat_A[8][12] * mat_B[12][29] +
                  mat_A[8][13] * mat_B[13][29] +
                  mat_A[8][14] * mat_B[14][29] +
                  mat_A[8][15] * mat_B[15][29] +
                  mat_A[8][16] * mat_B[16][29] +
                  mat_A[8][17] * mat_B[17][29] +
                  mat_A[8][18] * mat_B[18][29] +
                  mat_A[8][19] * mat_B[19][29] +
                  mat_A[8][20] * mat_B[20][29] +
                  mat_A[8][21] * mat_B[21][29] +
                  mat_A[8][22] * mat_B[22][29] +
                  mat_A[8][23] * mat_B[23][29] +
                  mat_A[8][24] * mat_B[24][29] +
                  mat_A[8][25] * mat_B[25][29] +
                  mat_A[8][26] * mat_B[26][29] +
                  mat_A[8][27] * mat_B[27][29] +
                  mat_A[8][28] * mat_B[28][29] +
                  mat_A[8][29] * mat_B[29][29] +
                  mat_A[8][30] * mat_B[30][29] +
                  mat_A[8][31] * mat_B[31][29];
    mat_C[8][30] <= 
                  mat_A[8][0] * mat_B[0][30] +
                  mat_A[8][1] * mat_B[1][30] +
                  mat_A[8][2] * mat_B[2][30] +
                  mat_A[8][3] * mat_B[3][30] +
                  mat_A[8][4] * mat_B[4][30] +
                  mat_A[8][5] * mat_B[5][30] +
                  mat_A[8][6] * mat_B[6][30] +
                  mat_A[8][7] * mat_B[7][30] +
                  mat_A[8][8] * mat_B[8][30] +
                  mat_A[8][9] * mat_B[9][30] +
                  mat_A[8][10] * mat_B[10][30] +
                  mat_A[8][11] * mat_B[11][30] +
                  mat_A[8][12] * mat_B[12][30] +
                  mat_A[8][13] * mat_B[13][30] +
                  mat_A[8][14] * mat_B[14][30] +
                  mat_A[8][15] * mat_B[15][30] +
                  mat_A[8][16] * mat_B[16][30] +
                  mat_A[8][17] * mat_B[17][30] +
                  mat_A[8][18] * mat_B[18][30] +
                  mat_A[8][19] * mat_B[19][30] +
                  mat_A[8][20] * mat_B[20][30] +
                  mat_A[8][21] * mat_B[21][30] +
                  mat_A[8][22] * mat_B[22][30] +
                  mat_A[8][23] * mat_B[23][30] +
                  mat_A[8][24] * mat_B[24][30] +
                  mat_A[8][25] * mat_B[25][30] +
                  mat_A[8][26] * mat_B[26][30] +
                  mat_A[8][27] * mat_B[27][30] +
                  mat_A[8][28] * mat_B[28][30] +
                  mat_A[8][29] * mat_B[29][30] +
                  mat_A[8][30] * mat_B[30][30] +
                  mat_A[8][31] * mat_B[31][30];
    mat_C[8][31] <= 
                  mat_A[8][0] * mat_B[0][31] +
                  mat_A[8][1] * mat_B[1][31] +
                  mat_A[8][2] * mat_B[2][31] +
                  mat_A[8][3] * mat_B[3][31] +
                  mat_A[8][4] * mat_B[4][31] +
                  mat_A[8][5] * mat_B[5][31] +
                  mat_A[8][6] * mat_B[6][31] +
                  mat_A[8][7] * mat_B[7][31] +
                  mat_A[8][8] * mat_B[8][31] +
                  mat_A[8][9] * mat_B[9][31] +
                  mat_A[8][10] * mat_B[10][31] +
                  mat_A[8][11] * mat_B[11][31] +
                  mat_A[8][12] * mat_B[12][31] +
                  mat_A[8][13] * mat_B[13][31] +
                  mat_A[8][14] * mat_B[14][31] +
                  mat_A[8][15] * mat_B[15][31] +
                  mat_A[8][16] * mat_B[16][31] +
                  mat_A[8][17] * mat_B[17][31] +
                  mat_A[8][18] * mat_B[18][31] +
                  mat_A[8][19] * mat_B[19][31] +
                  mat_A[8][20] * mat_B[20][31] +
                  mat_A[8][21] * mat_B[21][31] +
                  mat_A[8][22] * mat_B[22][31] +
                  mat_A[8][23] * mat_B[23][31] +
                  mat_A[8][24] * mat_B[24][31] +
                  mat_A[8][25] * mat_B[25][31] +
                  mat_A[8][26] * mat_B[26][31] +
                  mat_A[8][27] * mat_B[27][31] +
                  mat_A[8][28] * mat_B[28][31] +
                  mat_A[8][29] * mat_B[29][31] +
                  mat_A[8][30] * mat_B[30][31] +
                  mat_A[8][31] * mat_B[31][31];
    mat_C[9][0] <= 
                  mat_A[9][0] * mat_B[0][0] +
                  mat_A[9][1] * mat_B[1][0] +
                  mat_A[9][2] * mat_B[2][0] +
                  mat_A[9][3] * mat_B[3][0] +
                  mat_A[9][4] * mat_B[4][0] +
                  mat_A[9][5] * mat_B[5][0] +
                  mat_A[9][6] * mat_B[6][0] +
                  mat_A[9][7] * mat_B[7][0] +
                  mat_A[9][8] * mat_B[8][0] +
                  mat_A[9][9] * mat_B[9][0] +
                  mat_A[9][10] * mat_B[10][0] +
                  mat_A[9][11] * mat_B[11][0] +
                  mat_A[9][12] * mat_B[12][0] +
                  mat_A[9][13] * mat_B[13][0] +
                  mat_A[9][14] * mat_B[14][0] +
                  mat_A[9][15] * mat_B[15][0] +
                  mat_A[9][16] * mat_B[16][0] +
                  mat_A[9][17] * mat_B[17][0] +
                  mat_A[9][18] * mat_B[18][0] +
                  mat_A[9][19] * mat_B[19][0] +
                  mat_A[9][20] * mat_B[20][0] +
                  mat_A[9][21] * mat_B[21][0] +
                  mat_A[9][22] * mat_B[22][0] +
                  mat_A[9][23] * mat_B[23][0] +
                  mat_A[9][24] * mat_B[24][0] +
                  mat_A[9][25] * mat_B[25][0] +
                  mat_A[9][26] * mat_B[26][0] +
                  mat_A[9][27] * mat_B[27][0] +
                  mat_A[9][28] * mat_B[28][0] +
                  mat_A[9][29] * mat_B[29][0] +
                  mat_A[9][30] * mat_B[30][0] +
                  mat_A[9][31] * mat_B[31][0];
    mat_C[9][1] <= 
                  mat_A[9][0] * mat_B[0][1] +
                  mat_A[9][1] * mat_B[1][1] +
                  mat_A[9][2] * mat_B[2][1] +
                  mat_A[9][3] * mat_B[3][1] +
                  mat_A[9][4] * mat_B[4][1] +
                  mat_A[9][5] * mat_B[5][1] +
                  mat_A[9][6] * mat_B[6][1] +
                  mat_A[9][7] * mat_B[7][1] +
                  mat_A[9][8] * mat_B[8][1] +
                  mat_A[9][9] * mat_B[9][1] +
                  mat_A[9][10] * mat_B[10][1] +
                  mat_A[9][11] * mat_B[11][1] +
                  mat_A[9][12] * mat_B[12][1] +
                  mat_A[9][13] * mat_B[13][1] +
                  mat_A[9][14] * mat_B[14][1] +
                  mat_A[9][15] * mat_B[15][1] +
                  mat_A[9][16] * mat_B[16][1] +
                  mat_A[9][17] * mat_B[17][1] +
                  mat_A[9][18] * mat_B[18][1] +
                  mat_A[9][19] * mat_B[19][1] +
                  mat_A[9][20] * mat_B[20][1] +
                  mat_A[9][21] * mat_B[21][1] +
                  mat_A[9][22] * mat_B[22][1] +
                  mat_A[9][23] * mat_B[23][1] +
                  mat_A[9][24] * mat_B[24][1] +
                  mat_A[9][25] * mat_B[25][1] +
                  mat_A[9][26] * mat_B[26][1] +
                  mat_A[9][27] * mat_B[27][1] +
                  mat_A[9][28] * mat_B[28][1] +
                  mat_A[9][29] * mat_B[29][1] +
                  mat_A[9][30] * mat_B[30][1] +
                  mat_A[9][31] * mat_B[31][1];
    mat_C[9][2] <= 
                  mat_A[9][0] * mat_B[0][2] +
                  mat_A[9][1] * mat_B[1][2] +
                  mat_A[9][2] * mat_B[2][2] +
                  mat_A[9][3] * mat_B[3][2] +
                  mat_A[9][4] * mat_B[4][2] +
                  mat_A[9][5] * mat_B[5][2] +
                  mat_A[9][6] * mat_B[6][2] +
                  mat_A[9][7] * mat_B[7][2] +
                  mat_A[9][8] * mat_B[8][2] +
                  mat_A[9][9] * mat_B[9][2] +
                  mat_A[9][10] * mat_B[10][2] +
                  mat_A[9][11] * mat_B[11][2] +
                  mat_A[9][12] * mat_B[12][2] +
                  mat_A[9][13] * mat_B[13][2] +
                  mat_A[9][14] * mat_B[14][2] +
                  mat_A[9][15] * mat_B[15][2] +
                  mat_A[9][16] * mat_B[16][2] +
                  mat_A[9][17] * mat_B[17][2] +
                  mat_A[9][18] * mat_B[18][2] +
                  mat_A[9][19] * mat_B[19][2] +
                  mat_A[9][20] * mat_B[20][2] +
                  mat_A[9][21] * mat_B[21][2] +
                  mat_A[9][22] * mat_B[22][2] +
                  mat_A[9][23] * mat_B[23][2] +
                  mat_A[9][24] * mat_B[24][2] +
                  mat_A[9][25] * mat_B[25][2] +
                  mat_A[9][26] * mat_B[26][2] +
                  mat_A[9][27] * mat_B[27][2] +
                  mat_A[9][28] * mat_B[28][2] +
                  mat_A[9][29] * mat_B[29][2] +
                  mat_A[9][30] * mat_B[30][2] +
                  mat_A[9][31] * mat_B[31][2];
    mat_C[9][3] <= 
                  mat_A[9][0] * mat_B[0][3] +
                  mat_A[9][1] * mat_B[1][3] +
                  mat_A[9][2] * mat_B[2][3] +
                  mat_A[9][3] * mat_B[3][3] +
                  mat_A[9][4] * mat_B[4][3] +
                  mat_A[9][5] * mat_B[5][3] +
                  mat_A[9][6] * mat_B[6][3] +
                  mat_A[9][7] * mat_B[7][3] +
                  mat_A[9][8] * mat_B[8][3] +
                  mat_A[9][9] * mat_B[9][3] +
                  mat_A[9][10] * mat_B[10][3] +
                  mat_A[9][11] * mat_B[11][3] +
                  mat_A[9][12] * mat_B[12][3] +
                  mat_A[9][13] * mat_B[13][3] +
                  mat_A[9][14] * mat_B[14][3] +
                  mat_A[9][15] * mat_B[15][3] +
                  mat_A[9][16] * mat_B[16][3] +
                  mat_A[9][17] * mat_B[17][3] +
                  mat_A[9][18] * mat_B[18][3] +
                  mat_A[9][19] * mat_B[19][3] +
                  mat_A[9][20] * mat_B[20][3] +
                  mat_A[9][21] * mat_B[21][3] +
                  mat_A[9][22] * mat_B[22][3] +
                  mat_A[9][23] * mat_B[23][3] +
                  mat_A[9][24] * mat_B[24][3] +
                  mat_A[9][25] * mat_B[25][3] +
                  mat_A[9][26] * mat_B[26][3] +
                  mat_A[9][27] * mat_B[27][3] +
                  mat_A[9][28] * mat_B[28][3] +
                  mat_A[9][29] * mat_B[29][3] +
                  mat_A[9][30] * mat_B[30][3] +
                  mat_A[9][31] * mat_B[31][3];
    mat_C[9][4] <= 
                  mat_A[9][0] * mat_B[0][4] +
                  mat_A[9][1] * mat_B[1][4] +
                  mat_A[9][2] * mat_B[2][4] +
                  mat_A[9][3] * mat_B[3][4] +
                  mat_A[9][4] * mat_B[4][4] +
                  mat_A[9][5] * mat_B[5][4] +
                  mat_A[9][6] * mat_B[6][4] +
                  mat_A[9][7] * mat_B[7][4] +
                  mat_A[9][8] * mat_B[8][4] +
                  mat_A[9][9] * mat_B[9][4] +
                  mat_A[9][10] * mat_B[10][4] +
                  mat_A[9][11] * mat_B[11][4] +
                  mat_A[9][12] * mat_B[12][4] +
                  mat_A[9][13] * mat_B[13][4] +
                  mat_A[9][14] * mat_B[14][4] +
                  mat_A[9][15] * mat_B[15][4] +
                  mat_A[9][16] * mat_B[16][4] +
                  mat_A[9][17] * mat_B[17][4] +
                  mat_A[9][18] * mat_B[18][4] +
                  mat_A[9][19] * mat_B[19][4] +
                  mat_A[9][20] * mat_B[20][4] +
                  mat_A[9][21] * mat_B[21][4] +
                  mat_A[9][22] * mat_B[22][4] +
                  mat_A[9][23] * mat_B[23][4] +
                  mat_A[9][24] * mat_B[24][4] +
                  mat_A[9][25] * mat_B[25][4] +
                  mat_A[9][26] * mat_B[26][4] +
                  mat_A[9][27] * mat_B[27][4] +
                  mat_A[9][28] * mat_B[28][4] +
                  mat_A[9][29] * mat_B[29][4] +
                  mat_A[9][30] * mat_B[30][4] +
                  mat_A[9][31] * mat_B[31][4];
    mat_C[9][5] <= 
                  mat_A[9][0] * mat_B[0][5] +
                  mat_A[9][1] * mat_B[1][5] +
                  mat_A[9][2] * mat_B[2][5] +
                  mat_A[9][3] * mat_B[3][5] +
                  mat_A[9][4] * mat_B[4][5] +
                  mat_A[9][5] * mat_B[5][5] +
                  mat_A[9][6] * mat_B[6][5] +
                  mat_A[9][7] * mat_B[7][5] +
                  mat_A[9][8] * mat_B[8][5] +
                  mat_A[9][9] * mat_B[9][5] +
                  mat_A[9][10] * mat_B[10][5] +
                  mat_A[9][11] * mat_B[11][5] +
                  mat_A[9][12] * mat_B[12][5] +
                  mat_A[9][13] * mat_B[13][5] +
                  mat_A[9][14] * mat_B[14][5] +
                  mat_A[9][15] * mat_B[15][5] +
                  mat_A[9][16] * mat_B[16][5] +
                  mat_A[9][17] * mat_B[17][5] +
                  mat_A[9][18] * mat_B[18][5] +
                  mat_A[9][19] * mat_B[19][5] +
                  mat_A[9][20] * mat_B[20][5] +
                  mat_A[9][21] * mat_B[21][5] +
                  mat_A[9][22] * mat_B[22][5] +
                  mat_A[9][23] * mat_B[23][5] +
                  mat_A[9][24] * mat_B[24][5] +
                  mat_A[9][25] * mat_B[25][5] +
                  mat_A[9][26] * mat_B[26][5] +
                  mat_A[9][27] * mat_B[27][5] +
                  mat_A[9][28] * mat_B[28][5] +
                  mat_A[9][29] * mat_B[29][5] +
                  mat_A[9][30] * mat_B[30][5] +
                  mat_A[9][31] * mat_B[31][5];
    mat_C[9][6] <= 
                  mat_A[9][0] * mat_B[0][6] +
                  mat_A[9][1] * mat_B[1][6] +
                  mat_A[9][2] * mat_B[2][6] +
                  mat_A[9][3] * mat_B[3][6] +
                  mat_A[9][4] * mat_B[4][6] +
                  mat_A[9][5] * mat_B[5][6] +
                  mat_A[9][6] * mat_B[6][6] +
                  mat_A[9][7] * mat_B[7][6] +
                  mat_A[9][8] * mat_B[8][6] +
                  mat_A[9][9] * mat_B[9][6] +
                  mat_A[9][10] * mat_B[10][6] +
                  mat_A[9][11] * mat_B[11][6] +
                  mat_A[9][12] * mat_B[12][6] +
                  mat_A[9][13] * mat_B[13][6] +
                  mat_A[9][14] * mat_B[14][6] +
                  mat_A[9][15] * mat_B[15][6] +
                  mat_A[9][16] * mat_B[16][6] +
                  mat_A[9][17] * mat_B[17][6] +
                  mat_A[9][18] * mat_B[18][6] +
                  mat_A[9][19] * mat_B[19][6] +
                  mat_A[9][20] * mat_B[20][6] +
                  mat_A[9][21] * mat_B[21][6] +
                  mat_A[9][22] * mat_B[22][6] +
                  mat_A[9][23] * mat_B[23][6] +
                  mat_A[9][24] * mat_B[24][6] +
                  mat_A[9][25] * mat_B[25][6] +
                  mat_A[9][26] * mat_B[26][6] +
                  mat_A[9][27] * mat_B[27][6] +
                  mat_A[9][28] * mat_B[28][6] +
                  mat_A[9][29] * mat_B[29][6] +
                  mat_A[9][30] * mat_B[30][6] +
                  mat_A[9][31] * mat_B[31][6];
    mat_C[9][7] <= 
                  mat_A[9][0] * mat_B[0][7] +
                  mat_A[9][1] * mat_B[1][7] +
                  mat_A[9][2] * mat_B[2][7] +
                  mat_A[9][3] * mat_B[3][7] +
                  mat_A[9][4] * mat_B[4][7] +
                  mat_A[9][5] * mat_B[5][7] +
                  mat_A[9][6] * mat_B[6][7] +
                  mat_A[9][7] * mat_B[7][7] +
                  mat_A[9][8] * mat_B[8][7] +
                  mat_A[9][9] * mat_B[9][7] +
                  mat_A[9][10] * mat_B[10][7] +
                  mat_A[9][11] * mat_B[11][7] +
                  mat_A[9][12] * mat_B[12][7] +
                  mat_A[9][13] * mat_B[13][7] +
                  mat_A[9][14] * mat_B[14][7] +
                  mat_A[9][15] * mat_B[15][7] +
                  mat_A[9][16] * mat_B[16][7] +
                  mat_A[9][17] * mat_B[17][7] +
                  mat_A[9][18] * mat_B[18][7] +
                  mat_A[9][19] * mat_B[19][7] +
                  mat_A[9][20] * mat_B[20][7] +
                  mat_A[9][21] * mat_B[21][7] +
                  mat_A[9][22] * mat_B[22][7] +
                  mat_A[9][23] * mat_B[23][7] +
                  mat_A[9][24] * mat_B[24][7] +
                  mat_A[9][25] * mat_B[25][7] +
                  mat_A[9][26] * mat_B[26][7] +
                  mat_A[9][27] * mat_B[27][7] +
                  mat_A[9][28] * mat_B[28][7] +
                  mat_A[9][29] * mat_B[29][7] +
                  mat_A[9][30] * mat_B[30][7] +
                  mat_A[9][31] * mat_B[31][7];
    mat_C[9][8] <= 
                  mat_A[9][0] * mat_B[0][8] +
                  mat_A[9][1] * mat_B[1][8] +
                  mat_A[9][2] * mat_B[2][8] +
                  mat_A[9][3] * mat_B[3][8] +
                  mat_A[9][4] * mat_B[4][8] +
                  mat_A[9][5] * mat_B[5][8] +
                  mat_A[9][6] * mat_B[6][8] +
                  mat_A[9][7] * mat_B[7][8] +
                  mat_A[9][8] * mat_B[8][8] +
                  mat_A[9][9] * mat_B[9][8] +
                  mat_A[9][10] * mat_B[10][8] +
                  mat_A[9][11] * mat_B[11][8] +
                  mat_A[9][12] * mat_B[12][8] +
                  mat_A[9][13] * mat_B[13][8] +
                  mat_A[9][14] * mat_B[14][8] +
                  mat_A[9][15] * mat_B[15][8] +
                  mat_A[9][16] * mat_B[16][8] +
                  mat_A[9][17] * mat_B[17][8] +
                  mat_A[9][18] * mat_B[18][8] +
                  mat_A[9][19] * mat_B[19][8] +
                  mat_A[9][20] * mat_B[20][8] +
                  mat_A[9][21] * mat_B[21][8] +
                  mat_A[9][22] * mat_B[22][8] +
                  mat_A[9][23] * mat_B[23][8] +
                  mat_A[9][24] * mat_B[24][8] +
                  mat_A[9][25] * mat_B[25][8] +
                  mat_A[9][26] * mat_B[26][8] +
                  mat_A[9][27] * mat_B[27][8] +
                  mat_A[9][28] * mat_B[28][8] +
                  mat_A[9][29] * mat_B[29][8] +
                  mat_A[9][30] * mat_B[30][8] +
                  mat_A[9][31] * mat_B[31][8];
    mat_C[9][9] <= 
                  mat_A[9][0] * mat_B[0][9] +
                  mat_A[9][1] * mat_B[1][9] +
                  mat_A[9][2] * mat_B[2][9] +
                  mat_A[9][3] * mat_B[3][9] +
                  mat_A[9][4] * mat_B[4][9] +
                  mat_A[9][5] * mat_B[5][9] +
                  mat_A[9][6] * mat_B[6][9] +
                  mat_A[9][7] * mat_B[7][9] +
                  mat_A[9][8] * mat_B[8][9] +
                  mat_A[9][9] * mat_B[9][9] +
                  mat_A[9][10] * mat_B[10][9] +
                  mat_A[9][11] * mat_B[11][9] +
                  mat_A[9][12] * mat_B[12][9] +
                  mat_A[9][13] * mat_B[13][9] +
                  mat_A[9][14] * mat_B[14][9] +
                  mat_A[9][15] * mat_B[15][9] +
                  mat_A[9][16] * mat_B[16][9] +
                  mat_A[9][17] * mat_B[17][9] +
                  mat_A[9][18] * mat_B[18][9] +
                  mat_A[9][19] * mat_B[19][9] +
                  mat_A[9][20] * mat_B[20][9] +
                  mat_A[9][21] * mat_B[21][9] +
                  mat_A[9][22] * mat_B[22][9] +
                  mat_A[9][23] * mat_B[23][9] +
                  mat_A[9][24] * mat_B[24][9] +
                  mat_A[9][25] * mat_B[25][9] +
                  mat_A[9][26] * mat_B[26][9] +
                  mat_A[9][27] * mat_B[27][9] +
                  mat_A[9][28] * mat_B[28][9] +
                  mat_A[9][29] * mat_B[29][9] +
                  mat_A[9][30] * mat_B[30][9] +
                  mat_A[9][31] * mat_B[31][9];
    mat_C[9][10] <= 
                  mat_A[9][0] * mat_B[0][10] +
                  mat_A[9][1] * mat_B[1][10] +
                  mat_A[9][2] * mat_B[2][10] +
                  mat_A[9][3] * mat_B[3][10] +
                  mat_A[9][4] * mat_B[4][10] +
                  mat_A[9][5] * mat_B[5][10] +
                  mat_A[9][6] * mat_B[6][10] +
                  mat_A[9][7] * mat_B[7][10] +
                  mat_A[9][8] * mat_B[8][10] +
                  mat_A[9][9] * mat_B[9][10] +
                  mat_A[9][10] * mat_B[10][10] +
                  mat_A[9][11] * mat_B[11][10] +
                  mat_A[9][12] * mat_B[12][10] +
                  mat_A[9][13] * mat_B[13][10] +
                  mat_A[9][14] * mat_B[14][10] +
                  mat_A[9][15] * mat_B[15][10] +
                  mat_A[9][16] * mat_B[16][10] +
                  mat_A[9][17] * mat_B[17][10] +
                  mat_A[9][18] * mat_B[18][10] +
                  mat_A[9][19] * mat_B[19][10] +
                  mat_A[9][20] * mat_B[20][10] +
                  mat_A[9][21] * mat_B[21][10] +
                  mat_A[9][22] * mat_B[22][10] +
                  mat_A[9][23] * mat_B[23][10] +
                  mat_A[9][24] * mat_B[24][10] +
                  mat_A[9][25] * mat_B[25][10] +
                  mat_A[9][26] * mat_B[26][10] +
                  mat_A[9][27] * mat_B[27][10] +
                  mat_A[9][28] * mat_B[28][10] +
                  mat_A[9][29] * mat_B[29][10] +
                  mat_A[9][30] * mat_B[30][10] +
                  mat_A[9][31] * mat_B[31][10];
    mat_C[9][11] <= 
                  mat_A[9][0] * mat_B[0][11] +
                  mat_A[9][1] * mat_B[1][11] +
                  mat_A[9][2] * mat_B[2][11] +
                  mat_A[9][3] * mat_B[3][11] +
                  mat_A[9][4] * mat_B[4][11] +
                  mat_A[9][5] * mat_B[5][11] +
                  mat_A[9][6] * mat_B[6][11] +
                  mat_A[9][7] * mat_B[7][11] +
                  mat_A[9][8] * mat_B[8][11] +
                  mat_A[9][9] * mat_B[9][11] +
                  mat_A[9][10] * mat_B[10][11] +
                  mat_A[9][11] * mat_B[11][11] +
                  mat_A[9][12] * mat_B[12][11] +
                  mat_A[9][13] * mat_B[13][11] +
                  mat_A[9][14] * mat_B[14][11] +
                  mat_A[9][15] * mat_B[15][11] +
                  mat_A[9][16] * mat_B[16][11] +
                  mat_A[9][17] * mat_B[17][11] +
                  mat_A[9][18] * mat_B[18][11] +
                  mat_A[9][19] * mat_B[19][11] +
                  mat_A[9][20] * mat_B[20][11] +
                  mat_A[9][21] * mat_B[21][11] +
                  mat_A[9][22] * mat_B[22][11] +
                  mat_A[9][23] * mat_B[23][11] +
                  mat_A[9][24] * mat_B[24][11] +
                  mat_A[9][25] * mat_B[25][11] +
                  mat_A[9][26] * mat_B[26][11] +
                  mat_A[9][27] * mat_B[27][11] +
                  mat_A[9][28] * mat_B[28][11] +
                  mat_A[9][29] * mat_B[29][11] +
                  mat_A[9][30] * mat_B[30][11] +
                  mat_A[9][31] * mat_B[31][11];
    mat_C[9][12] <= 
                  mat_A[9][0] * mat_B[0][12] +
                  mat_A[9][1] * mat_B[1][12] +
                  mat_A[9][2] * mat_B[2][12] +
                  mat_A[9][3] * mat_B[3][12] +
                  mat_A[9][4] * mat_B[4][12] +
                  mat_A[9][5] * mat_B[5][12] +
                  mat_A[9][6] * mat_B[6][12] +
                  mat_A[9][7] * mat_B[7][12] +
                  mat_A[9][8] * mat_B[8][12] +
                  mat_A[9][9] * mat_B[9][12] +
                  mat_A[9][10] * mat_B[10][12] +
                  mat_A[9][11] * mat_B[11][12] +
                  mat_A[9][12] * mat_B[12][12] +
                  mat_A[9][13] * mat_B[13][12] +
                  mat_A[9][14] * mat_B[14][12] +
                  mat_A[9][15] * mat_B[15][12] +
                  mat_A[9][16] * mat_B[16][12] +
                  mat_A[9][17] * mat_B[17][12] +
                  mat_A[9][18] * mat_B[18][12] +
                  mat_A[9][19] * mat_B[19][12] +
                  mat_A[9][20] * mat_B[20][12] +
                  mat_A[9][21] * mat_B[21][12] +
                  mat_A[9][22] * mat_B[22][12] +
                  mat_A[9][23] * mat_B[23][12] +
                  mat_A[9][24] * mat_B[24][12] +
                  mat_A[9][25] * mat_B[25][12] +
                  mat_A[9][26] * mat_B[26][12] +
                  mat_A[9][27] * mat_B[27][12] +
                  mat_A[9][28] * mat_B[28][12] +
                  mat_A[9][29] * mat_B[29][12] +
                  mat_A[9][30] * mat_B[30][12] +
                  mat_A[9][31] * mat_B[31][12];
    mat_C[9][13] <= 
                  mat_A[9][0] * mat_B[0][13] +
                  mat_A[9][1] * mat_B[1][13] +
                  mat_A[9][2] * mat_B[2][13] +
                  mat_A[9][3] * mat_B[3][13] +
                  mat_A[9][4] * mat_B[4][13] +
                  mat_A[9][5] * mat_B[5][13] +
                  mat_A[9][6] * mat_B[6][13] +
                  mat_A[9][7] * mat_B[7][13] +
                  mat_A[9][8] * mat_B[8][13] +
                  mat_A[9][9] * mat_B[9][13] +
                  mat_A[9][10] * mat_B[10][13] +
                  mat_A[9][11] * mat_B[11][13] +
                  mat_A[9][12] * mat_B[12][13] +
                  mat_A[9][13] * mat_B[13][13] +
                  mat_A[9][14] * mat_B[14][13] +
                  mat_A[9][15] * mat_B[15][13] +
                  mat_A[9][16] * mat_B[16][13] +
                  mat_A[9][17] * mat_B[17][13] +
                  mat_A[9][18] * mat_B[18][13] +
                  mat_A[9][19] * mat_B[19][13] +
                  mat_A[9][20] * mat_B[20][13] +
                  mat_A[9][21] * mat_B[21][13] +
                  mat_A[9][22] * mat_B[22][13] +
                  mat_A[9][23] * mat_B[23][13] +
                  mat_A[9][24] * mat_B[24][13] +
                  mat_A[9][25] * mat_B[25][13] +
                  mat_A[9][26] * mat_B[26][13] +
                  mat_A[9][27] * mat_B[27][13] +
                  mat_A[9][28] * mat_B[28][13] +
                  mat_A[9][29] * mat_B[29][13] +
                  mat_A[9][30] * mat_B[30][13] +
                  mat_A[9][31] * mat_B[31][13];
    mat_C[9][14] <= 
                  mat_A[9][0] * mat_B[0][14] +
                  mat_A[9][1] * mat_B[1][14] +
                  mat_A[9][2] * mat_B[2][14] +
                  mat_A[9][3] * mat_B[3][14] +
                  mat_A[9][4] * mat_B[4][14] +
                  mat_A[9][5] * mat_B[5][14] +
                  mat_A[9][6] * mat_B[6][14] +
                  mat_A[9][7] * mat_B[7][14] +
                  mat_A[9][8] * mat_B[8][14] +
                  mat_A[9][9] * mat_B[9][14] +
                  mat_A[9][10] * mat_B[10][14] +
                  mat_A[9][11] * mat_B[11][14] +
                  mat_A[9][12] * mat_B[12][14] +
                  mat_A[9][13] * mat_B[13][14] +
                  mat_A[9][14] * mat_B[14][14] +
                  mat_A[9][15] * mat_B[15][14] +
                  mat_A[9][16] * mat_B[16][14] +
                  mat_A[9][17] * mat_B[17][14] +
                  mat_A[9][18] * mat_B[18][14] +
                  mat_A[9][19] * mat_B[19][14] +
                  mat_A[9][20] * mat_B[20][14] +
                  mat_A[9][21] * mat_B[21][14] +
                  mat_A[9][22] * mat_B[22][14] +
                  mat_A[9][23] * mat_B[23][14] +
                  mat_A[9][24] * mat_B[24][14] +
                  mat_A[9][25] * mat_B[25][14] +
                  mat_A[9][26] * mat_B[26][14] +
                  mat_A[9][27] * mat_B[27][14] +
                  mat_A[9][28] * mat_B[28][14] +
                  mat_A[9][29] * mat_B[29][14] +
                  mat_A[9][30] * mat_B[30][14] +
                  mat_A[9][31] * mat_B[31][14];
    mat_C[9][15] <= 
                  mat_A[9][0] * mat_B[0][15] +
                  mat_A[9][1] * mat_B[1][15] +
                  mat_A[9][2] * mat_B[2][15] +
                  mat_A[9][3] * mat_B[3][15] +
                  mat_A[9][4] * mat_B[4][15] +
                  mat_A[9][5] * mat_B[5][15] +
                  mat_A[9][6] * mat_B[6][15] +
                  mat_A[9][7] * mat_B[7][15] +
                  mat_A[9][8] * mat_B[8][15] +
                  mat_A[9][9] * mat_B[9][15] +
                  mat_A[9][10] * mat_B[10][15] +
                  mat_A[9][11] * mat_B[11][15] +
                  mat_A[9][12] * mat_B[12][15] +
                  mat_A[9][13] * mat_B[13][15] +
                  mat_A[9][14] * mat_B[14][15] +
                  mat_A[9][15] * mat_B[15][15] +
                  mat_A[9][16] * mat_B[16][15] +
                  mat_A[9][17] * mat_B[17][15] +
                  mat_A[9][18] * mat_B[18][15] +
                  mat_A[9][19] * mat_B[19][15] +
                  mat_A[9][20] * mat_B[20][15] +
                  mat_A[9][21] * mat_B[21][15] +
                  mat_A[9][22] * mat_B[22][15] +
                  mat_A[9][23] * mat_B[23][15] +
                  mat_A[9][24] * mat_B[24][15] +
                  mat_A[9][25] * mat_B[25][15] +
                  mat_A[9][26] * mat_B[26][15] +
                  mat_A[9][27] * mat_B[27][15] +
                  mat_A[9][28] * mat_B[28][15] +
                  mat_A[9][29] * mat_B[29][15] +
                  mat_A[9][30] * mat_B[30][15] +
                  mat_A[9][31] * mat_B[31][15];
    mat_C[9][16] <= 
                  mat_A[9][0] * mat_B[0][16] +
                  mat_A[9][1] * mat_B[1][16] +
                  mat_A[9][2] * mat_B[2][16] +
                  mat_A[9][3] * mat_B[3][16] +
                  mat_A[9][4] * mat_B[4][16] +
                  mat_A[9][5] * mat_B[5][16] +
                  mat_A[9][6] * mat_B[6][16] +
                  mat_A[9][7] * mat_B[7][16] +
                  mat_A[9][8] * mat_B[8][16] +
                  mat_A[9][9] * mat_B[9][16] +
                  mat_A[9][10] * mat_B[10][16] +
                  mat_A[9][11] * mat_B[11][16] +
                  mat_A[9][12] * mat_B[12][16] +
                  mat_A[9][13] * mat_B[13][16] +
                  mat_A[9][14] * mat_B[14][16] +
                  mat_A[9][15] * mat_B[15][16] +
                  mat_A[9][16] * mat_B[16][16] +
                  mat_A[9][17] * mat_B[17][16] +
                  mat_A[9][18] * mat_B[18][16] +
                  mat_A[9][19] * mat_B[19][16] +
                  mat_A[9][20] * mat_B[20][16] +
                  mat_A[9][21] * mat_B[21][16] +
                  mat_A[9][22] * mat_B[22][16] +
                  mat_A[9][23] * mat_B[23][16] +
                  mat_A[9][24] * mat_B[24][16] +
                  mat_A[9][25] * mat_B[25][16] +
                  mat_A[9][26] * mat_B[26][16] +
                  mat_A[9][27] * mat_B[27][16] +
                  mat_A[9][28] * mat_B[28][16] +
                  mat_A[9][29] * mat_B[29][16] +
                  mat_A[9][30] * mat_B[30][16] +
                  mat_A[9][31] * mat_B[31][16];
    mat_C[9][17] <= 
                  mat_A[9][0] * mat_B[0][17] +
                  mat_A[9][1] * mat_B[1][17] +
                  mat_A[9][2] * mat_B[2][17] +
                  mat_A[9][3] * mat_B[3][17] +
                  mat_A[9][4] * mat_B[4][17] +
                  mat_A[9][5] * mat_B[5][17] +
                  mat_A[9][6] * mat_B[6][17] +
                  mat_A[9][7] * mat_B[7][17] +
                  mat_A[9][8] * mat_B[8][17] +
                  mat_A[9][9] * mat_B[9][17] +
                  mat_A[9][10] * mat_B[10][17] +
                  mat_A[9][11] * mat_B[11][17] +
                  mat_A[9][12] * mat_B[12][17] +
                  mat_A[9][13] * mat_B[13][17] +
                  mat_A[9][14] * mat_B[14][17] +
                  mat_A[9][15] * mat_B[15][17] +
                  mat_A[9][16] * mat_B[16][17] +
                  mat_A[9][17] * mat_B[17][17] +
                  mat_A[9][18] * mat_B[18][17] +
                  mat_A[9][19] * mat_B[19][17] +
                  mat_A[9][20] * mat_B[20][17] +
                  mat_A[9][21] * mat_B[21][17] +
                  mat_A[9][22] * mat_B[22][17] +
                  mat_A[9][23] * mat_B[23][17] +
                  mat_A[9][24] * mat_B[24][17] +
                  mat_A[9][25] * mat_B[25][17] +
                  mat_A[9][26] * mat_B[26][17] +
                  mat_A[9][27] * mat_B[27][17] +
                  mat_A[9][28] * mat_B[28][17] +
                  mat_A[9][29] * mat_B[29][17] +
                  mat_A[9][30] * mat_B[30][17] +
                  mat_A[9][31] * mat_B[31][17];
    mat_C[9][18] <= 
                  mat_A[9][0] * mat_B[0][18] +
                  mat_A[9][1] * mat_B[1][18] +
                  mat_A[9][2] * mat_B[2][18] +
                  mat_A[9][3] * mat_B[3][18] +
                  mat_A[9][4] * mat_B[4][18] +
                  mat_A[9][5] * mat_B[5][18] +
                  mat_A[9][6] * mat_B[6][18] +
                  mat_A[9][7] * mat_B[7][18] +
                  mat_A[9][8] * mat_B[8][18] +
                  mat_A[9][9] * mat_B[9][18] +
                  mat_A[9][10] * mat_B[10][18] +
                  mat_A[9][11] * mat_B[11][18] +
                  mat_A[9][12] * mat_B[12][18] +
                  mat_A[9][13] * mat_B[13][18] +
                  mat_A[9][14] * mat_B[14][18] +
                  mat_A[9][15] * mat_B[15][18] +
                  mat_A[9][16] * mat_B[16][18] +
                  mat_A[9][17] * mat_B[17][18] +
                  mat_A[9][18] * mat_B[18][18] +
                  mat_A[9][19] * mat_B[19][18] +
                  mat_A[9][20] * mat_B[20][18] +
                  mat_A[9][21] * mat_B[21][18] +
                  mat_A[9][22] * mat_B[22][18] +
                  mat_A[9][23] * mat_B[23][18] +
                  mat_A[9][24] * mat_B[24][18] +
                  mat_A[9][25] * mat_B[25][18] +
                  mat_A[9][26] * mat_B[26][18] +
                  mat_A[9][27] * mat_B[27][18] +
                  mat_A[9][28] * mat_B[28][18] +
                  mat_A[9][29] * mat_B[29][18] +
                  mat_A[9][30] * mat_B[30][18] +
                  mat_A[9][31] * mat_B[31][18];
    mat_C[9][19] <= 
                  mat_A[9][0] * mat_B[0][19] +
                  mat_A[9][1] * mat_B[1][19] +
                  mat_A[9][2] * mat_B[2][19] +
                  mat_A[9][3] * mat_B[3][19] +
                  mat_A[9][4] * mat_B[4][19] +
                  mat_A[9][5] * mat_B[5][19] +
                  mat_A[9][6] * mat_B[6][19] +
                  mat_A[9][7] * mat_B[7][19] +
                  mat_A[9][8] * mat_B[8][19] +
                  mat_A[9][9] * mat_B[9][19] +
                  mat_A[9][10] * mat_B[10][19] +
                  mat_A[9][11] * mat_B[11][19] +
                  mat_A[9][12] * mat_B[12][19] +
                  mat_A[9][13] * mat_B[13][19] +
                  mat_A[9][14] * mat_B[14][19] +
                  mat_A[9][15] * mat_B[15][19] +
                  mat_A[9][16] * mat_B[16][19] +
                  mat_A[9][17] * mat_B[17][19] +
                  mat_A[9][18] * mat_B[18][19] +
                  mat_A[9][19] * mat_B[19][19] +
                  mat_A[9][20] * mat_B[20][19] +
                  mat_A[9][21] * mat_B[21][19] +
                  mat_A[9][22] * mat_B[22][19] +
                  mat_A[9][23] * mat_B[23][19] +
                  mat_A[9][24] * mat_B[24][19] +
                  mat_A[9][25] * mat_B[25][19] +
                  mat_A[9][26] * mat_B[26][19] +
                  mat_A[9][27] * mat_B[27][19] +
                  mat_A[9][28] * mat_B[28][19] +
                  mat_A[9][29] * mat_B[29][19] +
                  mat_A[9][30] * mat_B[30][19] +
                  mat_A[9][31] * mat_B[31][19];
    mat_C[9][20] <= 
                  mat_A[9][0] * mat_B[0][20] +
                  mat_A[9][1] * mat_B[1][20] +
                  mat_A[9][2] * mat_B[2][20] +
                  mat_A[9][3] * mat_B[3][20] +
                  mat_A[9][4] * mat_B[4][20] +
                  mat_A[9][5] * mat_B[5][20] +
                  mat_A[9][6] * mat_B[6][20] +
                  mat_A[9][7] * mat_B[7][20] +
                  mat_A[9][8] * mat_B[8][20] +
                  mat_A[9][9] * mat_B[9][20] +
                  mat_A[9][10] * mat_B[10][20] +
                  mat_A[9][11] * mat_B[11][20] +
                  mat_A[9][12] * mat_B[12][20] +
                  mat_A[9][13] * mat_B[13][20] +
                  mat_A[9][14] * mat_B[14][20] +
                  mat_A[9][15] * mat_B[15][20] +
                  mat_A[9][16] * mat_B[16][20] +
                  mat_A[9][17] * mat_B[17][20] +
                  mat_A[9][18] * mat_B[18][20] +
                  mat_A[9][19] * mat_B[19][20] +
                  mat_A[9][20] * mat_B[20][20] +
                  mat_A[9][21] * mat_B[21][20] +
                  mat_A[9][22] * mat_B[22][20] +
                  mat_A[9][23] * mat_B[23][20] +
                  mat_A[9][24] * mat_B[24][20] +
                  mat_A[9][25] * mat_B[25][20] +
                  mat_A[9][26] * mat_B[26][20] +
                  mat_A[9][27] * mat_B[27][20] +
                  mat_A[9][28] * mat_B[28][20] +
                  mat_A[9][29] * mat_B[29][20] +
                  mat_A[9][30] * mat_B[30][20] +
                  mat_A[9][31] * mat_B[31][20];
    mat_C[9][21] <= 
                  mat_A[9][0] * mat_B[0][21] +
                  mat_A[9][1] * mat_B[1][21] +
                  mat_A[9][2] * mat_B[2][21] +
                  mat_A[9][3] * mat_B[3][21] +
                  mat_A[9][4] * mat_B[4][21] +
                  mat_A[9][5] * mat_B[5][21] +
                  mat_A[9][6] * mat_B[6][21] +
                  mat_A[9][7] * mat_B[7][21] +
                  mat_A[9][8] * mat_B[8][21] +
                  mat_A[9][9] * mat_B[9][21] +
                  mat_A[9][10] * mat_B[10][21] +
                  mat_A[9][11] * mat_B[11][21] +
                  mat_A[9][12] * mat_B[12][21] +
                  mat_A[9][13] * mat_B[13][21] +
                  mat_A[9][14] * mat_B[14][21] +
                  mat_A[9][15] * mat_B[15][21] +
                  mat_A[9][16] * mat_B[16][21] +
                  mat_A[9][17] * mat_B[17][21] +
                  mat_A[9][18] * mat_B[18][21] +
                  mat_A[9][19] * mat_B[19][21] +
                  mat_A[9][20] * mat_B[20][21] +
                  mat_A[9][21] * mat_B[21][21] +
                  mat_A[9][22] * mat_B[22][21] +
                  mat_A[9][23] * mat_B[23][21] +
                  mat_A[9][24] * mat_B[24][21] +
                  mat_A[9][25] * mat_B[25][21] +
                  mat_A[9][26] * mat_B[26][21] +
                  mat_A[9][27] * mat_B[27][21] +
                  mat_A[9][28] * mat_B[28][21] +
                  mat_A[9][29] * mat_B[29][21] +
                  mat_A[9][30] * mat_B[30][21] +
                  mat_A[9][31] * mat_B[31][21];
    mat_C[9][22] <= 
                  mat_A[9][0] * mat_B[0][22] +
                  mat_A[9][1] * mat_B[1][22] +
                  mat_A[9][2] * mat_B[2][22] +
                  mat_A[9][3] * mat_B[3][22] +
                  mat_A[9][4] * mat_B[4][22] +
                  mat_A[9][5] * mat_B[5][22] +
                  mat_A[9][6] * mat_B[6][22] +
                  mat_A[9][7] * mat_B[7][22] +
                  mat_A[9][8] * mat_B[8][22] +
                  mat_A[9][9] * mat_B[9][22] +
                  mat_A[9][10] * mat_B[10][22] +
                  mat_A[9][11] * mat_B[11][22] +
                  mat_A[9][12] * mat_B[12][22] +
                  mat_A[9][13] * mat_B[13][22] +
                  mat_A[9][14] * mat_B[14][22] +
                  mat_A[9][15] * mat_B[15][22] +
                  mat_A[9][16] * mat_B[16][22] +
                  mat_A[9][17] * mat_B[17][22] +
                  mat_A[9][18] * mat_B[18][22] +
                  mat_A[9][19] * mat_B[19][22] +
                  mat_A[9][20] * mat_B[20][22] +
                  mat_A[9][21] * mat_B[21][22] +
                  mat_A[9][22] * mat_B[22][22] +
                  mat_A[9][23] * mat_B[23][22] +
                  mat_A[9][24] * mat_B[24][22] +
                  mat_A[9][25] * mat_B[25][22] +
                  mat_A[9][26] * mat_B[26][22] +
                  mat_A[9][27] * mat_B[27][22] +
                  mat_A[9][28] * mat_B[28][22] +
                  mat_A[9][29] * mat_B[29][22] +
                  mat_A[9][30] * mat_B[30][22] +
                  mat_A[9][31] * mat_B[31][22];
    mat_C[9][23] <= 
                  mat_A[9][0] * mat_B[0][23] +
                  mat_A[9][1] * mat_B[1][23] +
                  mat_A[9][2] * mat_B[2][23] +
                  mat_A[9][3] * mat_B[3][23] +
                  mat_A[9][4] * mat_B[4][23] +
                  mat_A[9][5] * mat_B[5][23] +
                  mat_A[9][6] * mat_B[6][23] +
                  mat_A[9][7] * mat_B[7][23] +
                  mat_A[9][8] * mat_B[8][23] +
                  mat_A[9][9] * mat_B[9][23] +
                  mat_A[9][10] * mat_B[10][23] +
                  mat_A[9][11] * mat_B[11][23] +
                  mat_A[9][12] * mat_B[12][23] +
                  mat_A[9][13] * mat_B[13][23] +
                  mat_A[9][14] * mat_B[14][23] +
                  mat_A[9][15] * mat_B[15][23] +
                  mat_A[9][16] * mat_B[16][23] +
                  mat_A[9][17] * mat_B[17][23] +
                  mat_A[9][18] * mat_B[18][23] +
                  mat_A[9][19] * mat_B[19][23] +
                  mat_A[9][20] * mat_B[20][23] +
                  mat_A[9][21] * mat_B[21][23] +
                  mat_A[9][22] * mat_B[22][23] +
                  mat_A[9][23] * mat_B[23][23] +
                  mat_A[9][24] * mat_B[24][23] +
                  mat_A[9][25] * mat_B[25][23] +
                  mat_A[9][26] * mat_B[26][23] +
                  mat_A[9][27] * mat_B[27][23] +
                  mat_A[9][28] * mat_B[28][23] +
                  mat_A[9][29] * mat_B[29][23] +
                  mat_A[9][30] * mat_B[30][23] +
                  mat_A[9][31] * mat_B[31][23];
    mat_C[9][24] <= 
                  mat_A[9][0] * mat_B[0][24] +
                  mat_A[9][1] * mat_B[1][24] +
                  mat_A[9][2] * mat_B[2][24] +
                  mat_A[9][3] * mat_B[3][24] +
                  mat_A[9][4] * mat_B[4][24] +
                  mat_A[9][5] * mat_B[5][24] +
                  mat_A[9][6] * mat_B[6][24] +
                  mat_A[9][7] * mat_B[7][24] +
                  mat_A[9][8] * mat_B[8][24] +
                  mat_A[9][9] * mat_B[9][24] +
                  mat_A[9][10] * mat_B[10][24] +
                  mat_A[9][11] * mat_B[11][24] +
                  mat_A[9][12] * mat_B[12][24] +
                  mat_A[9][13] * mat_B[13][24] +
                  mat_A[9][14] * mat_B[14][24] +
                  mat_A[9][15] * mat_B[15][24] +
                  mat_A[9][16] * mat_B[16][24] +
                  mat_A[9][17] * mat_B[17][24] +
                  mat_A[9][18] * mat_B[18][24] +
                  mat_A[9][19] * mat_B[19][24] +
                  mat_A[9][20] * mat_B[20][24] +
                  mat_A[9][21] * mat_B[21][24] +
                  mat_A[9][22] * mat_B[22][24] +
                  mat_A[9][23] * mat_B[23][24] +
                  mat_A[9][24] * mat_B[24][24] +
                  mat_A[9][25] * mat_B[25][24] +
                  mat_A[9][26] * mat_B[26][24] +
                  mat_A[9][27] * mat_B[27][24] +
                  mat_A[9][28] * mat_B[28][24] +
                  mat_A[9][29] * mat_B[29][24] +
                  mat_A[9][30] * mat_B[30][24] +
                  mat_A[9][31] * mat_B[31][24];
    mat_C[9][25] <= 
                  mat_A[9][0] * mat_B[0][25] +
                  mat_A[9][1] * mat_B[1][25] +
                  mat_A[9][2] * mat_B[2][25] +
                  mat_A[9][3] * mat_B[3][25] +
                  mat_A[9][4] * mat_B[4][25] +
                  mat_A[9][5] * mat_B[5][25] +
                  mat_A[9][6] * mat_B[6][25] +
                  mat_A[9][7] * mat_B[7][25] +
                  mat_A[9][8] * mat_B[8][25] +
                  mat_A[9][9] * mat_B[9][25] +
                  mat_A[9][10] * mat_B[10][25] +
                  mat_A[9][11] * mat_B[11][25] +
                  mat_A[9][12] * mat_B[12][25] +
                  mat_A[9][13] * mat_B[13][25] +
                  mat_A[9][14] * mat_B[14][25] +
                  mat_A[9][15] * mat_B[15][25] +
                  mat_A[9][16] * mat_B[16][25] +
                  mat_A[9][17] * mat_B[17][25] +
                  mat_A[9][18] * mat_B[18][25] +
                  mat_A[9][19] * mat_B[19][25] +
                  mat_A[9][20] * mat_B[20][25] +
                  mat_A[9][21] * mat_B[21][25] +
                  mat_A[9][22] * mat_B[22][25] +
                  mat_A[9][23] * mat_B[23][25] +
                  mat_A[9][24] * mat_B[24][25] +
                  mat_A[9][25] * mat_B[25][25] +
                  mat_A[9][26] * mat_B[26][25] +
                  mat_A[9][27] * mat_B[27][25] +
                  mat_A[9][28] * mat_B[28][25] +
                  mat_A[9][29] * mat_B[29][25] +
                  mat_A[9][30] * mat_B[30][25] +
                  mat_A[9][31] * mat_B[31][25];
    mat_C[9][26] <= 
                  mat_A[9][0] * mat_B[0][26] +
                  mat_A[9][1] * mat_B[1][26] +
                  mat_A[9][2] * mat_B[2][26] +
                  mat_A[9][3] * mat_B[3][26] +
                  mat_A[9][4] * mat_B[4][26] +
                  mat_A[9][5] * mat_B[5][26] +
                  mat_A[9][6] * mat_B[6][26] +
                  mat_A[9][7] * mat_B[7][26] +
                  mat_A[9][8] * mat_B[8][26] +
                  mat_A[9][9] * mat_B[9][26] +
                  mat_A[9][10] * mat_B[10][26] +
                  mat_A[9][11] * mat_B[11][26] +
                  mat_A[9][12] * mat_B[12][26] +
                  mat_A[9][13] * mat_B[13][26] +
                  mat_A[9][14] * mat_B[14][26] +
                  mat_A[9][15] * mat_B[15][26] +
                  mat_A[9][16] * mat_B[16][26] +
                  mat_A[9][17] * mat_B[17][26] +
                  mat_A[9][18] * mat_B[18][26] +
                  mat_A[9][19] * mat_B[19][26] +
                  mat_A[9][20] * mat_B[20][26] +
                  mat_A[9][21] * mat_B[21][26] +
                  mat_A[9][22] * mat_B[22][26] +
                  mat_A[9][23] * mat_B[23][26] +
                  mat_A[9][24] * mat_B[24][26] +
                  mat_A[9][25] * mat_B[25][26] +
                  mat_A[9][26] * mat_B[26][26] +
                  mat_A[9][27] * mat_B[27][26] +
                  mat_A[9][28] * mat_B[28][26] +
                  mat_A[9][29] * mat_B[29][26] +
                  mat_A[9][30] * mat_B[30][26] +
                  mat_A[9][31] * mat_B[31][26];
    mat_C[9][27] <= 
                  mat_A[9][0] * mat_B[0][27] +
                  mat_A[9][1] * mat_B[1][27] +
                  mat_A[9][2] * mat_B[2][27] +
                  mat_A[9][3] * mat_B[3][27] +
                  mat_A[9][4] * mat_B[4][27] +
                  mat_A[9][5] * mat_B[5][27] +
                  mat_A[9][6] * mat_B[6][27] +
                  mat_A[9][7] * mat_B[7][27] +
                  mat_A[9][8] * mat_B[8][27] +
                  mat_A[9][9] * mat_B[9][27] +
                  mat_A[9][10] * mat_B[10][27] +
                  mat_A[9][11] * mat_B[11][27] +
                  mat_A[9][12] * mat_B[12][27] +
                  mat_A[9][13] * mat_B[13][27] +
                  mat_A[9][14] * mat_B[14][27] +
                  mat_A[9][15] * mat_B[15][27] +
                  mat_A[9][16] * mat_B[16][27] +
                  mat_A[9][17] * mat_B[17][27] +
                  mat_A[9][18] * mat_B[18][27] +
                  mat_A[9][19] * mat_B[19][27] +
                  mat_A[9][20] * mat_B[20][27] +
                  mat_A[9][21] * mat_B[21][27] +
                  mat_A[9][22] * mat_B[22][27] +
                  mat_A[9][23] * mat_B[23][27] +
                  mat_A[9][24] * mat_B[24][27] +
                  mat_A[9][25] * mat_B[25][27] +
                  mat_A[9][26] * mat_B[26][27] +
                  mat_A[9][27] * mat_B[27][27] +
                  mat_A[9][28] * mat_B[28][27] +
                  mat_A[9][29] * mat_B[29][27] +
                  mat_A[9][30] * mat_B[30][27] +
                  mat_A[9][31] * mat_B[31][27];
    mat_C[9][28] <= 
                  mat_A[9][0] * mat_B[0][28] +
                  mat_A[9][1] * mat_B[1][28] +
                  mat_A[9][2] * mat_B[2][28] +
                  mat_A[9][3] * mat_B[3][28] +
                  mat_A[9][4] * mat_B[4][28] +
                  mat_A[9][5] * mat_B[5][28] +
                  mat_A[9][6] * mat_B[6][28] +
                  mat_A[9][7] * mat_B[7][28] +
                  mat_A[9][8] * mat_B[8][28] +
                  mat_A[9][9] * mat_B[9][28] +
                  mat_A[9][10] * mat_B[10][28] +
                  mat_A[9][11] * mat_B[11][28] +
                  mat_A[9][12] * mat_B[12][28] +
                  mat_A[9][13] * mat_B[13][28] +
                  mat_A[9][14] * mat_B[14][28] +
                  mat_A[9][15] * mat_B[15][28] +
                  mat_A[9][16] * mat_B[16][28] +
                  mat_A[9][17] * mat_B[17][28] +
                  mat_A[9][18] * mat_B[18][28] +
                  mat_A[9][19] * mat_B[19][28] +
                  mat_A[9][20] * mat_B[20][28] +
                  mat_A[9][21] * mat_B[21][28] +
                  mat_A[9][22] * mat_B[22][28] +
                  mat_A[9][23] * mat_B[23][28] +
                  mat_A[9][24] * mat_B[24][28] +
                  mat_A[9][25] * mat_B[25][28] +
                  mat_A[9][26] * mat_B[26][28] +
                  mat_A[9][27] * mat_B[27][28] +
                  mat_A[9][28] * mat_B[28][28] +
                  mat_A[9][29] * mat_B[29][28] +
                  mat_A[9][30] * mat_B[30][28] +
                  mat_A[9][31] * mat_B[31][28];
    mat_C[9][29] <= 
                  mat_A[9][0] * mat_B[0][29] +
                  mat_A[9][1] * mat_B[1][29] +
                  mat_A[9][2] * mat_B[2][29] +
                  mat_A[9][3] * mat_B[3][29] +
                  mat_A[9][4] * mat_B[4][29] +
                  mat_A[9][5] * mat_B[5][29] +
                  mat_A[9][6] * mat_B[6][29] +
                  mat_A[9][7] * mat_B[7][29] +
                  mat_A[9][8] * mat_B[8][29] +
                  mat_A[9][9] * mat_B[9][29] +
                  mat_A[9][10] * mat_B[10][29] +
                  mat_A[9][11] * mat_B[11][29] +
                  mat_A[9][12] * mat_B[12][29] +
                  mat_A[9][13] * mat_B[13][29] +
                  mat_A[9][14] * mat_B[14][29] +
                  mat_A[9][15] * mat_B[15][29] +
                  mat_A[9][16] * mat_B[16][29] +
                  mat_A[9][17] * mat_B[17][29] +
                  mat_A[9][18] * mat_B[18][29] +
                  mat_A[9][19] * mat_B[19][29] +
                  mat_A[9][20] * mat_B[20][29] +
                  mat_A[9][21] * mat_B[21][29] +
                  mat_A[9][22] * mat_B[22][29] +
                  mat_A[9][23] * mat_B[23][29] +
                  mat_A[9][24] * mat_B[24][29] +
                  mat_A[9][25] * mat_B[25][29] +
                  mat_A[9][26] * mat_B[26][29] +
                  mat_A[9][27] * mat_B[27][29] +
                  mat_A[9][28] * mat_B[28][29] +
                  mat_A[9][29] * mat_B[29][29] +
                  mat_A[9][30] * mat_B[30][29] +
                  mat_A[9][31] * mat_B[31][29];
    mat_C[9][30] <= 
                  mat_A[9][0] * mat_B[0][30] +
                  mat_A[9][1] * mat_B[1][30] +
                  mat_A[9][2] * mat_B[2][30] +
                  mat_A[9][3] * mat_B[3][30] +
                  mat_A[9][4] * mat_B[4][30] +
                  mat_A[9][5] * mat_B[5][30] +
                  mat_A[9][6] * mat_B[6][30] +
                  mat_A[9][7] * mat_B[7][30] +
                  mat_A[9][8] * mat_B[8][30] +
                  mat_A[9][9] * mat_B[9][30] +
                  mat_A[9][10] * mat_B[10][30] +
                  mat_A[9][11] * mat_B[11][30] +
                  mat_A[9][12] * mat_B[12][30] +
                  mat_A[9][13] * mat_B[13][30] +
                  mat_A[9][14] * mat_B[14][30] +
                  mat_A[9][15] * mat_B[15][30] +
                  mat_A[9][16] * mat_B[16][30] +
                  mat_A[9][17] * mat_B[17][30] +
                  mat_A[9][18] * mat_B[18][30] +
                  mat_A[9][19] * mat_B[19][30] +
                  mat_A[9][20] * mat_B[20][30] +
                  mat_A[9][21] * mat_B[21][30] +
                  mat_A[9][22] * mat_B[22][30] +
                  mat_A[9][23] * mat_B[23][30] +
                  mat_A[9][24] * mat_B[24][30] +
                  mat_A[9][25] * mat_B[25][30] +
                  mat_A[9][26] * mat_B[26][30] +
                  mat_A[9][27] * mat_B[27][30] +
                  mat_A[9][28] * mat_B[28][30] +
                  mat_A[9][29] * mat_B[29][30] +
                  mat_A[9][30] * mat_B[30][30] +
                  mat_A[9][31] * mat_B[31][30];
    mat_C[9][31] <= 
                  mat_A[9][0] * mat_B[0][31] +
                  mat_A[9][1] * mat_B[1][31] +
                  mat_A[9][2] * mat_B[2][31] +
                  mat_A[9][3] * mat_B[3][31] +
                  mat_A[9][4] * mat_B[4][31] +
                  mat_A[9][5] * mat_B[5][31] +
                  mat_A[9][6] * mat_B[6][31] +
                  mat_A[9][7] * mat_B[7][31] +
                  mat_A[9][8] * mat_B[8][31] +
                  mat_A[9][9] * mat_B[9][31] +
                  mat_A[9][10] * mat_B[10][31] +
                  mat_A[9][11] * mat_B[11][31] +
                  mat_A[9][12] * mat_B[12][31] +
                  mat_A[9][13] * mat_B[13][31] +
                  mat_A[9][14] * mat_B[14][31] +
                  mat_A[9][15] * mat_B[15][31] +
                  mat_A[9][16] * mat_B[16][31] +
                  mat_A[9][17] * mat_B[17][31] +
                  mat_A[9][18] * mat_B[18][31] +
                  mat_A[9][19] * mat_B[19][31] +
                  mat_A[9][20] * mat_B[20][31] +
                  mat_A[9][21] * mat_B[21][31] +
                  mat_A[9][22] * mat_B[22][31] +
                  mat_A[9][23] * mat_B[23][31] +
                  mat_A[9][24] * mat_B[24][31] +
                  mat_A[9][25] * mat_B[25][31] +
                  mat_A[9][26] * mat_B[26][31] +
                  mat_A[9][27] * mat_B[27][31] +
                  mat_A[9][28] * mat_B[28][31] +
                  mat_A[9][29] * mat_B[29][31] +
                  mat_A[9][30] * mat_B[30][31] +
                  mat_A[9][31] * mat_B[31][31];
    mat_C[10][0] <= 
                  mat_A[10][0] * mat_B[0][0] +
                  mat_A[10][1] * mat_B[1][0] +
                  mat_A[10][2] * mat_B[2][0] +
                  mat_A[10][3] * mat_B[3][0] +
                  mat_A[10][4] * mat_B[4][0] +
                  mat_A[10][5] * mat_B[5][0] +
                  mat_A[10][6] * mat_B[6][0] +
                  mat_A[10][7] * mat_B[7][0] +
                  mat_A[10][8] * mat_B[8][0] +
                  mat_A[10][9] * mat_B[9][0] +
                  mat_A[10][10] * mat_B[10][0] +
                  mat_A[10][11] * mat_B[11][0] +
                  mat_A[10][12] * mat_B[12][0] +
                  mat_A[10][13] * mat_B[13][0] +
                  mat_A[10][14] * mat_B[14][0] +
                  mat_A[10][15] * mat_B[15][0] +
                  mat_A[10][16] * mat_B[16][0] +
                  mat_A[10][17] * mat_B[17][0] +
                  mat_A[10][18] * mat_B[18][0] +
                  mat_A[10][19] * mat_B[19][0] +
                  mat_A[10][20] * mat_B[20][0] +
                  mat_A[10][21] * mat_B[21][0] +
                  mat_A[10][22] * mat_B[22][0] +
                  mat_A[10][23] * mat_B[23][0] +
                  mat_A[10][24] * mat_B[24][0] +
                  mat_A[10][25] * mat_B[25][0] +
                  mat_A[10][26] * mat_B[26][0] +
                  mat_A[10][27] * mat_B[27][0] +
                  mat_A[10][28] * mat_B[28][0] +
                  mat_A[10][29] * mat_B[29][0] +
                  mat_A[10][30] * mat_B[30][0] +
                  mat_A[10][31] * mat_B[31][0];
    mat_C[10][1] <= 
                  mat_A[10][0] * mat_B[0][1] +
                  mat_A[10][1] * mat_B[1][1] +
                  mat_A[10][2] * mat_B[2][1] +
                  mat_A[10][3] * mat_B[3][1] +
                  mat_A[10][4] * mat_B[4][1] +
                  mat_A[10][5] * mat_B[5][1] +
                  mat_A[10][6] * mat_B[6][1] +
                  mat_A[10][7] * mat_B[7][1] +
                  mat_A[10][8] * mat_B[8][1] +
                  mat_A[10][9] * mat_B[9][1] +
                  mat_A[10][10] * mat_B[10][1] +
                  mat_A[10][11] * mat_B[11][1] +
                  mat_A[10][12] * mat_B[12][1] +
                  mat_A[10][13] * mat_B[13][1] +
                  mat_A[10][14] * mat_B[14][1] +
                  mat_A[10][15] * mat_B[15][1] +
                  mat_A[10][16] * mat_B[16][1] +
                  mat_A[10][17] * mat_B[17][1] +
                  mat_A[10][18] * mat_B[18][1] +
                  mat_A[10][19] * mat_B[19][1] +
                  mat_A[10][20] * mat_B[20][1] +
                  mat_A[10][21] * mat_B[21][1] +
                  mat_A[10][22] * mat_B[22][1] +
                  mat_A[10][23] * mat_B[23][1] +
                  mat_A[10][24] * mat_B[24][1] +
                  mat_A[10][25] * mat_B[25][1] +
                  mat_A[10][26] * mat_B[26][1] +
                  mat_A[10][27] * mat_B[27][1] +
                  mat_A[10][28] * mat_B[28][1] +
                  mat_A[10][29] * mat_B[29][1] +
                  mat_A[10][30] * mat_B[30][1] +
                  mat_A[10][31] * mat_B[31][1];
    mat_C[10][2] <= 
                  mat_A[10][0] * mat_B[0][2] +
                  mat_A[10][1] * mat_B[1][2] +
                  mat_A[10][2] * mat_B[2][2] +
                  mat_A[10][3] * mat_B[3][2] +
                  mat_A[10][4] * mat_B[4][2] +
                  mat_A[10][5] * mat_B[5][2] +
                  mat_A[10][6] * mat_B[6][2] +
                  mat_A[10][7] * mat_B[7][2] +
                  mat_A[10][8] * mat_B[8][2] +
                  mat_A[10][9] * mat_B[9][2] +
                  mat_A[10][10] * mat_B[10][2] +
                  mat_A[10][11] * mat_B[11][2] +
                  mat_A[10][12] * mat_B[12][2] +
                  mat_A[10][13] * mat_B[13][2] +
                  mat_A[10][14] * mat_B[14][2] +
                  mat_A[10][15] * mat_B[15][2] +
                  mat_A[10][16] * mat_B[16][2] +
                  mat_A[10][17] * mat_B[17][2] +
                  mat_A[10][18] * mat_B[18][2] +
                  mat_A[10][19] * mat_B[19][2] +
                  mat_A[10][20] * mat_B[20][2] +
                  mat_A[10][21] * mat_B[21][2] +
                  mat_A[10][22] * mat_B[22][2] +
                  mat_A[10][23] * mat_B[23][2] +
                  mat_A[10][24] * mat_B[24][2] +
                  mat_A[10][25] * mat_B[25][2] +
                  mat_A[10][26] * mat_B[26][2] +
                  mat_A[10][27] * mat_B[27][2] +
                  mat_A[10][28] * mat_B[28][2] +
                  mat_A[10][29] * mat_B[29][2] +
                  mat_A[10][30] * mat_B[30][2] +
                  mat_A[10][31] * mat_B[31][2];
    mat_C[10][3] <= 
                  mat_A[10][0] * mat_B[0][3] +
                  mat_A[10][1] * mat_B[1][3] +
                  mat_A[10][2] * mat_B[2][3] +
                  mat_A[10][3] * mat_B[3][3] +
                  mat_A[10][4] * mat_B[4][3] +
                  mat_A[10][5] * mat_B[5][3] +
                  mat_A[10][6] * mat_B[6][3] +
                  mat_A[10][7] * mat_B[7][3] +
                  mat_A[10][8] * mat_B[8][3] +
                  mat_A[10][9] * mat_B[9][3] +
                  mat_A[10][10] * mat_B[10][3] +
                  mat_A[10][11] * mat_B[11][3] +
                  mat_A[10][12] * mat_B[12][3] +
                  mat_A[10][13] * mat_B[13][3] +
                  mat_A[10][14] * mat_B[14][3] +
                  mat_A[10][15] * mat_B[15][3] +
                  mat_A[10][16] * mat_B[16][3] +
                  mat_A[10][17] * mat_B[17][3] +
                  mat_A[10][18] * mat_B[18][3] +
                  mat_A[10][19] * mat_B[19][3] +
                  mat_A[10][20] * mat_B[20][3] +
                  mat_A[10][21] * mat_B[21][3] +
                  mat_A[10][22] * mat_B[22][3] +
                  mat_A[10][23] * mat_B[23][3] +
                  mat_A[10][24] * mat_B[24][3] +
                  mat_A[10][25] * mat_B[25][3] +
                  mat_A[10][26] * mat_B[26][3] +
                  mat_A[10][27] * mat_B[27][3] +
                  mat_A[10][28] * mat_B[28][3] +
                  mat_A[10][29] * mat_B[29][3] +
                  mat_A[10][30] * mat_B[30][3] +
                  mat_A[10][31] * mat_B[31][3];
    mat_C[10][4] <= 
                  mat_A[10][0] * mat_B[0][4] +
                  mat_A[10][1] * mat_B[1][4] +
                  mat_A[10][2] * mat_B[2][4] +
                  mat_A[10][3] * mat_B[3][4] +
                  mat_A[10][4] * mat_B[4][4] +
                  mat_A[10][5] * mat_B[5][4] +
                  mat_A[10][6] * mat_B[6][4] +
                  mat_A[10][7] * mat_B[7][4] +
                  mat_A[10][8] * mat_B[8][4] +
                  mat_A[10][9] * mat_B[9][4] +
                  mat_A[10][10] * mat_B[10][4] +
                  mat_A[10][11] * mat_B[11][4] +
                  mat_A[10][12] * mat_B[12][4] +
                  mat_A[10][13] * mat_B[13][4] +
                  mat_A[10][14] * mat_B[14][4] +
                  mat_A[10][15] * mat_B[15][4] +
                  mat_A[10][16] * mat_B[16][4] +
                  mat_A[10][17] * mat_B[17][4] +
                  mat_A[10][18] * mat_B[18][4] +
                  mat_A[10][19] * mat_B[19][4] +
                  mat_A[10][20] * mat_B[20][4] +
                  mat_A[10][21] * mat_B[21][4] +
                  mat_A[10][22] * mat_B[22][4] +
                  mat_A[10][23] * mat_B[23][4] +
                  mat_A[10][24] * mat_B[24][4] +
                  mat_A[10][25] * mat_B[25][4] +
                  mat_A[10][26] * mat_B[26][4] +
                  mat_A[10][27] * mat_B[27][4] +
                  mat_A[10][28] * mat_B[28][4] +
                  mat_A[10][29] * mat_B[29][4] +
                  mat_A[10][30] * mat_B[30][4] +
                  mat_A[10][31] * mat_B[31][4];
    mat_C[10][5] <= 
                  mat_A[10][0] * mat_B[0][5] +
                  mat_A[10][1] * mat_B[1][5] +
                  mat_A[10][2] * mat_B[2][5] +
                  mat_A[10][3] * mat_B[3][5] +
                  mat_A[10][4] * mat_B[4][5] +
                  mat_A[10][5] * mat_B[5][5] +
                  mat_A[10][6] * mat_B[6][5] +
                  mat_A[10][7] * mat_B[7][5] +
                  mat_A[10][8] * mat_B[8][5] +
                  mat_A[10][9] * mat_B[9][5] +
                  mat_A[10][10] * mat_B[10][5] +
                  mat_A[10][11] * mat_B[11][5] +
                  mat_A[10][12] * mat_B[12][5] +
                  mat_A[10][13] * mat_B[13][5] +
                  mat_A[10][14] * mat_B[14][5] +
                  mat_A[10][15] * mat_B[15][5] +
                  mat_A[10][16] * mat_B[16][5] +
                  mat_A[10][17] * mat_B[17][5] +
                  mat_A[10][18] * mat_B[18][5] +
                  mat_A[10][19] * mat_B[19][5] +
                  mat_A[10][20] * mat_B[20][5] +
                  mat_A[10][21] * mat_B[21][5] +
                  mat_A[10][22] * mat_B[22][5] +
                  mat_A[10][23] * mat_B[23][5] +
                  mat_A[10][24] * mat_B[24][5] +
                  mat_A[10][25] * mat_B[25][5] +
                  mat_A[10][26] * mat_B[26][5] +
                  mat_A[10][27] * mat_B[27][5] +
                  mat_A[10][28] * mat_B[28][5] +
                  mat_A[10][29] * mat_B[29][5] +
                  mat_A[10][30] * mat_B[30][5] +
                  mat_A[10][31] * mat_B[31][5];
    mat_C[10][6] <= 
                  mat_A[10][0] * mat_B[0][6] +
                  mat_A[10][1] * mat_B[1][6] +
                  mat_A[10][2] * mat_B[2][6] +
                  mat_A[10][3] * mat_B[3][6] +
                  mat_A[10][4] * mat_B[4][6] +
                  mat_A[10][5] * mat_B[5][6] +
                  mat_A[10][6] * mat_B[6][6] +
                  mat_A[10][7] * mat_B[7][6] +
                  mat_A[10][8] * mat_B[8][6] +
                  mat_A[10][9] * mat_B[9][6] +
                  mat_A[10][10] * mat_B[10][6] +
                  mat_A[10][11] * mat_B[11][6] +
                  mat_A[10][12] * mat_B[12][6] +
                  mat_A[10][13] * mat_B[13][6] +
                  mat_A[10][14] * mat_B[14][6] +
                  mat_A[10][15] * mat_B[15][6] +
                  mat_A[10][16] * mat_B[16][6] +
                  mat_A[10][17] * mat_B[17][6] +
                  mat_A[10][18] * mat_B[18][6] +
                  mat_A[10][19] * mat_B[19][6] +
                  mat_A[10][20] * mat_B[20][6] +
                  mat_A[10][21] * mat_B[21][6] +
                  mat_A[10][22] * mat_B[22][6] +
                  mat_A[10][23] * mat_B[23][6] +
                  mat_A[10][24] * mat_B[24][6] +
                  mat_A[10][25] * mat_B[25][6] +
                  mat_A[10][26] * mat_B[26][6] +
                  mat_A[10][27] * mat_B[27][6] +
                  mat_A[10][28] * mat_B[28][6] +
                  mat_A[10][29] * mat_B[29][6] +
                  mat_A[10][30] * mat_B[30][6] +
                  mat_A[10][31] * mat_B[31][6];
    mat_C[10][7] <= 
                  mat_A[10][0] * mat_B[0][7] +
                  mat_A[10][1] * mat_B[1][7] +
                  mat_A[10][2] * mat_B[2][7] +
                  mat_A[10][3] * mat_B[3][7] +
                  mat_A[10][4] * mat_B[4][7] +
                  mat_A[10][5] * mat_B[5][7] +
                  mat_A[10][6] * mat_B[6][7] +
                  mat_A[10][7] * mat_B[7][7] +
                  mat_A[10][8] * mat_B[8][7] +
                  mat_A[10][9] * mat_B[9][7] +
                  mat_A[10][10] * mat_B[10][7] +
                  mat_A[10][11] * mat_B[11][7] +
                  mat_A[10][12] * mat_B[12][7] +
                  mat_A[10][13] * mat_B[13][7] +
                  mat_A[10][14] * mat_B[14][7] +
                  mat_A[10][15] * mat_B[15][7] +
                  mat_A[10][16] * mat_B[16][7] +
                  mat_A[10][17] * mat_B[17][7] +
                  mat_A[10][18] * mat_B[18][7] +
                  mat_A[10][19] * mat_B[19][7] +
                  mat_A[10][20] * mat_B[20][7] +
                  mat_A[10][21] * mat_B[21][7] +
                  mat_A[10][22] * mat_B[22][7] +
                  mat_A[10][23] * mat_B[23][7] +
                  mat_A[10][24] * mat_B[24][7] +
                  mat_A[10][25] * mat_B[25][7] +
                  mat_A[10][26] * mat_B[26][7] +
                  mat_A[10][27] * mat_B[27][7] +
                  mat_A[10][28] * mat_B[28][7] +
                  mat_A[10][29] * mat_B[29][7] +
                  mat_A[10][30] * mat_B[30][7] +
                  mat_A[10][31] * mat_B[31][7];
    mat_C[10][8] <= 
                  mat_A[10][0] * mat_B[0][8] +
                  mat_A[10][1] * mat_B[1][8] +
                  mat_A[10][2] * mat_B[2][8] +
                  mat_A[10][3] * mat_B[3][8] +
                  mat_A[10][4] * mat_B[4][8] +
                  mat_A[10][5] * mat_B[5][8] +
                  mat_A[10][6] * mat_B[6][8] +
                  mat_A[10][7] * mat_B[7][8] +
                  mat_A[10][8] * mat_B[8][8] +
                  mat_A[10][9] * mat_B[9][8] +
                  mat_A[10][10] * mat_B[10][8] +
                  mat_A[10][11] * mat_B[11][8] +
                  mat_A[10][12] * mat_B[12][8] +
                  mat_A[10][13] * mat_B[13][8] +
                  mat_A[10][14] * mat_B[14][8] +
                  mat_A[10][15] * mat_B[15][8] +
                  mat_A[10][16] * mat_B[16][8] +
                  mat_A[10][17] * mat_B[17][8] +
                  mat_A[10][18] * mat_B[18][8] +
                  mat_A[10][19] * mat_B[19][8] +
                  mat_A[10][20] * mat_B[20][8] +
                  mat_A[10][21] * mat_B[21][8] +
                  mat_A[10][22] * mat_B[22][8] +
                  mat_A[10][23] * mat_B[23][8] +
                  mat_A[10][24] * mat_B[24][8] +
                  mat_A[10][25] * mat_B[25][8] +
                  mat_A[10][26] * mat_B[26][8] +
                  mat_A[10][27] * mat_B[27][8] +
                  mat_A[10][28] * mat_B[28][8] +
                  mat_A[10][29] * mat_B[29][8] +
                  mat_A[10][30] * mat_B[30][8] +
                  mat_A[10][31] * mat_B[31][8];
    mat_C[10][9] <= 
                  mat_A[10][0] * mat_B[0][9] +
                  mat_A[10][1] * mat_B[1][9] +
                  mat_A[10][2] * mat_B[2][9] +
                  mat_A[10][3] * mat_B[3][9] +
                  mat_A[10][4] * mat_B[4][9] +
                  mat_A[10][5] * mat_B[5][9] +
                  mat_A[10][6] * mat_B[6][9] +
                  mat_A[10][7] * mat_B[7][9] +
                  mat_A[10][8] * mat_B[8][9] +
                  mat_A[10][9] * mat_B[9][9] +
                  mat_A[10][10] * mat_B[10][9] +
                  mat_A[10][11] * mat_B[11][9] +
                  mat_A[10][12] * mat_B[12][9] +
                  mat_A[10][13] * mat_B[13][9] +
                  mat_A[10][14] * mat_B[14][9] +
                  mat_A[10][15] * mat_B[15][9] +
                  mat_A[10][16] * mat_B[16][9] +
                  mat_A[10][17] * mat_B[17][9] +
                  mat_A[10][18] * mat_B[18][9] +
                  mat_A[10][19] * mat_B[19][9] +
                  mat_A[10][20] * mat_B[20][9] +
                  mat_A[10][21] * mat_B[21][9] +
                  mat_A[10][22] * mat_B[22][9] +
                  mat_A[10][23] * mat_B[23][9] +
                  mat_A[10][24] * mat_B[24][9] +
                  mat_A[10][25] * mat_B[25][9] +
                  mat_A[10][26] * mat_B[26][9] +
                  mat_A[10][27] * mat_B[27][9] +
                  mat_A[10][28] * mat_B[28][9] +
                  mat_A[10][29] * mat_B[29][9] +
                  mat_A[10][30] * mat_B[30][9] +
                  mat_A[10][31] * mat_B[31][9];
    mat_C[10][10] <= 
                  mat_A[10][0] * mat_B[0][10] +
                  mat_A[10][1] * mat_B[1][10] +
                  mat_A[10][2] * mat_B[2][10] +
                  mat_A[10][3] * mat_B[3][10] +
                  mat_A[10][4] * mat_B[4][10] +
                  mat_A[10][5] * mat_B[5][10] +
                  mat_A[10][6] * mat_B[6][10] +
                  mat_A[10][7] * mat_B[7][10] +
                  mat_A[10][8] * mat_B[8][10] +
                  mat_A[10][9] * mat_B[9][10] +
                  mat_A[10][10] * mat_B[10][10] +
                  mat_A[10][11] * mat_B[11][10] +
                  mat_A[10][12] * mat_B[12][10] +
                  mat_A[10][13] * mat_B[13][10] +
                  mat_A[10][14] * mat_B[14][10] +
                  mat_A[10][15] * mat_B[15][10] +
                  mat_A[10][16] * mat_B[16][10] +
                  mat_A[10][17] * mat_B[17][10] +
                  mat_A[10][18] * mat_B[18][10] +
                  mat_A[10][19] * mat_B[19][10] +
                  mat_A[10][20] * mat_B[20][10] +
                  mat_A[10][21] * mat_B[21][10] +
                  mat_A[10][22] * mat_B[22][10] +
                  mat_A[10][23] * mat_B[23][10] +
                  mat_A[10][24] * mat_B[24][10] +
                  mat_A[10][25] * mat_B[25][10] +
                  mat_A[10][26] * mat_B[26][10] +
                  mat_A[10][27] * mat_B[27][10] +
                  mat_A[10][28] * mat_B[28][10] +
                  mat_A[10][29] * mat_B[29][10] +
                  mat_A[10][30] * mat_B[30][10] +
                  mat_A[10][31] * mat_B[31][10];
    mat_C[10][11] <= 
                  mat_A[10][0] * mat_B[0][11] +
                  mat_A[10][1] * mat_B[1][11] +
                  mat_A[10][2] * mat_B[2][11] +
                  mat_A[10][3] * mat_B[3][11] +
                  mat_A[10][4] * mat_B[4][11] +
                  mat_A[10][5] * mat_B[5][11] +
                  mat_A[10][6] * mat_B[6][11] +
                  mat_A[10][7] * mat_B[7][11] +
                  mat_A[10][8] * mat_B[8][11] +
                  mat_A[10][9] * mat_B[9][11] +
                  mat_A[10][10] * mat_B[10][11] +
                  mat_A[10][11] * mat_B[11][11] +
                  mat_A[10][12] * mat_B[12][11] +
                  mat_A[10][13] * mat_B[13][11] +
                  mat_A[10][14] * mat_B[14][11] +
                  mat_A[10][15] * mat_B[15][11] +
                  mat_A[10][16] * mat_B[16][11] +
                  mat_A[10][17] * mat_B[17][11] +
                  mat_A[10][18] * mat_B[18][11] +
                  mat_A[10][19] * mat_B[19][11] +
                  mat_A[10][20] * mat_B[20][11] +
                  mat_A[10][21] * mat_B[21][11] +
                  mat_A[10][22] * mat_B[22][11] +
                  mat_A[10][23] * mat_B[23][11] +
                  mat_A[10][24] * mat_B[24][11] +
                  mat_A[10][25] * mat_B[25][11] +
                  mat_A[10][26] * mat_B[26][11] +
                  mat_A[10][27] * mat_B[27][11] +
                  mat_A[10][28] * mat_B[28][11] +
                  mat_A[10][29] * mat_B[29][11] +
                  mat_A[10][30] * mat_B[30][11] +
                  mat_A[10][31] * mat_B[31][11];
    mat_C[10][12] <= 
                  mat_A[10][0] * mat_B[0][12] +
                  mat_A[10][1] * mat_B[1][12] +
                  mat_A[10][2] * mat_B[2][12] +
                  mat_A[10][3] * mat_B[3][12] +
                  mat_A[10][4] * mat_B[4][12] +
                  mat_A[10][5] * mat_B[5][12] +
                  mat_A[10][6] * mat_B[6][12] +
                  mat_A[10][7] * mat_B[7][12] +
                  mat_A[10][8] * mat_B[8][12] +
                  mat_A[10][9] * mat_B[9][12] +
                  mat_A[10][10] * mat_B[10][12] +
                  mat_A[10][11] * mat_B[11][12] +
                  mat_A[10][12] * mat_B[12][12] +
                  mat_A[10][13] * mat_B[13][12] +
                  mat_A[10][14] * mat_B[14][12] +
                  mat_A[10][15] * mat_B[15][12] +
                  mat_A[10][16] * mat_B[16][12] +
                  mat_A[10][17] * mat_B[17][12] +
                  mat_A[10][18] * mat_B[18][12] +
                  mat_A[10][19] * mat_B[19][12] +
                  mat_A[10][20] * mat_B[20][12] +
                  mat_A[10][21] * mat_B[21][12] +
                  mat_A[10][22] * mat_B[22][12] +
                  mat_A[10][23] * mat_B[23][12] +
                  mat_A[10][24] * mat_B[24][12] +
                  mat_A[10][25] * mat_B[25][12] +
                  mat_A[10][26] * mat_B[26][12] +
                  mat_A[10][27] * mat_B[27][12] +
                  mat_A[10][28] * mat_B[28][12] +
                  mat_A[10][29] * mat_B[29][12] +
                  mat_A[10][30] * mat_B[30][12] +
                  mat_A[10][31] * mat_B[31][12];
    mat_C[10][13] <= 
                  mat_A[10][0] * mat_B[0][13] +
                  mat_A[10][1] * mat_B[1][13] +
                  mat_A[10][2] * mat_B[2][13] +
                  mat_A[10][3] * mat_B[3][13] +
                  mat_A[10][4] * mat_B[4][13] +
                  mat_A[10][5] * mat_B[5][13] +
                  mat_A[10][6] * mat_B[6][13] +
                  mat_A[10][7] * mat_B[7][13] +
                  mat_A[10][8] * mat_B[8][13] +
                  mat_A[10][9] * mat_B[9][13] +
                  mat_A[10][10] * mat_B[10][13] +
                  mat_A[10][11] * mat_B[11][13] +
                  mat_A[10][12] * mat_B[12][13] +
                  mat_A[10][13] * mat_B[13][13] +
                  mat_A[10][14] * mat_B[14][13] +
                  mat_A[10][15] * mat_B[15][13] +
                  mat_A[10][16] * mat_B[16][13] +
                  mat_A[10][17] * mat_B[17][13] +
                  mat_A[10][18] * mat_B[18][13] +
                  mat_A[10][19] * mat_B[19][13] +
                  mat_A[10][20] * mat_B[20][13] +
                  mat_A[10][21] * mat_B[21][13] +
                  mat_A[10][22] * mat_B[22][13] +
                  mat_A[10][23] * mat_B[23][13] +
                  mat_A[10][24] * mat_B[24][13] +
                  mat_A[10][25] * mat_B[25][13] +
                  mat_A[10][26] * mat_B[26][13] +
                  mat_A[10][27] * mat_B[27][13] +
                  mat_A[10][28] * mat_B[28][13] +
                  mat_A[10][29] * mat_B[29][13] +
                  mat_A[10][30] * mat_B[30][13] +
                  mat_A[10][31] * mat_B[31][13];
    mat_C[10][14] <= 
                  mat_A[10][0] * mat_B[0][14] +
                  mat_A[10][1] * mat_B[1][14] +
                  mat_A[10][2] * mat_B[2][14] +
                  mat_A[10][3] * mat_B[3][14] +
                  mat_A[10][4] * mat_B[4][14] +
                  mat_A[10][5] * mat_B[5][14] +
                  mat_A[10][6] * mat_B[6][14] +
                  mat_A[10][7] * mat_B[7][14] +
                  mat_A[10][8] * mat_B[8][14] +
                  mat_A[10][9] * mat_B[9][14] +
                  mat_A[10][10] * mat_B[10][14] +
                  mat_A[10][11] * mat_B[11][14] +
                  mat_A[10][12] * mat_B[12][14] +
                  mat_A[10][13] * mat_B[13][14] +
                  mat_A[10][14] * mat_B[14][14] +
                  mat_A[10][15] * mat_B[15][14] +
                  mat_A[10][16] * mat_B[16][14] +
                  mat_A[10][17] * mat_B[17][14] +
                  mat_A[10][18] * mat_B[18][14] +
                  mat_A[10][19] * mat_B[19][14] +
                  mat_A[10][20] * mat_B[20][14] +
                  mat_A[10][21] * mat_B[21][14] +
                  mat_A[10][22] * mat_B[22][14] +
                  mat_A[10][23] * mat_B[23][14] +
                  mat_A[10][24] * mat_B[24][14] +
                  mat_A[10][25] * mat_B[25][14] +
                  mat_A[10][26] * mat_B[26][14] +
                  mat_A[10][27] * mat_B[27][14] +
                  mat_A[10][28] * mat_B[28][14] +
                  mat_A[10][29] * mat_B[29][14] +
                  mat_A[10][30] * mat_B[30][14] +
                  mat_A[10][31] * mat_B[31][14];
    mat_C[10][15] <= 
                  mat_A[10][0] * mat_B[0][15] +
                  mat_A[10][1] * mat_B[1][15] +
                  mat_A[10][2] * mat_B[2][15] +
                  mat_A[10][3] * mat_B[3][15] +
                  mat_A[10][4] * mat_B[4][15] +
                  mat_A[10][5] * mat_B[5][15] +
                  mat_A[10][6] * mat_B[6][15] +
                  mat_A[10][7] * mat_B[7][15] +
                  mat_A[10][8] * mat_B[8][15] +
                  mat_A[10][9] * mat_B[9][15] +
                  mat_A[10][10] * mat_B[10][15] +
                  mat_A[10][11] * mat_B[11][15] +
                  mat_A[10][12] * mat_B[12][15] +
                  mat_A[10][13] * mat_B[13][15] +
                  mat_A[10][14] * mat_B[14][15] +
                  mat_A[10][15] * mat_B[15][15] +
                  mat_A[10][16] * mat_B[16][15] +
                  mat_A[10][17] * mat_B[17][15] +
                  mat_A[10][18] * mat_B[18][15] +
                  mat_A[10][19] * mat_B[19][15] +
                  mat_A[10][20] * mat_B[20][15] +
                  mat_A[10][21] * mat_B[21][15] +
                  mat_A[10][22] * mat_B[22][15] +
                  mat_A[10][23] * mat_B[23][15] +
                  mat_A[10][24] * mat_B[24][15] +
                  mat_A[10][25] * mat_B[25][15] +
                  mat_A[10][26] * mat_B[26][15] +
                  mat_A[10][27] * mat_B[27][15] +
                  mat_A[10][28] * mat_B[28][15] +
                  mat_A[10][29] * mat_B[29][15] +
                  mat_A[10][30] * mat_B[30][15] +
                  mat_A[10][31] * mat_B[31][15];
    mat_C[10][16] <= 
                  mat_A[10][0] * mat_B[0][16] +
                  mat_A[10][1] * mat_B[1][16] +
                  mat_A[10][2] * mat_B[2][16] +
                  mat_A[10][3] * mat_B[3][16] +
                  mat_A[10][4] * mat_B[4][16] +
                  mat_A[10][5] * mat_B[5][16] +
                  mat_A[10][6] * mat_B[6][16] +
                  mat_A[10][7] * mat_B[7][16] +
                  mat_A[10][8] * mat_B[8][16] +
                  mat_A[10][9] * mat_B[9][16] +
                  mat_A[10][10] * mat_B[10][16] +
                  mat_A[10][11] * mat_B[11][16] +
                  mat_A[10][12] * mat_B[12][16] +
                  mat_A[10][13] * mat_B[13][16] +
                  mat_A[10][14] * mat_B[14][16] +
                  mat_A[10][15] * mat_B[15][16] +
                  mat_A[10][16] * mat_B[16][16] +
                  mat_A[10][17] * mat_B[17][16] +
                  mat_A[10][18] * mat_B[18][16] +
                  mat_A[10][19] * mat_B[19][16] +
                  mat_A[10][20] * mat_B[20][16] +
                  mat_A[10][21] * mat_B[21][16] +
                  mat_A[10][22] * mat_B[22][16] +
                  mat_A[10][23] * mat_B[23][16] +
                  mat_A[10][24] * mat_B[24][16] +
                  mat_A[10][25] * mat_B[25][16] +
                  mat_A[10][26] * mat_B[26][16] +
                  mat_A[10][27] * mat_B[27][16] +
                  mat_A[10][28] * mat_B[28][16] +
                  mat_A[10][29] * mat_B[29][16] +
                  mat_A[10][30] * mat_B[30][16] +
                  mat_A[10][31] * mat_B[31][16];
    mat_C[10][17] <= 
                  mat_A[10][0] * mat_B[0][17] +
                  mat_A[10][1] * mat_B[1][17] +
                  mat_A[10][2] * mat_B[2][17] +
                  mat_A[10][3] * mat_B[3][17] +
                  mat_A[10][4] * mat_B[4][17] +
                  mat_A[10][5] * mat_B[5][17] +
                  mat_A[10][6] * mat_B[6][17] +
                  mat_A[10][7] * mat_B[7][17] +
                  mat_A[10][8] * mat_B[8][17] +
                  mat_A[10][9] * mat_B[9][17] +
                  mat_A[10][10] * mat_B[10][17] +
                  mat_A[10][11] * mat_B[11][17] +
                  mat_A[10][12] * mat_B[12][17] +
                  mat_A[10][13] * mat_B[13][17] +
                  mat_A[10][14] * mat_B[14][17] +
                  mat_A[10][15] * mat_B[15][17] +
                  mat_A[10][16] * mat_B[16][17] +
                  mat_A[10][17] * mat_B[17][17] +
                  mat_A[10][18] * mat_B[18][17] +
                  mat_A[10][19] * mat_B[19][17] +
                  mat_A[10][20] * mat_B[20][17] +
                  mat_A[10][21] * mat_B[21][17] +
                  mat_A[10][22] * mat_B[22][17] +
                  mat_A[10][23] * mat_B[23][17] +
                  mat_A[10][24] * mat_B[24][17] +
                  mat_A[10][25] * mat_B[25][17] +
                  mat_A[10][26] * mat_B[26][17] +
                  mat_A[10][27] * mat_B[27][17] +
                  mat_A[10][28] * mat_B[28][17] +
                  mat_A[10][29] * mat_B[29][17] +
                  mat_A[10][30] * mat_B[30][17] +
                  mat_A[10][31] * mat_B[31][17];
    mat_C[10][18] <= 
                  mat_A[10][0] * mat_B[0][18] +
                  mat_A[10][1] * mat_B[1][18] +
                  mat_A[10][2] * mat_B[2][18] +
                  mat_A[10][3] * mat_B[3][18] +
                  mat_A[10][4] * mat_B[4][18] +
                  mat_A[10][5] * mat_B[5][18] +
                  mat_A[10][6] * mat_B[6][18] +
                  mat_A[10][7] * mat_B[7][18] +
                  mat_A[10][8] * mat_B[8][18] +
                  mat_A[10][9] * mat_B[9][18] +
                  mat_A[10][10] * mat_B[10][18] +
                  mat_A[10][11] * mat_B[11][18] +
                  mat_A[10][12] * mat_B[12][18] +
                  mat_A[10][13] * mat_B[13][18] +
                  mat_A[10][14] * mat_B[14][18] +
                  mat_A[10][15] * mat_B[15][18] +
                  mat_A[10][16] * mat_B[16][18] +
                  mat_A[10][17] * mat_B[17][18] +
                  mat_A[10][18] * mat_B[18][18] +
                  mat_A[10][19] * mat_B[19][18] +
                  mat_A[10][20] * mat_B[20][18] +
                  mat_A[10][21] * mat_B[21][18] +
                  mat_A[10][22] * mat_B[22][18] +
                  mat_A[10][23] * mat_B[23][18] +
                  mat_A[10][24] * mat_B[24][18] +
                  mat_A[10][25] * mat_B[25][18] +
                  mat_A[10][26] * mat_B[26][18] +
                  mat_A[10][27] * mat_B[27][18] +
                  mat_A[10][28] * mat_B[28][18] +
                  mat_A[10][29] * mat_B[29][18] +
                  mat_A[10][30] * mat_B[30][18] +
                  mat_A[10][31] * mat_B[31][18];
    mat_C[10][19] <= 
                  mat_A[10][0] * mat_B[0][19] +
                  mat_A[10][1] * mat_B[1][19] +
                  mat_A[10][2] * mat_B[2][19] +
                  mat_A[10][3] * mat_B[3][19] +
                  mat_A[10][4] * mat_B[4][19] +
                  mat_A[10][5] * mat_B[5][19] +
                  mat_A[10][6] * mat_B[6][19] +
                  mat_A[10][7] * mat_B[7][19] +
                  mat_A[10][8] * mat_B[8][19] +
                  mat_A[10][9] * mat_B[9][19] +
                  mat_A[10][10] * mat_B[10][19] +
                  mat_A[10][11] * mat_B[11][19] +
                  mat_A[10][12] * mat_B[12][19] +
                  mat_A[10][13] * mat_B[13][19] +
                  mat_A[10][14] * mat_B[14][19] +
                  mat_A[10][15] * mat_B[15][19] +
                  mat_A[10][16] * mat_B[16][19] +
                  mat_A[10][17] * mat_B[17][19] +
                  mat_A[10][18] * mat_B[18][19] +
                  mat_A[10][19] * mat_B[19][19] +
                  mat_A[10][20] * mat_B[20][19] +
                  mat_A[10][21] * mat_B[21][19] +
                  mat_A[10][22] * mat_B[22][19] +
                  mat_A[10][23] * mat_B[23][19] +
                  mat_A[10][24] * mat_B[24][19] +
                  mat_A[10][25] * mat_B[25][19] +
                  mat_A[10][26] * mat_B[26][19] +
                  mat_A[10][27] * mat_B[27][19] +
                  mat_A[10][28] * mat_B[28][19] +
                  mat_A[10][29] * mat_B[29][19] +
                  mat_A[10][30] * mat_B[30][19] +
                  mat_A[10][31] * mat_B[31][19];
    mat_C[10][20] <= 
                  mat_A[10][0] * mat_B[0][20] +
                  mat_A[10][1] * mat_B[1][20] +
                  mat_A[10][2] * mat_B[2][20] +
                  mat_A[10][3] * mat_B[3][20] +
                  mat_A[10][4] * mat_B[4][20] +
                  mat_A[10][5] * mat_B[5][20] +
                  mat_A[10][6] * mat_B[6][20] +
                  mat_A[10][7] * mat_B[7][20] +
                  mat_A[10][8] * mat_B[8][20] +
                  mat_A[10][9] * mat_B[9][20] +
                  mat_A[10][10] * mat_B[10][20] +
                  mat_A[10][11] * mat_B[11][20] +
                  mat_A[10][12] * mat_B[12][20] +
                  mat_A[10][13] * mat_B[13][20] +
                  mat_A[10][14] * mat_B[14][20] +
                  mat_A[10][15] * mat_B[15][20] +
                  mat_A[10][16] * mat_B[16][20] +
                  mat_A[10][17] * mat_B[17][20] +
                  mat_A[10][18] * mat_B[18][20] +
                  mat_A[10][19] * mat_B[19][20] +
                  mat_A[10][20] * mat_B[20][20] +
                  mat_A[10][21] * mat_B[21][20] +
                  mat_A[10][22] * mat_B[22][20] +
                  mat_A[10][23] * mat_B[23][20] +
                  mat_A[10][24] * mat_B[24][20] +
                  mat_A[10][25] * mat_B[25][20] +
                  mat_A[10][26] * mat_B[26][20] +
                  mat_A[10][27] * mat_B[27][20] +
                  mat_A[10][28] * mat_B[28][20] +
                  mat_A[10][29] * mat_B[29][20] +
                  mat_A[10][30] * mat_B[30][20] +
                  mat_A[10][31] * mat_B[31][20];
    mat_C[10][21] <= 
                  mat_A[10][0] * mat_B[0][21] +
                  mat_A[10][1] * mat_B[1][21] +
                  mat_A[10][2] * mat_B[2][21] +
                  mat_A[10][3] * mat_B[3][21] +
                  mat_A[10][4] * mat_B[4][21] +
                  mat_A[10][5] * mat_B[5][21] +
                  mat_A[10][6] * mat_B[6][21] +
                  mat_A[10][7] * mat_B[7][21] +
                  mat_A[10][8] * mat_B[8][21] +
                  mat_A[10][9] * mat_B[9][21] +
                  mat_A[10][10] * mat_B[10][21] +
                  mat_A[10][11] * mat_B[11][21] +
                  mat_A[10][12] * mat_B[12][21] +
                  mat_A[10][13] * mat_B[13][21] +
                  mat_A[10][14] * mat_B[14][21] +
                  mat_A[10][15] * mat_B[15][21] +
                  mat_A[10][16] * mat_B[16][21] +
                  mat_A[10][17] * mat_B[17][21] +
                  mat_A[10][18] * mat_B[18][21] +
                  mat_A[10][19] * mat_B[19][21] +
                  mat_A[10][20] * mat_B[20][21] +
                  mat_A[10][21] * mat_B[21][21] +
                  mat_A[10][22] * mat_B[22][21] +
                  mat_A[10][23] * mat_B[23][21] +
                  mat_A[10][24] * mat_B[24][21] +
                  mat_A[10][25] * mat_B[25][21] +
                  mat_A[10][26] * mat_B[26][21] +
                  mat_A[10][27] * mat_B[27][21] +
                  mat_A[10][28] * mat_B[28][21] +
                  mat_A[10][29] * mat_B[29][21] +
                  mat_A[10][30] * mat_B[30][21] +
                  mat_A[10][31] * mat_B[31][21];
    mat_C[10][22] <= 
                  mat_A[10][0] * mat_B[0][22] +
                  mat_A[10][1] * mat_B[1][22] +
                  mat_A[10][2] * mat_B[2][22] +
                  mat_A[10][3] * mat_B[3][22] +
                  mat_A[10][4] * mat_B[4][22] +
                  mat_A[10][5] * mat_B[5][22] +
                  mat_A[10][6] * mat_B[6][22] +
                  mat_A[10][7] * mat_B[7][22] +
                  mat_A[10][8] * mat_B[8][22] +
                  mat_A[10][9] * mat_B[9][22] +
                  mat_A[10][10] * mat_B[10][22] +
                  mat_A[10][11] * mat_B[11][22] +
                  mat_A[10][12] * mat_B[12][22] +
                  mat_A[10][13] * mat_B[13][22] +
                  mat_A[10][14] * mat_B[14][22] +
                  mat_A[10][15] * mat_B[15][22] +
                  mat_A[10][16] * mat_B[16][22] +
                  mat_A[10][17] * mat_B[17][22] +
                  mat_A[10][18] * mat_B[18][22] +
                  mat_A[10][19] * mat_B[19][22] +
                  mat_A[10][20] * mat_B[20][22] +
                  mat_A[10][21] * mat_B[21][22] +
                  mat_A[10][22] * mat_B[22][22] +
                  mat_A[10][23] * mat_B[23][22] +
                  mat_A[10][24] * mat_B[24][22] +
                  mat_A[10][25] * mat_B[25][22] +
                  mat_A[10][26] * mat_B[26][22] +
                  mat_A[10][27] * mat_B[27][22] +
                  mat_A[10][28] * mat_B[28][22] +
                  mat_A[10][29] * mat_B[29][22] +
                  mat_A[10][30] * mat_B[30][22] +
                  mat_A[10][31] * mat_B[31][22];
    mat_C[10][23] <= 
                  mat_A[10][0] * mat_B[0][23] +
                  mat_A[10][1] * mat_B[1][23] +
                  mat_A[10][2] * mat_B[2][23] +
                  mat_A[10][3] * mat_B[3][23] +
                  mat_A[10][4] * mat_B[4][23] +
                  mat_A[10][5] * mat_B[5][23] +
                  mat_A[10][6] * mat_B[6][23] +
                  mat_A[10][7] * mat_B[7][23] +
                  mat_A[10][8] * mat_B[8][23] +
                  mat_A[10][9] * mat_B[9][23] +
                  mat_A[10][10] * mat_B[10][23] +
                  mat_A[10][11] * mat_B[11][23] +
                  mat_A[10][12] * mat_B[12][23] +
                  mat_A[10][13] * mat_B[13][23] +
                  mat_A[10][14] * mat_B[14][23] +
                  mat_A[10][15] * mat_B[15][23] +
                  mat_A[10][16] * mat_B[16][23] +
                  mat_A[10][17] * mat_B[17][23] +
                  mat_A[10][18] * mat_B[18][23] +
                  mat_A[10][19] * mat_B[19][23] +
                  mat_A[10][20] * mat_B[20][23] +
                  mat_A[10][21] * mat_B[21][23] +
                  mat_A[10][22] * mat_B[22][23] +
                  mat_A[10][23] * mat_B[23][23] +
                  mat_A[10][24] * mat_B[24][23] +
                  mat_A[10][25] * mat_B[25][23] +
                  mat_A[10][26] * mat_B[26][23] +
                  mat_A[10][27] * mat_B[27][23] +
                  mat_A[10][28] * mat_B[28][23] +
                  mat_A[10][29] * mat_B[29][23] +
                  mat_A[10][30] * mat_B[30][23] +
                  mat_A[10][31] * mat_B[31][23];
    mat_C[10][24] <= 
                  mat_A[10][0] * mat_B[0][24] +
                  mat_A[10][1] * mat_B[1][24] +
                  mat_A[10][2] * mat_B[2][24] +
                  mat_A[10][3] * mat_B[3][24] +
                  mat_A[10][4] * mat_B[4][24] +
                  mat_A[10][5] * mat_B[5][24] +
                  mat_A[10][6] * mat_B[6][24] +
                  mat_A[10][7] * mat_B[7][24] +
                  mat_A[10][8] * mat_B[8][24] +
                  mat_A[10][9] * mat_B[9][24] +
                  mat_A[10][10] * mat_B[10][24] +
                  mat_A[10][11] * mat_B[11][24] +
                  mat_A[10][12] * mat_B[12][24] +
                  mat_A[10][13] * mat_B[13][24] +
                  mat_A[10][14] * mat_B[14][24] +
                  mat_A[10][15] * mat_B[15][24] +
                  mat_A[10][16] * mat_B[16][24] +
                  mat_A[10][17] * mat_B[17][24] +
                  mat_A[10][18] * mat_B[18][24] +
                  mat_A[10][19] * mat_B[19][24] +
                  mat_A[10][20] * mat_B[20][24] +
                  mat_A[10][21] * mat_B[21][24] +
                  mat_A[10][22] * mat_B[22][24] +
                  mat_A[10][23] * mat_B[23][24] +
                  mat_A[10][24] * mat_B[24][24] +
                  mat_A[10][25] * mat_B[25][24] +
                  mat_A[10][26] * mat_B[26][24] +
                  mat_A[10][27] * mat_B[27][24] +
                  mat_A[10][28] * mat_B[28][24] +
                  mat_A[10][29] * mat_B[29][24] +
                  mat_A[10][30] * mat_B[30][24] +
                  mat_A[10][31] * mat_B[31][24];
    mat_C[10][25] <= 
                  mat_A[10][0] * mat_B[0][25] +
                  mat_A[10][1] * mat_B[1][25] +
                  mat_A[10][2] * mat_B[2][25] +
                  mat_A[10][3] * mat_B[3][25] +
                  mat_A[10][4] * mat_B[4][25] +
                  mat_A[10][5] * mat_B[5][25] +
                  mat_A[10][6] * mat_B[6][25] +
                  mat_A[10][7] * mat_B[7][25] +
                  mat_A[10][8] * mat_B[8][25] +
                  mat_A[10][9] * mat_B[9][25] +
                  mat_A[10][10] * mat_B[10][25] +
                  mat_A[10][11] * mat_B[11][25] +
                  mat_A[10][12] * mat_B[12][25] +
                  mat_A[10][13] * mat_B[13][25] +
                  mat_A[10][14] * mat_B[14][25] +
                  mat_A[10][15] * mat_B[15][25] +
                  mat_A[10][16] * mat_B[16][25] +
                  mat_A[10][17] * mat_B[17][25] +
                  mat_A[10][18] * mat_B[18][25] +
                  mat_A[10][19] * mat_B[19][25] +
                  mat_A[10][20] * mat_B[20][25] +
                  mat_A[10][21] * mat_B[21][25] +
                  mat_A[10][22] * mat_B[22][25] +
                  mat_A[10][23] * mat_B[23][25] +
                  mat_A[10][24] * mat_B[24][25] +
                  mat_A[10][25] * mat_B[25][25] +
                  mat_A[10][26] * mat_B[26][25] +
                  mat_A[10][27] * mat_B[27][25] +
                  mat_A[10][28] * mat_B[28][25] +
                  mat_A[10][29] * mat_B[29][25] +
                  mat_A[10][30] * mat_B[30][25] +
                  mat_A[10][31] * mat_B[31][25];
    mat_C[10][26] <= 
                  mat_A[10][0] * mat_B[0][26] +
                  mat_A[10][1] * mat_B[1][26] +
                  mat_A[10][2] * mat_B[2][26] +
                  mat_A[10][3] * mat_B[3][26] +
                  mat_A[10][4] * mat_B[4][26] +
                  mat_A[10][5] * mat_B[5][26] +
                  mat_A[10][6] * mat_B[6][26] +
                  mat_A[10][7] * mat_B[7][26] +
                  mat_A[10][8] * mat_B[8][26] +
                  mat_A[10][9] * mat_B[9][26] +
                  mat_A[10][10] * mat_B[10][26] +
                  mat_A[10][11] * mat_B[11][26] +
                  mat_A[10][12] * mat_B[12][26] +
                  mat_A[10][13] * mat_B[13][26] +
                  mat_A[10][14] * mat_B[14][26] +
                  mat_A[10][15] * mat_B[15][26] +
                  mat_A[10][16] * mat_B[16][26] +
                  mat_A[10][17] * mat_B[17][26] +
                  mat_A[10][18] * mat_B[18][26] +
                  mat_A[10][19] * mat_B[19][26] +
                  mat_A[10][20] * mat_B[20][26] +
                  mat_A[10][21] * mat_B[21][26] +
                  mat_A[10][22] * mat_B[22][26] +
                  mat_A[10][23] * mat_B[23][26] +
                  mat_A[10][24] * mat_B[24][26] +
                  mat_A[10][25] * mat_B[25][26] +
                  mat_A[10][26] * mat_B[26][26] +
                  mat_A[10][27] * mat_B[27][26] +
                  mat_A[10][28] * mat_B[28][26] +
                  mat_A[10][29] * mat_B[29][26] +
                  mat_A[10][30] * mat_B[30][26] +
                  mat_A[10][31] * mat_B[31][26];
    mat_C[10][27] <= 
                  mat_A[10][0] * mat_B[0][27] +
                  mat_A[10][1] * mat_B[1][27] +
                  mat_A[10][2] * mat_B[2][27] +
                  mat_A[10][3] * mat_B[3][27] +
                  mat_A[10][4] * mat_B[4][27] +
                  mat_A[10][5] * mat_B[5][27] +
                  mat_A[10][6] * mat_B[6][27] +
                  mat_A[10][7] * mat_B[7][27] +
                  mat_A[10][8] * mat_B[8][27] +
                  mat_A[10][9] * mat_B[9][27] +
                  mat_A[10][10] * mat_B[10][27] +
                  mat_A[10][11] * mat_B[11][27] +
                  mat_A[10][12] * mat_B[12][27] +
                  mat_A[10][13] * mat_B[13][27] +
                  mat_A[10][14] * mat_B[14][27] +
                  mat_A[10][15] * mat_B[15][27] +
                  mat_A[10][16] * mat_B[16][27] +
                  mat_A[10][17] * mat_B[17][27] +
                  mat_A[10][18] * mat_B[18][27] +
                  mat_A[10][19] * mat_B[19][27] +
                  mat_A[10][20] * mat_B[20][27] +
                  mat_A[10][21] * mat_B[21][27] +
                  mat_A[10][22] * mat_B[22][27] +
                  mat_A[10][23] * mat_B[23][27] +
                  mat_A[10][24] * mat_B[24][27] +
                  mat_A[10][25] * mat_B[25][27] +
                  mat_A[10][26] * mat_B[26][27] +
                  mat_A[10][27] * mat_B[27][27] +
                  mat_A[10][28] * mat_B[28][27] +
                  mat_A[10][29] * mat_B[29][27] +
                  mat_A[10][30] * mat_B[30][27] +
                  mat_A[10][31] * mat_B[31][27];
    mat_C[10][28] <= 
                  mat_A[10][0] * mat_B[0][28] +
                  mat_A[10][1] * mat_B[1][28] +
                  mat_A[10][2] * mat_B[2][28] +
                  mat_A[10][3] * mat_B[3][28] +
                  mat_A[10][4] * mat_B[4][28] +
                  mat_A[10][5] * mat_B[5][28] +
                  mat_A[10][6] * mat_B[6][28] +
                  mat_A[10][7] * mat_B[7][28] +
                  mat_A[10][8] * mat_B[8][28] +
                  mat_A[10][9] * mat_B[9][28] +
                  mat_A[10][10] * mat_B[10][28] +
                  mat_A[10][11] * mat_B[11][28] +
                  mat_A[10][12] * mat_B[12][28] +
                  mat_A[10][13] * mat_B[13][28] +
                  mat_A[10][14] * mat_B[14][28] +
                  mat_A[10][15] * mat_B[15][28] +
                  mat_A[10][16] * mat_B[16][28] +
                  mat_A[10][17] * mat_B[17][28] +
                  mat_A[10][18] * mat_B[18][28] +
                  mat_A[10][19] * mat_B[19][28] +
                  mat_A[10][20] * mat_B[20][28] +
                  mat_A[10][21] * mat_B[21][28] +
                  mat_A[10][22] * mat_B[22][28] +
                  mat_A[10][23] * mat_B[23][28] +
                  mat_A[10][24] * mat_B[24][28] +
                  mat_A[10][25] * mat_B[25][28] +
                  mat_A[10][26] * mat_B[26][28] +
                  mat_A[10][27] * mat_B[27][28] +
                  mat_A[10][28] * mat_B[28][28] +
                  mat_A[10][29] * mat_B[29][28] +
                  mat_A[10][30] * mat_B[30][28] +
                  mat_A[10][31] * mat_B[31][28];
    mat_C[10][29] <= 
                  mat_A[10][0] * mat_B[0][29] +
                  mat_A[10][1] * mat_B[1][29] +
                  mat_A[10][2] * mat_B[2][29] +
                  mat_A[10][3] * mat_B[3][29] +
                  mat_A[10][4] * mat_B[4][29] +
                  mat_A[10][5] * mat_B[5][29] +
                  mat_A[10][6] * mat_B[6][29] +
                  mat_A[10][7] * mat_B[7][29] +
                  mat_A[10][8] * mat_B[8][29] +
                  mat_A[10][9] * mat_B[9][29] +
                  mat_A[10][10] * mat_B[10][29] +
                  mat_A[10][11] * mat_B[11][29] +
                  mat_A[10][12] * mat_B[12][29] +
                  mat_A[10][13] * mat_B[13][29] +
                  mat_A[10][14] * mat_B[14][29] +
                  mat_A[10][15] * mat_B[15][29] +
                  mat_A[10][16] * mat_B[16][29] +
                  mat_A[10][17] * mat_B[17][29] +
                  mat_A[10][18] * mat_B[18][29] +
                  mat_A[10][19] * mat_B[19][29] +
                  mat_A[10][20] * mat_B[20][29] +
                  mat_A[10][21] * mat_B[21][29] +
                  mat_A[10][22] * mat_B[22][29] +
                  mat_A[10][23] * mat_B[23][29] +
                  mat_A[10][24] * mat_B[24][29] +
                  mat_A[10][25] * mat_B[25][29] +
                  mat_A[10][26] * mat_B[26][29] +
                  mat_A[10][27] * mat_B[27][29] +
                  mat_A[10][28] * mat_B[28][29] +
                  mat_A[10][29] * mat_B[29][29] +
                  mat_A[10][30] * mat_B[30][29] +
                  mat_A[10][31] * mat_B[31][29];
    mat_C[10][30] <= 
                  mat_A[10][0] * mat_B[0][30] +
                  mat_A[10][1] * mat_B[1][30] +
                  mat_A[10][2] * mat_B[2][30] +
                  mat_A[10][3] * mat_B[3][30] +
                  mat_A[10][4] * mat_B[4][30] +
                  mat_A[10][5] * mat_B[5][30] +
                  mat_A[10][6] * mat_B[6][30] +
                  mat_A[10][7] * mat_B[7][30] +
                  mat_A[10][8] * mat_B[8][30] +
                  mat_A[10][9] * mat_B[9][30] +
                  mat_A[10][10] * mat_B[10][30] +
                  mat_A[10][11] * mat_B[11][30] +
                  mat_A[10][12] * mat_B[12][30] +
                  mat_A[10][13] * mat_B[13][30] +
                  mat_A[10][14] * mat_B[14][30] +
                  mat_A[10][15] * mat_B[15][30] +
                  mat_A[10][16] * mat_B[16][30] +
                  mat_A[10][17] * mat_B[17][30] +
                  mat_A[10][18] * mat_B[18][30] +
                  mat_A[10][19] * mat_B[19][30] +
                  mat_A[10][20] * mat_B[20][30] +
                  mat_A[10][21] * mat_B[21][30] +
                  mat_A[10][22] * mat_B[22][30] +
                  mat_A[10][23] * mat_B[23][30] +
                  mat_A[10][24] * mat_B[24][30] +
                  mat_A[10][25] * mat_B[25][30] +
                  mat_A[10][26] * mat_B[26][30] +
                  mat_A[10][27] * mat_B[27][30] +
                  mat_A[10][28] * mat_B[28][30] +
                  mat_A[10][29] * mat_B[29][30] +
                  mat_A[10][30] * mat_B[30][30] +
                  mat_A[10][31] * mat_B[31][30];
    mat_C[10][31] <= 
                  mat_A[10][0] * mat_B[0][31] +
                  mat_A[10][1] * mat_B[1][31] +
                  mat_A[10][2] * mat_B[2][31] +
                  mat_A[10][3] * mat_B[3][31] +
                  mat_A[10][4] * mat_B[4][31] +
                  mat_A[10][5] * mat_B[5][31] +
                  mat_A[10][6] * mat_B[6][31] +
                  mat_A[10][7] * mat_B[7][31] +
                  mat_A[10][8] * mat_B[8][31] +
                  mat_A[10][9] * mat_B[9][31] +
                  mat_A[10][10] * mat_B[10][31] +
                  mat_A[10][11] * mat_B[11][31] +
                  mat_A[10][12] * mat_B[12][31] +
                  mat_A[10][13] * mat_B[13][31] +
                  mat_A[10][14] * mat_B[14][31] +
                  mat_A[10][15] * mat_B[15][31] +
                  mat_A[10][16] * mat_B[16][31] +
                  mat_A[10][17] * mat_B[17][31] +
                  mat_A[10][18] * mat_B[18][31] +
                  mat_A[10][19] * mat_B[19][31] +
                  mat_A[10][20] * mat_B[20][31] +
                  mat_A[10][21] * mat_B[21][31] +
                  mat_A[10][22] * mat_B[22][31] +
                  mat_A[10][23] * mat_B[23][31] +
                  mat_A[10][24] * mat_B[24][31] +
                  mat_A[10][25] * mat_B[25][31] +
                  mat_A[10][26] * mat_B[26][31] +
                  mat_A[10][27] * mat_B[27][31] +
                  mat_A[10][28] * mat_B[28][31] +
                  mat_A[10][29] * mat_B[29][31] +
                  mat_A[10][30] * mat_B[30][31] +
                  mat_A[10][31] * mat_B[31][31];
    mat_C[11][0] <= 
                  mat_A[11][0] * mat_B[0][0] +
                  mat_A[11][1] * mat_B[1][0] +
                  mat_A[11][2] * mat_B[2][0] +
                  mat_A[11][3] * mat_B[3][0] +
                  mat_A[11][4] * mat_B[4][0] +
                  mat_A[11][5] * mat_B[5][0] +
                  mat_A[11][6] * mat_B[6][0] +
                  mat_A[11][7] * mat_B[7][0] +
                  mat_A[11][8] * mat_B[8][0] +
                  mat_A[11][9] * mat_B[9][0] +
                  mat_A[11][10] * mat_B[10][0] +
                  mat_A[11][11] * mat_B[11][0] +
                  mat_A[11][12] * mat_B[12][0] +
                  mat_A[11][13] * mat_B[13][0] +
                  mat_A[11][14] * mat_B[14][0] +
                  mat_A[11][15] * mat_B[15][0] +
                  mat_A[11][16] * mat_B[16][0] +
                  mat_A[11][17] * mat_B[17][0] +
                  mat_A[11][18] * mat_B[18][0] +
                  mat_A[11][19] * mat_B[19][0] +
                  mat_A[11][20] * mat_B[20][0] +
                  mat_A[11][21] * mat_B[21][0] +
                  mat_A[11][22] * mat_B[22][0] +
                  mat_A[11][23] * mat_B[23][0] +
                  mat_A[11][24] * mat_B[24][0] +
                  mat_A[11][25] * mat_B[25][0] +
                  mat_A[11][26] * mat_B[26][0] +
                  mat_A[11][27] * mat_B[27][0] +
                  mat_A[11][28] * mat_B[28][0] +
                  mat_A[11][29] * mat_B[29][0] +
                  mat_A[11][30] * mat_B[30][0] +
                  mat_A[11][31] * mat_B[31][0];
    mat_C[11][1] <= 
                  mat_A[11][0] * mat_B[0][1] +
                  mat_A[11][1] * mat_B[1][1] +
                  mat_A[11][2] * mat_B[2][1] +
                  mat_A[11][3] * mat_B[3][1] +
                  mat_A[11][4] * mat_B[4][1] +
                  mat_A[11][5] * mat_B[5][1] +
                  mat_A[11][6] * mat_B[6][1] +
                  mat_A[11][7] * mat_B[7][1] +
                  mat_A[11][8] * mat_B[8][1] +
                  mat_A[11][9] * mat_B[9][1] +
                  mat_A[11][10] * mat_B[10][1] +
                  mat_A[11][11] * mat_B[11][1] +
                  mat_A[11][12] * mat_B[12][1] +
                  mat_A[11][13] * mat_B[13][1] +
                  mat_A[11][14] * mat_B[14][1] +
                  mat_A[11][15] * mat_B[15][1] +
                  mat_A[11][16] * mat_B[16][1] +
                  mat_A[11][17] * mat_B[17][1] +
                  mat_A[11][18] * mat_B[18][1] +
                  mat_A[11][19] * mat_B[19][1] +
                  mat_A[11][20] * mat_B[20][1] +
                  mat_A[11][21] * mat_B[21][1] +
                  mat_A[11][22] * mat_B[22][1] +
                  mat_A[11][23] * mat_B[23][1] +
                  mat_A[11][24] * mat_B[24][1] +
                  mat_A[11][25] * mat_B[25][1] +
                  mat_A[11][26] * mat_B[26][1] +
                  mat_A[11][27] * mat_B[27][1] +
                  mat_A[11][28] * mat_B[28][1] +
                  mat_A[11][29] * mat_B[29][1] +
                  mat_A[11][30] * mat_B[30][1] +
                  mat_A[11][31] * mat_B[31][1];
    mat_C[11][2] <= 
                  mat_A[11][0] * mat_B[0][2] +
                  mat_A[11][1] * mat_B[1][2] +
                  mat_A[11][2] * mat_B[2][2] +
                  mat_A[11][3] * mat_B[3][2] +
                  mat_A[11][4] * mat_B[4][2] +
                  mat_A[11][5] * mat_B[5][2] +
                  mat_A[11][6] * mat_B[6][2] +
                  mat_A[11][7] * mat_B[7][2] +
                  mat_A[11][8] * mat_B[8][2] +
                  mat_A[11][9] * mat_B[9][2] +
                  mat_A[11][10] * mat_B[10][2] +
                  mat_A[11][11] * mat_B[11][2] +
                  mat_A[11][12] * mat_B[12][2] +
                  mat_A[11][13] * mat_B[13][2] +
                  mat_A[11][14] * mat_B[14][2] +
                  mat_A[11][15] * mat_B[15][2] +
                  mat_A[11][16] * mat_B[16][2] +
                  mat_A[11][17] * mat_B[17][2] +
                  mat_A[11][18] * mat_B[18][2] +
                  mat_A[11][19] * mat_B[19][2] +
                  mat_A[11][20] * mat_B[20][2] +
                  mat_A[11][21] * mat_B[21][2] +
                  mat_A[11][22] * mat_B[22][2] +
                  mat_A[11][23] * mat_B[23][2] +
                  mat_A[11][24] * mat_B[24][2] +
                  mat_A[11][25] * mat_B[25][2] +
                  mat_A[11][26] * mat_B[26][2] +
                  mat_A[11][27] * mat_B[27][2] +
                  mat_A[11][28] * mat_B[28][2] +
                  mat_A[11][29] * mat_B[29][2] +
                  mat_A[11][30] * mat_B[30][2] +
                  mat_A[11][31] * mat_B[31][2];
    mat_C[11][3] <= 
                  mat_A[11][0] * mat_B[0][3] +
                  mat_A[11][1] * mat_B[1][3] +
                  mat_A[11][2] * mat_B[2][3] +
                  mat_A[11][3] * mat_B[3][3] +
                  mat_A[11][4] * mat_B[4][3] +
                  mat_A[11][5] * mat_B[5][3] +
                  mat_A[11][6] * mat_B[6][3] +
                  mat_A[11][7] * mat_B[7][3] +
                  mat_A[11][8] * mat_B[8][3] +
                  mat_A[11][9] * mat_B[9][3] +
                  mat_A[11][10] * mat_B[10][3] +
                  mat_A[11][11] * mat_B[11][3] +
                  mat_A[11][12] * mat_B[12][3] +
                  mat_A[11][13] * mat_B[13][3] +
                  mat_A[11][14] * mat_B[14][3] +
                  mat_A[11][15] * mat_B[15][3] +
                  mat_A[11][16] * mat_B[16][3] +
                  mat_A[11][17] * mat_B[17][3] +
                  mat_A[11][18] * mat_B[18][3] +
                  mat_A[11][19] * mat_B[19][3] +
                  mat_A[11][20] * mat_B[20][3] +
                  mat_A[11][21] * mat_B[21][3] +
                  mat_A[11][22] * mat_B[22][3] +
                  mat_A[11][23] * mat_B[23][3] +
                  mat_A[11][24] * mat_B[24][3] +
                  mat_A[11][25] * mat_B[25][3] +
                  mat_A[11][26] * mat_B[26][3] +
                  mat_A[11][27] * mat_B[27][3] +
                  mat_A[11][28] * mat_B[28][3] +
                  mat_A[11][29] * mat_B[29][3] +
                  mat_A[11][30] * mat_B[30][3] +
                  mat_A[11][31] * mat_B[31][3];
    mat_C[11][4] <= 
                  mat_A[11][0] * mat_B[0][4] +
                  mat_A[11][1] * mat_B[1][4] +
                  mat_A[11][2] * mat_B[2][4] +
                  mat_A[11][3] * mat_B[3][4] +
                  mat_A[11][4] * mat_B[4][4] +
                  mat_A[11][5] * mat_B[5][4] +
                  mat_A[11][6] * mat_B[6][4] +
                  mat_A[11][7] * mat_B[7][4] +
                  mat_A[11][8] * mat_B[8][4] +
                  mat_A[11][9] * mat_B[9][4] +
                  mat_A[11][10] * mat_B[10][4] +
                  mat_A[11][11] * mat_B[11][4] +
                  mat_A[11][12] * mat_B[12][4] +
                  mat_A[11][13] * mat_B[13][4] +
                  mat_A[11][14] * mat_B[14][4] +
                  mat_A[11][15] * mat_B[15][4] +
                  mat_A[11][16] * mat_B[16][4] +
                  mat_A[11][17] * mat_B[17][4] +
                  mat_A[11][18] * mat_B[18][4] +
                  mat_A[11][19] * mat_B[19][4] +
                  mat_A[11][20] * mat_B[20][4] +
                  mat_A[11][21] * mat_B[21][4] +
                  mat_A[11][22] * mat_B[22][4] +
                  mat_A[11][23] * mat_B[23][4] +
                  mat_A[11][24] * mat_B[24][4] +
                  mat_A[11][25] * mat_B[25][4] +
                  mat_A[11][26] * mat_B[26][4] +
                  mat_A[11][27] * mat_B[27][4] +
                  mat_A[11][28] * mat_B[28][4] +
                  mat_A[11][29] * mat_B[29][4] +
                  mat_A[11][30] * mat_B[30][4] +
                  mat_A[11][31] * mat_B[31][4];
    mat_C[11][5] <= 
                  mat_A[11][0] * mat_B[0][5] +
                  mat_A[11][1] * mat_B[1][5] +
                  mat_A[11][2] * mat_B[2][5] +
                  mat_A[11][3] * mat_B[3][5] +
                  mat_A[11][4] * mat_B[4][5] +
                  mat_A[11][5] * mat_B[5][5] +
                  mat_A[11][6] * mat_B[6][5] +
                  mat_A[11][7] * mat_B[7][5] +
                  mat_A[11][8] * mat_B[8][5] +
                  mat_A[11][9] * mat_B[9][5] +
                  mat_A[11][10] * mat_B[10][5] +
                  mat_A[11][11] * mat_B[11][5] +
                  mat_A[11][12] * mat_B[12][5] +
                  mat_A[11][13] * mat_B[13][5] +
                  mat_A[11][14] * mat_B[14][5] +
                  mat_A[11][15] * mat_B[15][5] +
                  mat_A[11][16] * mat_B[16][5] +
                  mat_A[11][17] * mat_B[17][5] +
                  mat_A[11][18] * mat_B[18][5] +
                  mat_A[11][19] * mat_B[19][5] +
                  mat_A[11][20] * mat_B[20][5] +
                  mat_A[11][21] * mat_B[21][5] +
                  mat_A[11][22] * mat_B[22][5] +
                  mat_A[11][23] * mat_B[23][5] +
                  mat_A[11][24] * mat_B[24][5] +
                  mat_A[11][25] * mat_B[25][5] +
                  mat_A[11][26] * mat_B[26][5] +
                  mat_A[11][27] * mat_B[27][5] +
                  mat_A[11][28] * mat_B[28][5] +
                  mat_A[11][29] * mat_B[29][5] +
                  mat_A[11][30] * mat_B[30][5] +
                  mat_A[11][31] * mat_B[31][5];
    mat_C[11][6] <= 
                  mat_A[11][0] * mat_B[0][6] +
                  mat_A[11][1] * mat_B[1][6] +
                  mat_A[11][2] * mat_B[2][6] +
                  mat_A[11][3] * mat_B[3][6] +
                  mat_A[11][4] * mat_B[4][6] +
                  mat_A[11][5] * mat_B[5][6] +
                  mat_A[11][6] * mat_B[6][6] +
                  mat_A[11][7] * mat_B[7][6] +
                  mat_A[11][8] * mat_B[8][6] +
                  mat_A[11][9] * mat_B[9][6] +
                  mat_A[11][10] * mat_B[10][6] +
                  mat_A[11][11] * mat_B[11][6] +
                  mat_A[11][12] * mat_B[12][6] +
                  mat_A[11][13] * mat_B[13][6] +
                  mat_A[11][14] * mat_B[14][6] +
                  mat_A[11][15] * mat_B[15][6] +
                  mat_A[11][16] * mat_B[16][6] +
                  mat_A[11][17] * mat_B[17][6] +
                  mat_A[11][18] * mat_B[18][6] +
                  mat_A[11][19] * mat_B[19][6] +
                  mat_A[11][20] * mat_B[20][6] +
                  mat_A[11][21] * mat_B[21][6] +
                  mat_A[11][22] * mat_B[22][6] +
                  mat_A[11][23] * mat_B[23][6] +
                  mat_A[11][24] * mat_B[24][6] +
                  mat_A[11][25] * mat_B[25][6] +
                  mat_A[11][26] * mat_B[26][6] +
                  mat_A[11][27] * mat_B[27][6] +
                  mat_A[11][28] * mat_B[28][6] +
                  mat_A[11][29] * mat_B[29][6] +
                  mat_A[11][30] * mat_B[30][6] +
                  mat_A[11][31] * mat_B[31][6];
    mat_C[11][7] <= 
                  mat_A[11][0] * mat_B[0][7] +
                  mat_A[11][1] * mat_B[1][7] +
                  mat_A[11][2] * mat_B[2][7] +
                  mat_A[11][3] * mat_B[3][7] +
                  mat_A[11][4] * mat_B[4][7] +
                  mat_A[11][5] * mat_B[5][7] +
                  mat_A[11][6] * mat_B[6][7] +
                  mat_A[11][7] * mat_B[7][7] +
                  mat_A[11][8] * mat_B[8][7] +
                  mat_A[11][9] * mat_B[9][7] +
                  mat_A[11][10] * mat_B[10][7] +
                  mat_A[11][11] * mat_B[11][7] +
                  mat_A[11][12] * mat_B[12][7] +
                  mat_A[11][13] * mat_B[13][7] +
                  mat_A[11][14] * mat_B[14][7] +
                  mat_A[11][15] * mat_B[15][7] +
                  mat_A[11][16] * mat_B[16][7] +
                  mat_A[11][17] * mat_B[17][7] +
                  mat_A[11][18] * mat_B[18][7] +
                  mat_A[11][19] * mat_B[19][7] +
                  mat_A[11][20] * mat_B[20][7] +
                  mat_A[11][21] * mat_B[21][7] +
                  mat_A[11][22] * mat_B[22][7] +
                  mat_A[11][23] * mat_B[23][7] +
                  mat_A[11][24] * mat_B[24][7] +
                  mat_A[11][25] * mat_B[25][7] +
                  mat_A[11][26] * mat_B[26][7] +
                  mat_A[11][27] * mat_B[27][7] +
                  mat_A[11][28] * mat_B[28][7] +
                  mat_A[11][29] * mat_B[29][7] +
                  mat_A[11][30] * mat_B[30][7] +
                  mat_A[11][31] * mat_B[31][7];
    mat_C[11][8] <= 
                  mat_A[11][0] * mat_B[0][8] +
                  mat_A[11][1] * mat_B[1][8] +
                  mat_A[11][2] * mat_B[2][8] +
                  mat_A[11][3] * mat_B[3][8] +
                  mat_A[11][4] * mat_B[4][8] +
                  mat_A[11][5] * mat_B[5][8] +
                  mat_A[11][6] * mat_B[6][8] +
                  mat_A[11][7] * mat_B[7][8] +
                  mat_A[11][8] * mat_B[8][8] +
                  mat_A[11][9] * mat_B[9][8] +
                  mat_A[11][10] * mat_B[10][8] +
                  mat_A[11][11] * mat_B[11][8] +
                  mat_A[11][12] * mat_B[12][8] +
                  mat_A[11][13] * mat_B[13][8] +
                  mat_A[11][14] * mat_B[14][8] +
                  mat_A[11][15] * mat_B[15][8] +
                  mat_A[11][16] * mat_B[16][8] +
                  mat_A[11][17] * mat_B[17][8] +
                  mat_A[11][18] * mat_B[18][8] +
                  mat_A[11][19] * mat_B[19][8] +
                  mat_A[11][20] * mat_B[20][8] +
                  mat_A[11][21] * mat_B[21][8] +
                  mat_A[11][22] * mat_B[22][8] +
                  mat_A[11][23] * mat_B[23][8] +
                  mat_A[11][24] * mat_B[24][8] +
                  mat_A[11][25] * mat_B[25][8] +
                  mat_A[11][26] * mat_B[26][8] +
                  mat_A[11][27] * mat_B[27][8] +
                  mat_A[11][28] * mat_B[28][8] +
                  mat_A[11][29] * mat_B[29][8] +
                  mat_A[11][30] * mat_B[30][8] +
                  mat_A[11][31] * mat_B[31][8];
    mat_C[11][9] <= 
                  mat_A[11][0] * mat_B[0][9] +
                  mat_A[11][1] * mat_B[1][9] +
                  mat_A[11][2] * mat_B[2][9] +
                  mat_A[11][3] * mat_B[3][9] +
                  mat_A[11][4] * mat_B[4][9] +
                  mat_A[11][5] * mat_B[5][9] +
                  mat_A[11][6] * mat_B[6][9] +
                  mat_A[11][7] * mat_B[7][9] +
                  mat_A[11][8] * mat_B[8][9] +
                  mat_A[11][9] * mat_B[9][9] +
                  mat_A[11][10] * mat_B[10][9] +
                  mat_A[11][11] * mat_B[11][9] +
                  mat_A[11][12] * mat_B[12][9] +
                  mat_A[11][13] * mat_B[13][9] +
                  mat_A[11][14] * mat_B[14][9] +
                  mat_A[11][15] * mat_B[15][9] +
                  mat_A[11][16] * mat_B[16][9] +
                  mat_A[11][17] * mat_B[17][9] +
                  mat_A[11][18] * mat_B[18][9] +
                  mat_A[11][19] * mat_B[19][9] +
                  mat_A[11][20] * mat_B[20][9] +
                  mat_A[11][21] * mat_B[21][9] +
                  mat_A[11][22] * mat_B[22][9] +
                  mat_A[11][23] * mat_B[23][9] +
                  mat_A[11][24] * mat_B[24][9] +
                  mat_A[11][25] * mat_B[25][9] +
                  mat_A[11][26] * mat_B[26][9] +
                  mat_A[11][27] * mat_B[27][9] +
                  mat_A[11][28] * mat_B[28][9] +
                  mat_A[11][29] * mat_B[29][9] +
                  mat_A[11][30] * mat_B[30][9] +
                  mat_A[11][31] * mat_B[31][9];
    mat_C[11][10] <= 
                  mat_A[11][0] * mat_B[0][10] +
                  mat_A[11][1] * mat_B[1][10] +
                  mat_A[11][2] * mat_B[2][10] +
                  mat_A[11][3] * mat_B[3][10] +
                  mat_A[11][4] * mat_B[4][10] +
                  mat_A[11][5] * mat_B[5][10] +
                  mat_A[11][6] * mat_B[6][10] +
                  mat_A[11][7] * mat_B[7][10] +
                  mat_A[11][8] * mat_B[8][10] +
                  mat_A[11][9] * mat_B[9][10] +
                  mat_A[11][10] * mat_B[10][10] +
                  mat_A[11][11] * mat_B[11][10] +
                  mat_A[11][12] * mat_B[12][10] +
                  mat_A[11][13] * mat_B[13][10] +
                  mat_A[11][14] * mat_B[14][10] +
                  mat_A[11][15] * mat_B[15][10] +
                  mat_A[11][16] * mat_B[16][10] +
                  mat_A[11][17] * mat_B[17][10] +
                  mat_A[11][18] * mat_B[18][10] +
                  mat_A[11][19] * mat_B[19][10] +
                  mat_A[11][20] * mat_B[20][10] +
                  mat_A[11][21] * mat_B[21][10] +
                  mat_A[11][22] * mat_B[22][10] +
                  mat_A[11][23] * mat_B[23][10] +
                  mat_A[11][24] * mat_B[24][10] +
                  mat_A[11][25] * mat_B[25][10] +
                  mat_A[11][26] * mat_B[26][10] +
                  mat_A[11][27] * mat_B[27][10] +
                  mat_A[11][28] * mat_B[28][10] +
                  mat_A[11][29] * mat_B[29][10] +
                  mat_A[11][30] * mat_B[30][10] +
                  mat_A[11][31] * mat_B[31][10];
    mat_C[11][11] <= 
                  mat_A[11][0] * mat_B[0][11] +
                  mat_A[11][1] * mat_B[1][11] +
                  mat_A[11][2] * mat_B[2][11] +
                  mat_A[11][3] * mat_B[3][11] +
                  mat_A[11][4] * mat_B[4][11] +
                  mat_A[11][5] * mat_B[5][11] +
                  mat_A[11][6] * mat_B[6][11] +
                  mat_A[11][7] * mat_B[7][11] +
                  mat_A[11][8] * mat_B[8][11] +
                  mat_A[11][9] * mat_B[9][11] +
                  mat_A[11][10] * mat_B[10][11] +
                  mat_A[11][11] * mat_B[11][11] +
                  mat_A[11][12] * mat_B[12][11] +
                  mat_A[11][13] * mat_B[13][11] +
                  mat_A[11][14] * mat_B[14][11] +
                  mat_A[11][15] * mat_B[15][11] +
                  mat_A[11][16] * mat_B[16][11] +
                  mat_A[11][17] * mat_B[17][11] +
                  mat_A[11][18] * mat_B[18][11] +
                  mat_A[11][19] * mat_B[19][11] +
                  mat_A[11][20] * mat_B[20][11] +
                  mat_A[11][21] * mat_B[21][11] +
                  mat_A[11][22] * mat_B[22][11] +
                  mat_A[11][23] * mat_B[23][11] +
                  mat_A[11][24] * mat_B[24][11] +
                  mat_A[11][25] * mat_B[25][11] +
                  mat_A[11][26] * mat_B[26][11] +
                  mat_A[11][27] * mat_B[27][11] +
                  mat_A[11][28] * mat_B[28][11] +
                  mat_A[11][29] * mat_B[29][11] +
                  mat_A[11][30] * mat_B[30][11] +
                  mat_A[11][31] * mat_B[31][11];
    mat_C[11][12] <= 
                  mat_A[11][0] * mat_B[0][12] +
                  mat_A[11][1] * mat_B[1][12] +
                  mat_A[11][2] * mat_B[2][12] +
                  mat_A[11][3] * mat_B[3][12] +
                  mat_A[11][4] * mat_B[4][12] +
                  mat_A[11][5] * mat_B[5][12] +
                  mat_A[11][6] * mat_B[6][12] +
                  mat_A[11][7] * mat_B[7][12] +
                  mat_A[11][8] * mat_B[8][12] +
                  mat_A[11][9] * mat_B[9][12] +
                  mat_A[11][10] * mat_B[10][12] +
                  mat_A[11][11] * mat_B[11][12] +
                  mat_A[11][12] * mat_B[12][12] +
                  mat_A[11][13] * mat_B[13][12] +
                  mat_A[11][14] * mat_B[14][12] +
                  mat_A[11][15] * mat_B[15][12] +
                  mat_A[11][16] * mat_B[16][12] +
                  mat_A[11][17] * mat_B[17][12] +
                  mat_A[11][18] * mat_B[18][12] +
                  mat_A[11][19] * mat_B[19][12] +
                  mat_A[11][20] * mat_B[20][12] +
                  mat_A[11][21] * mat_B[21][12] +
                  mat_A[11][22] * mat_B[22][12] +
                  mat_A[11][23] * mat_B[23][12] +
                  mat_A[11][24] * mat_B[24][12] +
                  mat_A[11][25] * mat_B[25][12] +
                  mat_A[11][26] * mat_B[26][12] +
                  mat_A[11][27] * mat_B[27][12] +
                  mat_A[11][28] * mat_B[28][12] +
                  mat_A[11][29] * mat_B[29][12] +
                  mat_A[11][30] * mat_B[30][12] +
                  mat_A[11][31] * mat_B[31][12];
    mat_C[11][13] <= 
                  mat_A[11][0] * mat_B[0][13] +
                  mat_A[11][1] * mat_B[1][13] +
                  mat_A[11][2] * mat_B[2][13] +
                  mat_A[11][3] * mat_B[3][13] +
                  mat_A[11][4] * mat_B[4][13] +
                  mat_A[11][5] * mat_B[5][13] +
                  mat_A[11][6] * mat_B[6][13] +
                  mat_A[11][7] * mat_B[7][13] +
                  mat_A[11][8] * mat_B[8][13] +
                  mat_A[11][9] * mat_B[9][13] +
                  mat_A[11][10] * mat_B[10][13] +
                  mat_A[11][11] * mat_B[11][13] +
                  mat_A[11][12] * mat_B[12][13] +
                  mat_A[11][13] * mat_B[13][13] +
                  mat_A[11][14] * mat_B[14][13] +
                  mat_A[11][15] * mat_B[15][13] +
                  mat_A[11][16] * mat_B[16][13] +
                  mat_A[11][17] * mat_B[17][13] +
                  mat_A[11][18] * mat_B[18][13] +
                  mat_A[11][19] * mat_B[19][13] +
                  mat_A[11][20] * mat_B[20][13] +
                  mat_A[11][21] * mat_B[21][13] +
                  mat_A[11][22] * mat_B[22][13] +
                  mat_A[11][23] * mat_B[23][13] +
                  mat_A[11][24] * mat_B[24][13] +
                  mat_A[11][25] * mat_B[25][13] +
                  mat_A[11][26] * mat_B[26][13] +
                  mat_A[11][27] * mat_B[27][13] +
                  mat_A[11][28] * mat_B[28][13] +
                  mat_A[11][29] * mat_B[29][13] +
                  mat_A[11][30] * mat_B[30][13] +
                  mat_A[11][31] * mat_B[31][13];
    mat_C[11][14] <= 
                  mat_A[11][0] * mat_B[0][14] +
                  mat_A[11][1] * mat_B[1][14] +
                  mat_A[11][2] * mat_B[2][14] +
                  mat_A[11][3] * mat_B[3][14] +
                  mat_A[11][4] * mat_B[4][14] +
                  mat_A[11][5] * mat_B[5][14] +
                  mat_A[11][6] * mat_B[6][14] +
                  mat_A[11][7] * mat_B[7][14] +
                  mat_A[11][8] * mat_B[8][14] +
                  mat_A[11][9] * mat_B[9][14] +
                  mat_A[11][10] * mat_B[10][14] +
                  mat_A[11][11] * mat_B[11][14] +
                  mat_A[11][12] * mat_B[12][14] +
                  mat_A[11][13] * mat_B[13][14] +
                  mat_A[11][14] * mat_B[14][14] +
                  mat_A[11][15] * mat_B[15][14] +
                  mat_A[11][16] * mat_B[16][14] +
                  mat_A[11][17] * mat_B[17][14] +
                  mat_A[11][18] * mat_B[18][14] +
                  mat_A[11][19] * mat_B[19][14] +
                  mat_A[11][20] * mat_B[20][14] +
                  mat_A[11][21] * mat_B[21][14] +
                  mat_A[11][22] * mat_B[22][14] +
                  mat_A[11][23] * mat_B[23][14] +
                  mat_A[11][24] * mat_B[24][14] +
                  mat_A[11][25] * mat_B[25][14] +
                  mat_A[11][26] * mat_B[26][14] +
                  mat_A[11][27] * mat_B[27][14] +
                  mat_A[11][28] * mat_B[28][14] +
                  mat_A[11][29] * mat_B[29][14] +
                  mat_A[11][30] * mat_B[30][14] +
                  mat_A[11][31] * mat_B[31][14];
    mat_C[11][15] <= 
                  mat_A[11][0] * mat_B[0][15] +
                  mat_A[11][1] * mat_B[1][15] +
                  mat_A[11][2] * mat_B[2][15] +
                  mat_A[11][3] * mat_B[3][15] +
                  mat_A[11][4] * mat_B[4][15] +
                  mat_A[11][5] * mat_B[5][15] +
                  mat_A[11][6] * mat_B[6][15] +
                  mat_A[11][7] * mat_B[7][15] +
                  mat_A[11][8] * mat_B[8][15] +
                  mat_A[11][9] * mat_B[9][15] +
                  mat_A[11][10] * mat_B[10][15] +
                  mat_A[11][11] * mat_B[11][15] +
                  mat_A[11][12] * mat_B[12][15] +
                  mat_A[11][13] * mat_B[13][15] +
                  mat_A[11][14] * mat_B[14][15] +
                  mat_A[11][15] * mat_B[15][15] +
                  mat_A[11][16] * mat_B[16][15] +
                  mat_A[11][17] * mat_B[17][15] +
                  mat_A[11][18] * mat_B[18][15] +
                  mat_A[11][19] * mat_B[19][15] +
                  mat_A[11][20] * mat_B[20][15] +
                  mat_A[11][21] * mat_B[21][15] +
                  mat_A[11][22] * mat_B[22][15] +
                  mat_A[11][23] * mat_B[23][15] +
                  mat_A[11][24] * mat_B[24][15] +
                  mat_A[11][25] * mat_B[25][15] +
                  mat_A[11][26] * mat_B[26][15] +
                  mat_A[11][27] * mat_B[27][15] +
                  mat_A[11][28] * mat_B[28][15] +
                  mat_A[11][29] * mat_B[29][15] +
                  mat_A[11][30] * mat_B[30][15] +
                  mat_A[11][31] * mat_B[31][15];
    mat_C[11][16] <= 
                  mat_A[11][0] * mat_B[0][16] +
                  mat_A[11][1] * mat_B[1][16] +
                  mat_A[11][2] * mat_B[2][16] +
                  mat_A[11][3] * mat_B[3][16] +
                  mat_A[11][4] * mat_B[4][16] +
                  mat_A[11][5] * mat_B[5][16] +
                  mat_A[11][6] * mat_B[6][16] +
                  mat_A[11][7] * mat_B[7][16] +
                  mat_A[11][8] * mat_B[8][16] +
                  mat_A[11][9] * mat_B[9][16] +
                  mat_A[11][10] * mat_B[10][16] +
                  mat_A[11][11] * mat_B[11][16] +
                  mat_A[11][12] * mat_B[12][16] +
                  mat_A[11][13] * mat_B[13][16] +
                  mat_A[11][14] * mat_B[14][16] +
                  mat_A[11][15] * mat_B[15][16] +
                  mat_A[11][16] * mat_B[16][16] +
                  mat_A[11][17] * mat_B[17][16] +
                  mat_A[11][18] * mat_B[18][16] +
                  mat_A[11][19] * mat_B[19][16] +
                  mat_A[11][20] * mat_B[20][16] +
                  mat_A[11][21] * mat_B[21][16] +
                  mat_A[11][22] * mat_B[22][16] +
                  mat_A[11][23] * mat_B[23][16] +
                  mat_A[11][24] * mat_B[24][16] +
                  mat_A[11][25] * mat_B[25][16] +
                  mat_A[11][26] * mat_B[26][16] +
                  mat_A[11][27] * mat_B[27][16] +
                  mat_A[11][28] * mat_B[28][16] +
                  mat_A[11][29] * mat_B[29][16] +
                  mat_A[11][30] * mat_B[30][16] +
                  mat_A[11][31] * mat_B[31][16];
    mat_C[11][17] <= 
                  mat_A[11][0] * mat_B[0][17] +
                  mat_A[11][1] * mat_B[1][17] +
                  mat_A[11][2] * mat_B[2][17] +
                  mat_A[11][3] * mat_B[3][17] +
                  mat_A[11][4] * mat_B[4][17] +
                  mat_A[11][5] * mat_B[5][17] +
                  mat_A[11][6] * mat_B[6][17] +
                  mat_A[11][7] * mat_B[7][17] +
                  mat_A[11][8] * mat_B[8][17] +
                  mat_A[11][9] * mat_B[9][17] +
                  mat_A[11][10] * mat_B[10][17] +
                  mat_A[11][11] * mat_B[11][17] +
                  mat_A[11][12] * mat_B[12][17] +
                  mat_A[11][13] * mat_B[13][17] +
                  mat_A[11][14] * mat_B[14][17] +
                  mat_A[11][15] * mat_B[15][17] +
                  mat_A[11][16] * mat_B[16][17] +
                  mat_A[11][17] * mat_B[17][17] +
                  mat_A[11][18] * mat_B[18][17] +
                  mat_A[11][19] * mat_B[19][17] +
                  mat_A[11][20] * mat_B[20][17] +
                  mat_A[11][21] * mat_B[21][17] +
                  mat_A[11][22] * mat_B[22][17] +
                  mat_A[11][23] * mat_B[23][17] +
                  mat_A[11][24] * mat_B[24][17] +
                  mat_A[11][25] * mat_B[25][17] +
                  mat_A[11][26] * mat_B[26][17] +
                  mat_A[11][27] * mat_B[27][17] +
                  mat_A[11][28] * mat_B[28][17] +
                  mat_A[11][29] * mat_B[29][17] +
                  mat_A[11][30] * mat_B[30][17] +
                  mat_A[11][31] * mat_B[31][17];
    mat_C[11][18] <= 
                  mat_A[11][0] * mat_B[0][18] +
                  mat_A[11][1] * mat_B[1][18] +
                  mat_A[11][2] * mat_B[2][18] +
                  mat_A[11][3] * mat_B[3][18] +
                  mat_A[11][4] * mat_B[4][18] +
                  mat_A[11][5] * mat_B[5][18] +
                  mat_A[11][6] * mat_B[6][18] +
                  mat_A[11][7] * mat_B[7][18] +
                  mat_A[11][8] * mat_B[8][18] +
                  mat_A[11][9] * mat_B[9][18] +
                  mat_A[11][10] * mat_B[10][18] +
                  mat_A[11][11] * mat_B[11][18] +
                  mat_A[11][12] * mat_B[12][18] +
                  mat_A[11][13] * mat_B[13][18] +
                  mat_A[11][14] * mat_B[14][18] +
                  mat_A[11][15] * mat_B[15][18] +
                  mat_A[11][16] * mat_B[16][18] +
                  mat_A[11][17] * mat_B[17][18] +
                  mat_A[11][18] * mat_B[18][18] +
                  mat_A[11][19] * mat_B[19][18] +
                  mat_A[11][20] * mat_B[20][18] +
                  mat_A[11][21] * mat_B[21][18] +
                  mat_A[11][22] * mat_B[22][18] +
                  mat_A[11][23] * mat_B[23][18] +
                  mat_A[11][24] * mat_B[24][18] +
                  mat_A[11][25] * mat_B[25][18] +
                  mat_A[11][26] * mat_B[26][18] +
                  mat_A[11][27] * mat_B[27][18] +
                  mat_A[11][28] * mat_B[28][18] +
                  mat_A[11][29] * mat_B[29][18] +
                  mat_A[11][30] * mat_B[30][18] +
                  mat_A[11][31] * mat_B[31][18];
    mat_C[11][19] <= 
                  mat_A[11][0] * mat_B[0][19] +
                  mat_A[11][1] * mat_B[1][19] +
                  mat_A[11][2] * mat_B[2][19] +
                  mat_A[11][3] * mat_B[3][19] +
                  mat_A[11][4] * mat_B[4][19] +
                  mat_A[11][5] * mat_B[5][19] +
                  mat_A[11][6] * mat_B[6][19] +
                  mat_A[11][7] * mat_B[7][19] +
                  mat_A[11][8] * mat_B[8][19] +
                  mat_A[11][9] * mat_B[9][19] +
                  mat_A[11][10] * mat_B[10][19] +
                  mat_A[11][11] * mat_B[11][19] +
                  mat_A[11][12] * mat_B[12][19] +
                  mat_A[11][13] * mat_B[13][19] +
                  mat_A[11][14] * mat_B[14][19] +
                  mat_A[11][15] * mat_B[15][19] +
                  mat_A[11][16] * mat_B[16][19] +
                  mat_A[11][17] * mat_B[17][19] +
                  mat_A[11][18] * mat_B[18][19] +
                  mat_A[11][19] * mat_B[19][19] +
                  mat_A[11][20] * mat_B[20][19] +
                  mat_A[11][21] * mat_B[21][19] +
                  mat_A[11][22] * mat_B[22][19] +
                  mat_A[11][23] * mat_B[23][19] +
                  mat_A[11][24] * mat_B[24][19] +
                  mat_A[11][25] * mat_B[25][19] +
                  mat_A[11][26] * mat_B[26][19] +
                  mat_A[11][27] * mat_B[27][19] +
                  mat_A[11][28] * mat_B[28][19] +
                  mat_A[11][29] * mat_B[29][19] +
                  mat_A[11][30] * mat_B[30][19] +
                  mat_A[11][31] * mat_B[31][19];
    mat_C[11][20] <= 
                  mat_A[11][0] * mat_B[0][20] +
                  mat_A[11][1] * mat_B[1][20] +
                  mat_A[11][2] * mat_B[2][20] +
                  mat_A[11][3] * mat_B[3][20] +
                  mat_A[11][4] * mat_B[4][20] +
                  mat_A[11][5] * mat_B[5][20] +
                  mat_A[11][6] * mat_B[6][20] +
                  mat_A[11][7] * mat_B[7][20] +
                  mat_A[11][8] * mat_B[8][20] +
                  mat_A[11][9] * mat_B[9][20] +
                  mat_A[11][10] * mat_B[10][20] +
                  mat_A[11][11] * mat_B[11][20] +
                  mat_A[11][12] * mat_B[12][20] +
                  mat_A[11][13] * mat_B[13][20] +
                  mat_A[11][14] * mat_B[14][20] +
                  mat_A[11][15] * mat_B[15][20] +
                  mat_A[11][16] * mat_B[16][20] +
                  mat_A[11][17] * mat_B[17][20] +
                  mat_A[11][18] * mat_B[18][20] +
                  mat_A[11][19] * mat_B[19][20] +
                  mat_A[11][20] * mat_B[20][20] +
                  mat_A[11][21] * mat_B[21][20] +
                  mat_A[11][22] * mat_B[22][20] +
                  mat_A[11][23] * mat_B[23][20] +
                  mat_A[11][24] * mat_B[24][20] +
                  mat_A[11][25] * mat_B[25][20] +
                  mat_A[11][26] * mat_B[26][20] +
                  mat_A[11][27] * mat_B[27][20] +
                  mat_A[11][28] * mat_B[28][20] +
                  mat_A[11][29] * mat_B[29][20] +
                  mat_A[11][30] * mat_B[30][20] +
                  mat_A[11][31] * mat_B[31][20];
    mat_C[11][21] <= 
                  mat_A[11][0] * mat_B[0][21] +
                  mat_A[11][1] * mat_B[1][21] +
                  mat_A[11][2] * mat_B[2][21] +
                  mat_A[11][3] * mat_B[3][21] +
                  mat_A[11][4] * mat_B[4][21] +
                  mat_A[11][5] * mat_B[5][21] +
                  mat_A[11][6] * mat_B[6][21] +
                  mat_A[11][7] * mat_B[7][21] +
                  mat_A[11][8] * mat_B[8][21] +
                  mat_A[11][9] * mat_B[9][21] +
                  mat_A[11][10] * mat_B[10][21] +
                  mat_A[11][11] * mat_B[11][21] +
                  mat_A[11][12] * mat_B[12][21] +
                  mat_A[11][13] * mat_B[13][21] +
                  mat_A[11][14] * mat_B[14][21] +
                  mat_A[11][15] * mat_B[15][21] +
                  mat_A[11][16] * mat_B[16][21] +
                  mat_A[11][17] * mat_B[17][21] +
                  mat_A[11][18] * mat_B[18][21] +
                  mat_A[11][19] * mat_B[19][21] +
                  mat_A[11][20] * mat_B[20][21] +
                  mat_A[11][21] * mat_B[21][21] +
                  mat_A[11][22] * mat_B[22][21] +
                  mat_A[11][23] * mat_B[23][21] +
                  mat_A[11][24] * mat_B[24][21] +
                  mat_A[11][25] * mat_B[25][21] +
                  mat_A[11][26] * mat_B[26][21] +
                  mat_A[11][27] * mat_B[27][21] +
                  mat_A[11][28] * mat_B[28][21] +
                  mat_A[11][29] * mat_B[29][21] +
                  mat_A[11][30] * mat_B[30][21] +
                  mat_A[11][31] * mat_B[31][21];
    mat_C[11][22] <= 
                  mat_A[11][0] * mat_B[0][22] +
                  mat_A[11][1] * mat_B[1][22] +
                  mat_A[11][2] * mat_B[2][22] +
                  mat_A[11][3] * mat_B[3][22] +
                  mat_A[11][4] * mat_B[4][22] +
                  mat_A[11][5] * mat_B[5][22] +
                  mat_A[11][6] * mat_B[6][22] +
                  mat_A[11][7] * mat_B[7][22] +
                  mat_A[11][8] * mat_B[8][22] +
                  mat_A[11][9] * mat_B[9][22] +
                  mat_A[11][10] * mat_B[10][22] +
                  mat_A[11][11] * mat_B[11][22] +
                  mat_A[11][12] * mat_B[12][22] +
                  mat_A[11][13] * mat_B[13][22] +
                  mat_A[11][14] * mat_B[14][22] +
                  mat_A[11][15] * mat_B[15][22] +
                  mat_A[11][16] * mat_B[16][22] +
                  mat_A[11][17] * mat_B[17][22] +
                  mat_A[11][18] * mat_B[18][22] +
                  mat_A[11][19] * mat_B[19][22] +
                  mat_A[11][20] * mat_B[20][22] +
                  mat_A[11][21] * mat_B[21][22] +
                  mat_A[11][22] * mat_B[22][22] +
                  mat_A[11][23] * mat_B[23][22] +
                  mat_A[11][24] * mat_B[24][22] +
                  mat_A[11][25] * mat_B[25][22] +
                  mat_A[11][26] * mat_B[26][22] +
                  mat_A[11][27] * mat_B[27][22] +
                  mat_A[11][28] * mat_B[28][22] +
                  mat_A[11][29] * mat_B[29][22] +
                  mat_A[11][30] * mat_B[30][22] +
                  mat_A[11][31] * mat_B[31][22];
    mat_C[11][23] <= 
                  mat_A[11][0] * mat_B[0][23] +
                  mat_A[11][1] * mat_B[1][23] +
                  mat_A[11][2] * mat_B[2][23] +
                  mat_A[11][3] * mat_B[3][23] +
                  mat_A[11][4] * mat_B[4][23] +
                  mat_A[11][5] * mat_B[5][23] +
                  mat_A[11][6] * mat_B[6][23] +
                  mat_A[11][7] * mat_B[7][23] +
                  mat_A[11][8] * mat_B[8][23] +
                  mat_A[11][9] * mat_B[9][23] +
                  mat_A[11][10] * mat_B[10][23] +
                  mat_A[11][11] * mat_B[11][23] +
                  mat_A[11][12] * mat_B[12][23] +
                  mat_A[11][13] * mat_B[13][23] +
                  mat_A[11][14] * mat_B[14][23] +
                  mat_A[11][15] * mat_B[15][23] +
                  mat_A[11][16] * mat_B[16][23] +
                  mat_A[11][17] * mat_B[17][23] +
                  mat_A[11][18] * mat_B[18][23] +
                  mat_A[11][19] * mat_B[19][23] +
                  mat_A[11][20] * mat_B[20][23] +
                  mat_A[11][21] * mat_B[21][23] +
                  mat_A[11][22] * mat_B[22][23] +
                  mat_A[11][23] * mat_B[23][23] +
                  mat_A[11][24] * mat_B[24][23] +
                  mat_A[11][25] * mat_B[25][23] +
                  mat_A[11][26] * mat_B[26][23] +
                  mat_A[11][27] * mat_B[27][23] +
                  mat_A[11][28] * mat_B[28][23] +
                  mat_A[11][29] * mat_B[29][23] +
                  mat_A[11][30] * mat_B[30][23] +
                  mat_A[11][31] * mat_B[31][23];
    mat_C[11][24] <= 
                  mat_A[11][0] * mat_B[0][24] +
                  mat_A[11][1] * mat_B[1][24] +
                  mat_A[11][2] * mat_B[2][24] +
                  mat_A[11][3] * mat_B[3][24] +
                  mat_A[11][4] * mat_B[4][24] +
                  mat_A[11][5] * mat_B[5][24] +
                  mat_A[11][6] * mat_B[6][24] +
                  mat_A[11][7] * mat_B[7][24] +
                  mat_A[11][8] * mat_B[8][24] +
                  mat_A[11][9] * mat_B[9][24] +
                  mat_A[11][10] * mat_B[10][24] +
                  mat_A[11][11] * mat_B[11][24] +
                  mat_A[11][12] * mat_B[12][24] +
                  mat_A[11][13] * mat_B[13][24] +
                  mat_A[11][14] * mat_B[14][24] +
                  mat_A[11][15] * mat_B[15][24] +
                  mat_A[11][16] * mat_B[16][24] +
                  mat_A[11][17] * mat_B[17][24] +
                  mat_A[11][18] * mat_B[18][24] +
                  mat_A[11][19] * mat_B[19][24] +
                  mat_A[11][20] * mat_B[20][24] +
                  mat_A[11][21] * mat_B[21][24] +
                  mat_A[11][22] * mat_B[22][24] +
                  mat_A[11][23] * mat_B[23][24] +
                  mat_A[11][24] * mat_B[24][24] +
                  mat_A[11][25] * mat_B[25][24] +
                  mat_A[11][26] * mat_B[26][24] +
                  mat_A[11][27] * mat_B[27][24] +
                  mat_A[11][28] * mat_B[28][24] +
                  mat_A[11][29] * mat_B[29][24] +
                  mat_A[11][30] * mat_B[30][24] +
                  mat_A[11][31] * mat_B[31][24];
    mat_C[11][25] <= 
                  mat_A[11][0] * mat_B[0][25] +
                  mat_A[11][1] * mat_B[1][25] +
                  mat_A[11][2] * mat_B[2][25] +
                  mat_A[11][3] * mat_B[3][25] +
                  mat_A[11][4] * mat_B[4][25] +
                  mat_A[11][5] * mat_B[5][25] +
                  mat_A[11][6] * mat_B[6][25] +
                  mat_A[11][7] * mat_B[7][25] +
                  mat_A[11][8] * mat_B[8][25] +
                  mat_A[11][9] * mat_B[9][25] +
                  mat_A[11][10] * mat_B[10][25] +
                  mat_A[11][11] * mat_B[11][25] +
                  mat_A[11][12] * mat_B[12][25] +
                  mat_A[11][13] * mat_B[13][25] +
                  mat_A[11][14] * mat_B[14][25] +
                  mat_A[11][15] * mat_B[15][25] +
                  mat_A[11][16] * mat_B[16][25] +
                  mat_A[11][17] * mat_B[17][25] +
                  mat_A[11][18] * mat_B[18][25] +
                  mat_A[11][19] * mat_B[19][25] +
                  mat_A[11][20] * mat_B[20][25] +
                  mat_A[11][21] * mat_B[21][25] +
                  mat_A[11][22] * mat_B[22][25] +
                  mat_A[11][23] * mat_B[23][25] +
                  mat_A[11][24] * mat_B[24][25] +
                  mat_A[11][25] * mat_B[25][25] +
                  mat_A[11][26] * mat_B[26][25] +
                  mat_A[11][27] * mat_B[27][25] +
                  mat_A[11][28] * mat_B[28][25] +
                  mat_A[11][29] * mat_B[29][25] +
                  mat_A[11][30] * mat_B[30][25] +
                  mat_A[11][31] * mat_B[31][25];
    mat_C[11][26] <= 
                  mat_A[11][0] * mat_B[0][26] +
                  mat_A[11][1] * mat_B[1][26] +
                  mat_A[11][2] * mat_B[2][26] +
                  mat_A[11][3] * mat_B[3][26] +
                  mat_A[11][4] * mat_B[4][26] +
                  mat_A[11][5] * mat_B[5][26] +
                  mat_A[11][6] * mat_B[6][26] +
                  mat_A[11][7] * mat_B[7][26] +
                  mat_A[11][8] * mat_B[8][26] +
                  mat_A[11][9] * mat_B[9][26] +
                  mat_A[11][10] * mat_B[10][26] +
                  mat_A[11][11] * mat_B[11][26] +
                  mat_A[11][12] * mat_B[12][26] +
                  mat_A[11][13] * mat_B[13][26] +
                  mat_A[11][14] * mat_B[14][26] +
                  mat_A[11][15] * mat_B[15][26] +
                  mat_A[11][16] * mat_B[16][26] +
                  mat_A[11][17] * mat_B[17][26] +
                  mat_A[11][18] * mat_B[18][26] +
                  mat_A[11][19] * mat_B[19][26] +
                  mat_A[11][20] * mat_B[20][26] +
                  mat_A[11][21] * mat_B[21][26] +
                  mat_A[11][22] * mat_B[22][26] +
                  mat_A[11][23] * mat_B[23][26] +
                  mat_A[11][24] * mat_B[24][26] +
                  mat_A[11][25] * mat_B[25][26] +
                  mat_A[11][26] * mat_B[26][26] +
                  mat_A[11][27] * mat_B[27][26] +
                  mat_A[11][28] * mat_B[28][26] +
                  mat_A[11][29] * mat_B[29][26] +
                  mat_A[11][30] * mat_B[30][26] +
                  mat_A[11][31] * mat_B[31][26];
    mat_C[11][27] <= 
                  mat_A[11][0] * mat_B[0][27] +
                  mat_A[11][1] * mat_B[1][27] +
                  mat_A[11][2] * mat_B[2][27] +
                  mat_A[11][3] * mat_B[3][27] +
                  mat_A[11][4] * mat_B[4][27] +
                  mat_A[11][5] * mat_B[5][27] +
                  mat_A[11][6] * mat_B[6][27] +
                  mat_A[11][7] * mat_B[7][27] +
                  mat_A[11][8] * mat_B[8][27] +
                  mat_A[11][9] * mat_B[9][27] +
                  mat_A[11][10] * mat_B[10][27] +
                  mat_A[11][11] * mat_B[11][27] +
                  mat_A[11][12] * mat_B[12][27] +
                  mat_A[11][13] * mat_B[13][27] +
                  mat_A[11][14] * mat_B[14][27] +
                  mat_A[11][15] * mat_B[15][27] +
                  mat_A[11][16] * mat_B[16][27] +
                  mat_A[11][17] * mat_B[17][27] +
                  mat_A[11][18] * mat_B[18][27] +
                  mat_A[11][19] * mat_B[19][27] +
                  mat_A[11][20] * mat_B[20][27] +
                  mat_A[11][21] * mat_B[21][27] +
                  mat_A[11][22] * mat_B[22][27] +
                  mat_A[11][23] * mat_B[23][27] +
                  mat_A[11][24] * mat_B[24][27] +
                  mat_A[11][25] * mat_B[25][27] +
                  mat_A[11][26] * mat_B[26][27] +
                  mat_A[11][27] * mat_B[27][27] +
                  mat_A[11][28] * mat_B[28][27] +
                  mat_A[11][29] * mat_B[29][27] +
                  mat_A[11][30] * mat_B[30][27] +
                  mat_A[11][31] * mat_B[31][27];
    mat_C[11][28] <= 
                  mat_A[11][0] * mat_B[0][28] +
                  mat_A[11][1] * mat_B[1][28] +
                  mat_A[11][2] * mat_B[2][28] +
                  mat_A[11][3] * mat_B[3][28] +
                  mat_A[11][4] * mat_B[4][28] +
                  mat_A[11][5] * mat_B[5][28] +
                  mat_A[11][6] * mat_B[6][28] +
                  mat_A[11][7] * mat_B[7][28] +
                  mat_A[11][8] * mat_B[8][28] +
                  mat_A[11][9] * mat_B[9][28] +
                  mat_A[11][10] * mat_B[10][28] +
                  mat_A[11][11] * mat_B[11][28] +
                  mat_A[11][12] * mat_B[12][28] +
                  mat_A[11][13] * mat_B[13][28] +
                  mat_A[11][14] * mat_B[14][28] +
                  mat_A[11][15] * mat_B[15][28] +
                  mat_A[11][16] * mat_B[16][28] +
                  mat_A[11][17] * mat_B[17][28] +
                  mat_A[11][18] * mat_B[18][28] +
                  mat_A[11][19] * mat_B[19][28] +
                  mat_A[11][20] * mat_B[20][28] +
                  mat_A[11][21] * mat_B[21][28] +
                  mat_A[11][22] * mat_B[22][28] +
                  mat_A[11][23] * mat_B[23][28] +
                  mat_A[11][24] * mat_B[24][28] +
                  mat_A[11][25] * mat_B[25][28] +
                  mat_A[11][26] * mat_B[26][28] +
                  mat_A[11][27] * mat_B[27][28] +
                  mat_A[11][28] * mat_B[28][28] +
                  mat_A[11][29] * mat_B[29][28] +
                  mat_A[11][30] * mat_B[30][28] +
                  mat_A[11][31] * mat_B[31][28];
    mat_C[11][29] <= 
                  mat_A[11][0] * mat_B[0][29] +
                  mat_A[11][1] * mat_B[1][29] +
                  mat_A[11][2] * mat_B[2][29] +
                  mat_A[11][3] * mat_B[3][29] +
                  mat_A[11][4] * mat_B[4][29] +
                  mat_A[11][5] * mat_B[5][29] +
                  mat_A[11][6] * mat_B[6][29] +
                  mat_A[11][7] * mat_B[7][29] +
                  mat_A[11][8] * mat_B[8][29] +
                  mat_A[11][9] * mat_B[9][29] +
                  mat_A[11][10] * mat_B[10][29] +
                  mat_A[11][11] * mat_B[11][29] +
                  mat_A[11][12] * mat_B[12][29] +
                  mat_A[11][13] * mat_B[13][29] +
                  mat_A[11][14] * mat_B[14][29] +
                  mat_A[11][15] * mat_B[15][29] +
                  mat_A[11][16] * mat_B[16][29] +
                  mat_A[11][17] * mat_B[17][29] +
                  mat_A[11][18] * mat_B[18][29] +
                  mat_A[11][19] * mat_B[19][29] +
                  mat_A[11][20] * mat_B[20][29] +
                  mat_A[11][21] * mat_B[21][29] +
                  mat_A[11][22] * mat_B[22][29] +
                  mat_A[11][23] * mat_B[23][29] +
                  mat_A[11][24] * mat_B[24][29] +
                  mat_A[11][25] * mat_B[25][29] +
                  mat_A[11][26] * mat_B[26][29] +
                  mat_A[11][27] * mat_B[27][29] +
                  mat_A[11][28] * mat_B[28][29] +
                  mat_A[11][29] * mat_B[29][29] +
                  mat_A[11][30] * mat_B[30][29] +
                  mat_A[11][31] * mat_B[31][29];
    mat_C[11][30] <= 
                  mat_A[11][0] * mat_B[0][30] +
                  mat_A[11][1] * mat_B[1][30] +
                  mat_A[11][2] * mat_B[2][30] +
                  mat_A[11][3] * mat_B[3][30] +
                  mat_A[11][4] * mat_B[4][30] +
                  mat_A[11][5] * mat_B[5][30] +
                  mat_A[11][6] * mat_B[6][30] +
                  mat_A[11][7] * mat_B[7][30] +
                  mat_A[11][8] * mat_B[8][30] +
                  mat_A[11][9] * mat_B[9][30] +
                  mat_A[11][10] * mat_B[10][30] +
                  mat_A[11][11] * mat_B[11][30] +
                  mat_A[11][12] * mat_B[12][30] +
                  mat_A[11][13] * mat_B[13][30] +
                  mat_A[11][14] * mat_B[14][30] +
                  mat_A[11][15] * mat_B[15][30] +
                  mat_A[11][16] * mat_B[16][30] +
                  mat_A[11][17] * mat_B[17][30] +
                  mat_A[11][18] * mat_B[18][30] +
                  mat_A[11][19] * mat_B[19][30] +
                  mat_A[11][20] * mat_B[20][30] +
                  mat_A[11][21] * mat_B[21][30] +
                  mat_A[11][22] * mat_B[22][30] +
                  mat_A[11][23] * mat_B[23][30] +
                  mat_A[11][24] * mat_B[24][30] +
                  mat_A[11][25] * mat_B[25][30] +
                  mat_A[11][26] * mat_B[26][30] +
                  mat_A[11][27] * mat_B[27][30] +
                  mat_A[11][28] * mat_B[28][30] +
                  mat_A[11][29] * mat_B[29][30] +
                  mat_A[11][30] * mat_B[30][30] +
                  mat_A[11][31] * mat_B[31][30];
    mat_C[11][31] <= 
                  mat_A[11][0] * mat_B[0][31] +
                  mat_A[11][1] * mat_B[1][31] +
                  mat_A[11][2] * mat_B[2][31] +
                  mat_A[11][3] * mat_B[3][31] +
                  mat_A[11][4] * mat_B[4][31] +
                  mat_A[11][5] * mat_B[5][31] +
                  mat_A[11][6] * mat_B[6][31] +
                  mat_A[11][7] * mat_B[7][31] +
                  mat_A[11][8] * mat_B[8][31] +
                  mat_A[11][9] * mat_B[9][31] +
                  mat_A[11][10] * mat_B[10][31] +
                  mat_A[11][11] * mat_B[11][31] +
                  mat_A[11][12] * mat_B[12][31] +
                  mat_A[11][13] * mat_B[13][31] +
                  mat_A[11][14] * mat_B[14][31] +
                  mat_A[11][15] * mat_B[15][31] +
                  mat_A[11][16] * mat_B[16][31] +
                  mat_A[11][17] * mat_B[17][31] +
                  mat_A[11][18] * mat_B[18][31] +
                  mat_A[11][19] * mat_B[19][31] +
                  mat_A[11][20] * mat_B[20][31] +
                  mat_A[11][21] * mat_B[21][31] +
                  mat_A[11][22] * mat_B[22][31] +
                  mat_A[11][23] * mat_B[23][31] +
                  mat_A[11][24] * mat_B[24][31] +
                  mat_A[11][25] * mat_B[25][31] +
                  mat_A[11][26] * mat_B[26][31] +
                  mat_A[11][27] * mat_B[27][31] +
                  mat_A[11][28] * mat_B[28][31] +
                  mat_A[11][29] * mat_B[29][31] +
                  mat_A[11][30] * mat_B[30][31] +
                  mat_A[11][31] * mat_B[31][31];
    mat_C[12][0] <= 
                  mat_A[12][0] * mat_B[0][0] +
                  mat_A[12][1] * mat_B[1][0] +
                  mat_A[12][2] * mat_B[2][0] +
                  mat_A[12][3] * mat_B[3][0] +
                  mat_A[12][4] * mat_B[4][0] +
                  mat_A[12][5] * mat_B[5][0] +
                  mat_A[12][6] * mat_B[6][0] +
                  mat_A[12][7] * mat_B[7][0] +
                  mat_A[12][8] * mat_B[8][0] +
                  mat_A[12][9] * mat_B[9][0] +
                  mat_A[12][10] * mat_B[10][0] +
                  mat_A[12][11] * mat_B[11][0] +
                  mat_A[12][12] * mat_B[12][0] +
                  mat_A[12][13] * mat_B[13][0] +
                  mat_A[12][14] * mat_B[14][0] +
                  mat_A[12][15] * mat_B[15][0] +
                  mat_A[12][16] * mat_B[16][0] +
                  mat_A[12][17] * mat_B[17][0] +
                  mat_A[12][18] * mat_B[18][0] +
                  mat_A[12][19] * mat_B[19][0] +
                  mat_A[12][20] * mat_B[20][0] +
                  mat_A[12][21] * mat_B[21][0] +
                  mat_A[12][22] * mat_B[22][0] +
                  mat_A[12][23] * mat_B[23][0] +
                  mat_A[12][24] * mat_B[24][0] +
                  mat_A[12][25] * mat_B[25][0] +
                  mat_A[12][26] * mat_B[26][0] +
                  mat_A[12][27] * mat_B[27][0] +
                  mat_A[12][28] * mat_B[28][0] +
                  mat_A[12][29] * mat_B[29][0] +
                  mat_A[12][30] * mat_B[30][0] +
                  mat_A[12][31] * mat_B[31][0];
    mat_C[12][1] <= 
                  mat_A[12][0] * mat_B[0][1] +
                  mat_A[12][1] * mat_B[1][1] +
                  mat_A[12][2] * mat_B[2][1] +
                  mat_A[12][3] * mat_B[3][1] +
                  mat_A[12][4] * mat_B[4][1] +
                  mat_A[12][5] * mat_B[5][1] +
                  mat_A[12][6] * mat_B[6][1] +
                  mat_A[12][7] * mat_B[7][1] +
                  mat_A[12][8] * mat_B[8][1] +
                  mat_A[12][9] * mat_B[9][1] +
                  mat_A[12][10] * mat_B[10][1] +
                  mat_A[12][11] * mat_B[11][1] +
                  mat_A[12][12] * mat_B[12][1] +
                  mat_A[12][13] * mat_B[13][1] +
                  mat_A[12][14] * mat_B[14][1] +
                  mat_A[12][15] * mat_B[15][1] +
                  mat_A[12][16] * mat_B[16][1] +
                  mat_A[12][17] * mat_B[17][1] +
                  mat_A[12][18] * mat_B[18][1] +
                  mat_A[12][19] * mat_B[19][1] +
                  mat_A[12][20] * mat_B[20][1] +
                  mat_A[12][21] * mat_B[21][1] +
                  mat_A[12][22] * mat_B[22][1] +
                  mat_A[12][23] * mat_B[23][1] +
                  mat_A[12][24] * mat_B[24][1] +
                  mat_A[12][25] * mat_B[25][1] +
                  mat_A[12][26] * mat_B[26][1] +
                  mat_A[12][27] * mat_B[27][1] +
                  mat_A[12][28] * mat_B[28][1] +
                  mat_A[12][29] * mat_B[29][1] +
                  mat_A[12][30] * mat_B[30][1] +
                  mat_A[12][31] * mat_B[31][1];
    mat_C[12][2] <= 
                  mat_A[12][0] * mat_B[0][2] +
                  mat_A[12][1] * mat_B[1][2] +
                  mat_A[12][2] * mat_B[2][2] +
                  mat_A[12][3] * mat_B[3][2] +
                  mat_A[12][4] * mat_B[4][2] +
                  mat_A[12][5] * mat_B[5][2] +
                  mat_A[12][6] * mat_B[6][2] +
                  mat_A[12][7] * mat_B[7][2] +
                  mat_A[12][8] * mat_B[8][2] +
                  mat_A[12][9] * mat_B[9][2] +
                  mat_A[12][10] * mat_B[10][2] +
                  mat_A[12][11] * mat_B[11][2] +
                  mat_A[12][12] * mat_B[12][2] +
                  mat_A[12][13] * mat_B[13][2] +
                  mat_A[12][14] * mat_B[14][2] +
                  mat_A[12][15] * mat_B[15][2] +
                  mat_A[12][16] * mat_B[16][2] +
                  mat_A[12][17] * mat_B[17][2] +
                  mat_A[12][18] * mat_B[18][2] +
                  mat_A[12][19] * mat_B[19][2] +
                  mat_A[12][20] * mat_B[20][2] +
                  mat_A[12][21] * mat_B[21][2] +
                  mat_A[12][22] * mat_B[22][2] +
                  mat_A[12][23] * mat_B[23][2] +
                  mat_A[12][24] * mat_B[24][2] +
                  mat_A[12][25] * mat_B[25][2] +
                  mat_A[12][26] * mat_B[26][2] +
                  mat_A[12][27] * mat_B[27][2] +
                  mat_A[12][28] * mat_B[28][2] +
                  mat_A[12][29] * mat_B[29][2] +
                  mat_A[12][30] * mat_B[30][2] +
                  mat_A[12][31] * mat_B[31][2];
    mat_C[12][3] <= 
                  mat_A[12][0] * mat_B[0][3] +
                  mat_A[12][1] * mat_B[1][3] +
                  mat_A[12][2] * mat_B[2][3] +
                  mat_A[12][3] * mat_B[3][3] +
                  mat_A[12][4] * mat_B[4][3] +
                  mat_A[12][5] * mat_B[5][3] +
                  mat_A[12][6] * mat_B[6][3] +
                  mat_A[12][7] * mat_B[7][3] +
                  mat_A[12][8] * mat_B[8][3] +
                  mat_A[12][9] * mat_B[9][3] +
                  mat_A[12][10] * mat_B[10][3] +
                  mat_A[12][11] * mat_B[11][3] +
                  mat_A[12][12] * mat_B[12][3] +
                  mat_A[12][13] * mat_B[13][3] +
                  mat_A[12][14] * mat_B[14][3] +
                  mat_A[12][15] * mat_B[15][3] +
                  mat_A[12][16] * mat_B[16][3] +
                  mat_A[12][17] * mat_B[17][3] +
                  mat_A[12][18] * mat_B[18][3] +
                  mat_A[12][19] * mat_B[19][3] +
                  mat_A[12][20] * mat_B[20][3] +
                  mat_A[12][21] * mat_B[21][3] +
                  mat_A[12][22] * mat_B[22][3] +
                  mat_A[12][23] * mat_B[23][3] +
                  mat_A[12][24] * mat_B[24][3] +
                  mat_A[12][25] * mat_B[25][3] +
                  mat_A[12][26] * mat_B[26][3] +
                  mat_A[12][27] * mat_B[27][3] +
                  mat_A[12][28] * mat_B[28][3] +
                  mat_A[12][29] * mat_B[29][3] +
                  mat_A[12][30] * mat_B[30][3] +
                  mat_A[12][31] * mat_B[31][3];
    mat_C[12][4] <= 
                  mat_A[12][0] * mat_B[0][4] +
                  mat_A[12][1] * mat_B[1][4] +
                  mat_A[12][2] * mat_B[2][4] +
                  mat_A[12][3] * mat_B[3][4] +
                  mat_A[12][4] * mat_B[4][4] +
                  mat_A[12][5] * mat_B[5][4] +
                  mat_A[12][6] * mat_B[6][4] +
                  mat_A[12][7] * mat_B[7][4] +
                  mat_A[12][8] * mat_B[8][4] +
                  mat_A[12][9] * mat_B[9][4] +
                  mat_A[12][10] * mat_B[10][4] +
                  mat_A[12][11] * mat_B[11][4] +
                  mat_A[12][12] * mat_B[12][4] +
                  mat_A[12][13] * mat_B[13][4] +
                  mat_A[12][14] * mat_B[14][4] +
                  mat_A[12][15] * mat_B[15][4] +
                  mat_A[12][16] * mat_B[16][4] +
                  mat_A[12][17] * mat_B[17][4] +
                  mat_A[12][18] * mat_B[18][4] +
                  mat_A[12][19] * mat_B[19][4] +
                  mat_A[12][20] * mat_B[20][4] +
                  mat_A[12][21] * mat_B[21][4] +
                  mat_A[12][22] * mat_B[22][4] +
                  mat_A[12][23] * mat_B[23][4] +
                  mat_A[12][24] * mat_B[24][4] +
                  mat_A[12][25] * mat_B[25][4] +
                  mat_A[12][26] * mat_B[26][4] +
                  mat_A[12][27] * mat_B[27][4] +
                  mat_A[12][28] * mat_B[28][4] +
                  mat_A[12][29] * mat_B[29][4] +
                  mat_A[12][30] * mat_B[30][4] +
                  mat_A[12][31] * mat_B[31][4];
    mat_C[12][5] <= 
                  mat_A[12][0] * mat_B[0][5] +
                  mat_A[12][1] * mat_B[1][5] +
                  mat_A[12][2] * mat_B[2][5] +
                  mat_A[12][3] * mat_B[3][5] +
                  mat_A[12][4] * mat_B[4][5] +
                  mat_A[12][5] * mat_B[5][5] +
                  mat_A[12][6] * mat_B[6][5] +
                  mat_A[12][7] * mat_B[7][5] +
                  mat_A[12][8] * mat_B[8][5] +
                  mat_A[12][9] * mat_B[9][5] +
                  mat_A[12][10] * mat_B[10][5] +
                  mat_A[12][11] * mat_B[11][5] +
                  mat_A[12][12] * mat_B[12][5] +
                  mat_A[12][13] * mat_B[13][5] +
                  mat_A[12][14] * mat_B[14][5] +
                  mat_A[12][15] * mat_B[15][5] +
                  mat_A[12][16] * mat_B[16][5] +
                  mat_A[12][17] * mat_B[17][5] +
                  mat_A[12][18] * mat_B[18][5] +
                  mat_A[12][19] * mat_B[19][5] +
                  mat_A[12][20] * mat_B[20][5] +
                  mat_A[12][21] * mat_B[21][5] +
                  mat_A[12][22] * mat_B[22][5] +
                  mat_A[12][23] * mat_B[23][5] +
                  mat_A[12][24] * mat_B[24][5] +
                  mat_A[12][25] * mat_B[25][5] +
                  mat_A[12][26] * mat_B[26][5] +
                  mat_A[12][27] * mat_B[27][5] +
                  mat_A[12][28] * mat_B[28][5] +
                  mat_A[12][29] * mat_B[29][5] +
                  mat_A[12][30] * mat_B[30][5] +
                  mat_A[12][31] * mat_B[31][5];
    mat_C[12][6] <= 
                  mat_A[12][0] * mat_B[0][6] +
                  mat_A[12][1] * mat_B[1][6] +
                  mat_A[12][2] * mat_B[2][6] +
                  mat_A[12][3] * mat_B[3][6] +
                  mat_A[12][4] * mat_B[4][6] +
                  mat_A[12][5] * mat_B[5][6] +
                  mat_A[12][6] * mat_B[6][6] +
                  mat_A[12][7] * mat_B[7][6] +
                  mat_A[12][8] * mat_B[8][6] +
                  mat_A[12][9] * mat_B[9][6] +
                  mat_A[12][10] * mat_B[10][6] +
                  mat_A[12][11] * mat_B[11][6] +
                  mat_A[12][12] * mat_B[12][6] +
                  mat_A[12][13] * mat_B[13][6] +
                  mat_A[12][14] * mat_B[14][6] +
                  mat_A[12][15] * mat_B[15][6] +
                  mat_A[12][16] * mat_B[16][6] +
                  mat_A[12][17] * mat_B[17][6] +
                  mat_A[12][18] * mat_B[18][6] +
                  mat_A[12][19] * mat_B[19][6] +
                  mat_A[12][20] * mat_B[20][6] +
                  mat_A[12][21] * mat_B[21][6] +
                  mat_A[12][22] * mat_B[22][6] +
                  mat_A[12][23] * mat_B[23][6] +
                  mat_A[12][24] * mat_B[24][6] +
                  mat_A[12][25] * mat_B[25][6] +
                  mat_A[12][26] * mat_B[26][6] +
                  mat_A[12][27] * mat_B[27][6] +
                  mat_A[12][28] * mat_B[28][6] +
                  mat_A[12][29] * mat_B[29][6] +
                  mat_A[12][30] * mat_B[30][6] +
                  mat_A[12][31] * mat_B[31][6];
    mat_C[12][7] <= 
                  mat_A[12][0] * mat_B[0][7] +
                  mat_A[12][1] * mat_B[1][7] +
                  mat_A[12][2] * mat_B[2][7] +
                  mat_A[12][3] * mat_B[3][7] +
                  mat_A[12][4] * mat_B[4][7] +
                  mat_A[12][5] * mat_B[5][7] +
                  mat_A[12][6] * mat_B[6][7] +
                  mat_A[12][7] * mat_B[7][7] +
                  mat_A[12][8] * mat_B[8][7] +
                  mat_A[12][9] * mat_B[9][7] +
                  mat_A[12][10] * mat_B[10][7] +
                  mat_A[12][11] * mat_B[11][7] +
                  mat_A[12][12] * mat_B[12][7] +
                  mat_A[12][13] * mat_B[13][7] +
                  mat_A[12][14] * mat_B[14][7] +
                  mat_A[12][15] * mat_B[15][7] +
                  mat_A[12][16] * mat_B[16][7] +
                  mat_A[12][17] * mat_B[17][7] +
                  mat_A[12][18] * mat_B[18][7] +
                  mat_A[12][19] * mat_B[19][7] +
                  mat_A[12][20] * mat_B[20][7] +
                  mat_A[12][21] * mat_B[21][7] +
                  mat_A[12][22] * mat_B[22][7] +
                  mat_A[12][23] * mat_B[23][7] +
                  mat_A[12][24] * mat_B[24][7] +
                  mat_A[12][25] * mat_B[25][7] +
                  mat_A[12][26] * mat_B[26][7] +
                  mat_A[12][27] * mat_B[27][7] +
                  mat_A[12][28] * mat_B[28][7] +
                  mat_A[12][29] * mat_B[29][7] +
                  mat_A[12][30] * mat_B[30][7] +
                  mat_A[12][31] * mat_B[31][7];
    mat_C[12][8] <= 
                  mat_A[12][0] * mat_B[0][8] +
                  mat_A[12][1] * mat_B[1][8] +
                  mat_A[12][2] * mat_B[2][8] +
                  mat_A[12][3] * mat_B[3][8] +
                  mat_A[12][4] * mat_B[4][8] +
                  mat_A[12][5] * mat_B[5][8] +
                  mat_A[12][6] * mat_B[6][8] +
                  mat_A[12][7] * mat_B[7][8] +
                  mat_A[12][8] * mat_B[8][8] +
                  mat_A[12][9] * mat_B[9][8] +
                  mat_A[12][10] * mat_B[10][8] +
                  mat_A[12][11] * mat_B[11][8] +
                  mat_A[12][12] * mat_B[12][8] +
                  mat_A[12][13] * mat_B[13][8] +
                  mat_A[12][14] * mat_B[14][8] +
                  mat_A[12][15] * mat_B[15][8] +
                  mat_A[12][16] * mat_B[16][8] +
                  mat_A[12][17] * mat_B[17][8] +
                  mat_A[12][18] * mat_B[18][8] +
                  mat_A[12][19] * mat_B[19][8] +
                  mat_A[12][20] * mat_B[20][8] +
                  mat_A[12][21] * mat_B[21][8] +
                  mat_A[12][22] * mat_B[22][8] +
                  mat_A[12][23] * mat_B[23][8] +
                  mat_A[12][24] * mat_B[24][8] +
                  mat_A[12][25] * mat_B[25][8] +
                  mat_A[12][26] * mat_B[26][8] +
                  mat_A[12][27] * mat_B[27][8] +
                  mat_A[12][28] * mat_B[28][8] +
                  mat_A[12][29] * mat_B[29][8] +
                  mat_A[12][30] * mat_B[30][8] +
                  mat_A[12][31] * mat_B[31][8];
    mat_C[12][9] <= 
                  mat_A[12][0] * mat_B[0][9] +
                  mat_A[12][1] * mat_B[1][9] +
                  mat_A[12][2] * mat_B[2][9] +
                  mat_A[12][3] * mat_B[3][9] +
                  mat_A[12][4] * mat_B[4][9] +
                  mat_A[12][5] * mat_B[5][9] +
                  mat_A[12][6] * mat_B[6][9] +
                  mat_A[12][7] * mat_B[7][9] +
                  mat_A[12][8] * mat_B[8][9] +
                  mat_A[12][9] * mat_B[9][9] +
                  mat_A[12][10] * mat_B[10][9] +
                  mat_A[12][11] * mat_B[11][9] +
                  mat_A[12][12] * mat_B[12][9] +
                  mat_A[12][13] * mat_B[13][9] +
                  mat_A[12][14] * mat_B[14][9] +
                  mat_A[12][15] * mat_B[15][9] +
                  mat_A[12][16] * mat_B[16][9] +
                  mat_A[12][17] * mat_B[17][9] +
                  mat_A[12][18] * mat_B[18][9] +
                  mat_A[12][19] * mat_B[19][9] +
                  mat_A[12][20] * mat_B[20][9] +
                  mat_A[12][21] * mat_B[21][9] +
                  mat_A[12][22] * mat_B[22][9] +
                  mat_A[12][23] * mat_B[23][9] +
                  mat_A[12][24] * mat_B[24][9] +
                  mat_A[12][25] * mat_B[25][9] +
                  mat_A[12][26] * mat_B[26][9] +
                  mat_A[12][27] * mat_B[27][9] +
                  mat_A[12][28] * mat_B[28][9] +
                  mat_A[12][29] * mat_B[29][9] +
                  mat_A[12][30] * mat_B[30][9] +
                  mat_A[12][31] * mat_B[31][9];
    mat_C[12][10] <= 
                  mat_A[12][0] * mat_B[0][10] +
                  mat_A[12][1] * mat_B[1][10] +
                  mat_A[12][2] * mat_B[2][10] +
                  mat_A[12][3] * mat_B[3][10] +
                  mat_A[12][4] * mat_B[4][10] +
                  mat_A[12][5] * mat_B[5][10] +
                  mat_A[12][6] * mat_B[6][10] +
                  mat_A[12][7] * mat_B[7][10] +
                  mat_A[12][8] * mat_B[8][10] +
                  mat_A[12][9] * mat_B[9][10] +
                  mat_A[12][10] * mat_B[10][10] +
                  mat_A[12][11] * mat_B[11][10] +
                  mat_A[12][12] * mat_B[12][10] +
                  mat_A[12][13] * mat_B[13][10] +
                  mat_A[12][14] * mat_B[14][10] +
                  mat_A[12][15] * mat_B[15][10] +
                  mat_A[12][16] * mat_B[16][10] +
                  mat_A[12][17] * mat_B[17][10] +
                  mat_A[12][18] * mat_B[18][10] +
                  mat_A[12][19] * mat_B[19][10] +
                  mat_A[12][20] * mat_B[20][10] +
                  mat_A[12][21] * mat_B[21][10] +
                  mat_A[12][22] * mat_B[22][10] +
                  mat_A[12][23] * mat_B[23][10] +
                  mat_A[12][24] * mat_B[24][10] +
                  mat_A[12][25] * mat_B[25][10] +
                  mat_A[12][26] * mat_B[26][10] +
                  mat_A[12][27] * mat_B[27][10] +
                  mat_A[12][28] * mat_B[28][10] +
                  mat_A[12][29] * mat_B[29][10] +
                  mat_A[12][30] * mat_B[30][10] +
                  mat_A[12][31] * mat_B[31][10];
    mat_C[12][11] <= 
                  mat_A[12][0] * mat_B[0][11] +
                  mat_A[12][1] * mat_B[1][11] +
                  mat_A[12][2] * mat_B[2][11] +
                  mat_A[12][3] * mat_B[3][11] +
                  mat_A[12][4] * mat_B[4][11] +
                  mat_A[12][5] * mat_B[5][11] +
                  mat_A[12][6] * mat_B[6][11] +
                  mat_A[12][7] * mat_B[7][11] +
                  mat_A[12][8] * mat_B[8][11] +
                  mat_A[12][9] * mat_B[9][11] +
                  mat_A[12][10] * mat_B[10][11] +
                  mat_A[12][11] * mat_B[11][11] +
                  mat_A[12][12] * mat_B[12][11] +
                  mat_A[12][13] * mat_B[13][11] +
                  mat_A[12][14] * mat_B[14][11] +
                  mat_A[12][15] * mat_B[15][11] +
                  mat_A[12][16] * mat_B[16][11] +
                  mat_A[12][17] * mat_B[17][11] +
                  mat_A[12][18] * mat_B[18][11] +
                  mat_A[12][19] * mat_B[19][11] +
                  mat_A[12][20] * mat_B[20][11] +
                  mat_A[12][21] * mat_B[21][11] +
                  mat_A[12][22] * mat_B[22][11] +
                  mat_A[12][23] * mat_B[23][11] +
                  mat_A[12][24] * mat_B[24][11] +
                  mat_A[12][25] * mat_B[25][11] +
                  mat_A[12][26] * mat_B[26][11] +
                  mat_A[12][27] * mat_B[27][11] +
                  mat_A[12][28] * mat_B[28][11] +
                  mat_A[12][29] * mat_B[29][11] +
                  mat_A[12][30] * mat_B[30][11] +
                  mat_A[12][31] * mat_B[31][11];
    mat_C[12][12] <= 
                  mat_A[12][0] * mat_B[0][12] +
                  mat_A[12][1] * mat_B[1][12] +
                  mat_A[12][2] * mat_B[2][12] +
                  mat_A[12][3] * mat_B[3][12] +
                  mat_A[12][4] * mat_B[4][12] +
                  mat_A[12][5] * mat_B[5][12] +
                  mat_A[12][6] * mat_B[6][12] +
                  mat_A[12][7] * mat_B[7][12] +
                  mat_A[12][8] * mat_B[8][12] +
                  mat_A[12][9] * mat_B[9][12] +
                  mat_A[12][10] * mat_B[10][12] +
                  mat_A[12][11] * mat_B[11][12] +
                  mat_A[12][12] * mat_B[12][12] +
                  mat_A[12][13] * mat_B[13][12] +
                  mat_A[12][14] * mat_B[14][12] +
                  mat_A[12][15] * mat_B[15][12] +
                  mat_A[12][16] * mat_B[16][12] +
                  mat_A[12][17] * mat_B[17][12] +
                  mat_A[12][18] * mat_B[18][12] +
                  mat_A[12][19] * mat_B[19][12] +
                  mat_A[12][20] * mat_B[20][12] +
                  mat_A[12][21] * mat_B[21][12] +
                  mat_A[12][22] * mat_B[22][12] +
                  mat_A[12][23] * mat_B[23][12] +
                  mat_A[12][24] * mat_B[24][12] +
                  mat_A[12][25] * mat_B[25][12] +
                  mat_A[12][26] * mat_B[26][12] +
                  mat_A[12][27] * mat_B[27][12] +
                  mat_A[12][28] * mat_B[28][12] +
                  mat_A[12][29] * mat_B[29][12] +
                  mat_A[12][30] * mat_B[30][12] +
                  mat_A[12][31] * mat_B[31][12];
    mat_C[12][13] <= 
                  mat_A[12][0] * mat_B[0][13] +
                  mat_A[12][1] * mat_B[1][13] +
                  mat_A[12][2] * mat_B[2][13] +
                  mat_A[12][3] * mat_B[3][13] +
                  mat_A[12][4] * mat_B[4][13] +
                  mat_A[12][5] * mat_B[5][13] +
                  mat_A[12][6] * mat_B[6][13] +
                  mat_A[12][7] * mat_B[7][13] +
                  mat_A[12][8] * mat_B[8][13] +
                  mat_A[12][9] * mat_B[9][13] +
                  mat_A[12][10] * mat_B[10][13] +
                  mat_A[12][11] * mat_B[11][13] +
                  mat_A[12][12] * mat_B[12][13] +
                  mat_A[12][13] * mat_B[13][13] +
                  mat_A[12][14] * mat_B[14][13] +
                  mat_A[12][15] * mat_B[15][13] +
                  mat_A[12][16] * mat_B[16][13] +
                  mat_A[12][17] * mat_B[17][13] +
                  mat_A[12][18] * mat_B[18][13] +
                  mat_A[12][19] * mat_B[19][13] +
                  mat_A[12][20] * mat_B[20][13] +
                  mat_A[12][21] * mat_B[21][13] +
                  mat_A[12][22] * mat_B[22][13] +
                  mat_A[12][23] * mat_B[23][13] +
                  mat_A[12][24] * mat_B[24][13] +
                  mat_A[12][25] * mat_B[25][13] +
                  mat_A[12][26] * mat_B[26][13] +
                  mat_A[12][27] * mat_B[27][13] +
                  mat_A[12][28] * mat_B[28][13] +
                  mat_A[12][29] * mat_B[29][13] +
                  mat_A[12][30] * mat_B[30][13] +
                  mat_A[12][31] * mat_B[31][13];
    mat_C[12][14] <= 
                  mat_A[12][0] * mat_B[0][14] +
                  mat_A[12][1] * mat_B[1][14] +
                  mat_A[12][2] * mat_B[2][14] +
                  mat_A[12][3] * mat_B[3][14] +
                  mat_A[12][4] * mat_B[4][14] +
                  mat_A[12][5] * mat_B[5][14] +
                  mat_A[12][6] * mat_B[6][14] +
                  mat_A[12][7] * mat_B[7][14] +
                  mat_A[12][8] * mat_B[8][14] +
                  mat_A[12][9] * mat_B[9][14] +
                  mat_A[12][10] * mat_B[10][14] +
                  mat_A[12][11] * mat_B[11][14] +
                  mat_A[12][12] * mat_B[12][14] +
                  mat_A[12][13] * mat_B[13][14] +
                  mat_A[12][14] * mat_B[14][14] +
                  mat_A[12][15] * mat_B[15][14] +
                  mat_A[12][16] * mat_B[16][14] +
                  mat_A[12][17] * mat_B[17][14] +
                  mat_A[12][18] * mat_B[18][14] +
                  mat_A[12][19] * mat_B[19][14] +
                  mat_A[12][20] * mat_B[20][14] +
                  mat_A[12][21] * mat_B[21][14] +
                  mat_A[12][22] * mat_B[22][14] +
                  mat_A[12][23] * mat_B[23][14] +
                  mat_A[12][24] * mat_B[24][14] +
                  mat_A[12][25] * mat_B[25][14] +
                  mat_A[12][26] * mat_B[26][14] +
                  mat_A[12][27] * mat_B[27][14] +
                  mat_A[12][28] * mat_B[28][14] +
                  mat_A[12][29] * mat_B[29][14] +
                  mat_A[12][30] * mat_B[30][14] +
                  mat_A[12][31] * mat_B[31][14];
    mat_C[12][15] <= 
                  mat_A[12][0] * mat_B[0][15] +
                  mat_A[12][1] * mat_B[1][15] +
                  mat_A[12][2] * mat_B[2][15] +
                  mat_A[12][3] * mat_B[3][15] +
                  mat_A[12][4] * mat_B[4][15] +
                  mat_A[12][5] * mat_B[5][15] +
                  mat_A[12][6] * mat_B[6][15] +
                  mat_A[12][7] * mat_B[7][15] +
                  mat_A[12][8] * mat_B[8][15] +
                  mat_A[12][9] * mat_B[9][15] +
                  mat_A[12][10] * mat_B[10][15] +
                  mat_A[12][11] * mat_B[11][15] +
                  mat_A[12][12] * mat_B[12][15] +
                  mat_A[12][13] * mat_B[13][15] +
                  mat_A[12][14] * mat_B[14][15] +
                  mat_A[12][15] * mat_B[15][15] +
                  mat_A[12][16] * mat_B[16][15] +
                  mat_A[12][17] * mat_B[17][15] +
                  mat_A[12][18] * mat_B[18][15] +
                  mat_A[12][19] * mat_B[19][15] +
                  mat_A[12][20] * mat_B[20][15] +
                  mat_A[12][21] * mat_B[21][15] +
                  mat_A[12][22] * mat_B[22][15] +
                  mat_A[12][23] * mat_B[23][15] +
                  mat_A[12][24] * mat_B[24][15] +
                  mat_A[12][25] * mat_B[25][15] +
                  mat_A[12][26] * mat_B[26][15] +
                  mat_A[12][27] * mat_B[27][15] +
                  mat_A[12][28] * mat_B[28][15] +
                  mat_A[12][29] * mat_B[29][15] +
                  mat_A[12][30] * mat_B[30][15] +
                  mat_A[12][31] * mat_B[31][15];
    mat_C[12][16] <= 
                  mat_A[12][0] * mat_B[0][16] +
                  mat_A[12][1] * mat_B[1][16] +
                  mat_A[12][2] * mat_B[2][16] +
                  mat_A[12][3] * mat_B[3][16] +
                  mat_A[12][4] * mat_B[4][16] +
                  mat_A[12][5] * mat_B[5][16] +
                  mat_A[12][6] * mat_B[6][16] +
                  mat_A[12][7] * mat_B[7][16] +
                  mat_A[12][8] * mat_B[8][16] +
                  mat_A[12][9] * mat_B[9][16] +
                  mat_A[12][10] * mat_B[10][16] +
                  mat_A[12][11] * mat_B[11][16] +
                  mat_A[12][12] * mat_B[12][16] +
                  mat_A[12][13] * mat_B[13][16] +
                  mat_A[12][14] * mat_B[14][16] +
                  mat_A[12][15] * mat_B[15][16] +
                  mat_A[12][16] * mat_B[16][16] +
                  mat_A[12][17] * mat_B[17][16] +
                  mat_A[12][18] * mat_B[18][16] +
                  mat_A[12][19] * mat_B[19][16] +
                  mat_A[12][20] * mat_B[20][16] +
                  mat_A[12][21] * mat_B[21][16] +
                  mat_A[12][22] * mat_B[22][16] +
                  mat_A[12][23] * mat_B[23][16] +
                  mat_A[12][24] * mat_B[24][16] +
                  mat_A[12][25] * mat_B[25][16] +
                  mat_A[12][26] * mat_B[26][16] +
                  mat_A[12][27] * mat_B[27][16] +
                  mat_A[12][28] * mat_B[28][16] +
                  mat_A[12][29] * mat_B[29][16] +
                  mat_A[12][30] * mat_B[30][16] +
                  mat_A[12][31] * mat_B[31][16];
    mat_C[12][17] <= 
                  mat_A[12][0] * mat_B[0][17] +
                  mat_A[12][1] * mat_B[1][17] +
                  mat_A[12][2] * mat_B[2][17] +
                  mat_A[12][3] * mat_B[3][17] +
                  mat_A[12][4] * mat_B[4][17] +
                  mat_A[12][5] * mat_B[5][17] +
                  mat_A[12][6] * mat_B[6][17] +
                  mat_A[12][7] * mat_B[7][17] +
                  mat_A[12][8] * mat_B[8][17] +
                  mat_A[12][9] * mat_B[9][17] +
                  mat_A[12][10] * mat_B[10][17] +
                  mat_A[12][11] * mat_B[11][17] +
                  mat_A[12][12] * mat_B[12][17] +
                  mat_A[12][13] * mat_B[13][17] +
                  mat_A[12][14] * mat_B[14][17] +
                  mat_A[12][15] * mat_B[15][17] +
                  mat_A[12][16] * mat_B[16][17] +
                  mat_A[12][17] * mat_B[17][17] +
                  mat_A[12][18] * mat_B[18][17] +
                  mat_A[12][19] * mat_B[19][17] +
                  mat_A[12][20] * mat_B[20][17] +
                  mat_A[12][21] * mat_B[21][17] +
                  mat_A[12][22] * mat_B[22][17] +
                  mat_A[12][23] * mat_B[23][17] +
                  mat_A[12][24] * mat_B[24][17] +
                  mat_A[12][25] * mat_B[25][17] +
                  mat_A[12][26] * mat_B[26][17] +
                  mat_A[12][27] * mat_B[27][17] +
                  mat_A[12][28] * mat_B[28][17] +
                  mat_A[12][29] * mat_B[29][17] +
                  mat_A[12][30] * mat_B[30][17] +
                  mat_A[12][31] * mat_B[31][17];
    mat_C[12][18] <= 
                  mat_A[12][0] * mat_B[0][18] +
                  mat_A[12][1] * mat_B[1][18] +
                  mat_A[12][2] * mat_B[2][18] +
                  mat_A[12][3] * mat_B[3][18] +
                  mat_A[12][4] * mat_B[4][18] +
                  mat_A[12][5] * mat_B[5][18] +
                  mat_A[12][6] * mat_B[6][18] +
                  mat_A[12][7] * mat_B[7][18] +
                  mat_A[12][8] * mat_B[8][18] +
                  mat_A[12][9] * mat_B[9][18] +
                  mat_A[12][10] * mat_B[10][18] +
                  mat_A[12][11] * mat_B[11][18] +
                  mat_A[12][12] * mat_B[12][18] +
                  mat_A[12][13] * mat_B[13][18] +
                  mat_A[12][14] * mat_B[14][18] +
                  mat_A[12][15] * mat_B[15][18] +
                  mat_A[12][16] * mat_B[16][18] +
                  mat_A[12][17] * mat_B[17][18] +
                  mat_A[12][18] * mat_B[18][18] +
                  mat_A[12][19] * mat_B[19][18] +
                  mat_A[12][20] * mat_B[20][18] +
                  mat_A[12][21] * mat_B[21][18] +
                  mat_A[12][22] * mat_B[22][18] +
                  mat_A[12][23] * mat_B[23][18] +
                  mat_A[12][24] * mat_B[24][18] +
                  mat_A[12][25] * mat_B[25][18] +
                  mat_A[12][26] * mat_B[26][18] +
                  mat_A[12][27] * mat_B[27][18] +
                  mat_A[12][28] * mat_B[28][18] +
                  mat_A[12][29] * mat_B[29][18] +
                  mat_A[12][30] * mat_B[30][18] +
                  mat_A[12][31] * mat_B[31][18];
    mat_C[12][19] <= 
                  mat_A[12][0] * mat_B[0][19] +
                  mat_A[12][1] * mat_B[1][19] +
                  mat_A[12][2] * mat_B[2][19] +
                  mat_A[12][3] * mat_B[3][19] +
                  mat_A[12][4] * mat_B[4][19] +
                  mat_A[12][5] * mat_B[5][19] +
                  mat_A[12][6] * mat_B[6][19] +
                  mat_A[12][7] * mat_B[7][19] +
                  mat_A[12][8] * mat_B[8][19] +
                  mat_A[12][9] * mat_B[9][19] +
                  mat_A[12][10] * mat_B[10][19] +
                  mat_A[12][11] * mat_B[11][19] +
                  mat_A[12][12] * mat_B[12][19] +
                  mat_A[12][13] * mat_B[13][19] +
                  mat_A[12][14] * mat_B[14][19] +
                  mat_A[12][15] * mat_B[15][19] +
                  mat_A[12][16] * mat_B[16][19] +
                  mat_A[12][17] * mat_B[17][19] +
                  mat_A[12][18] * mat_B[18][19] +
                  mat_A[12][19] * mat_B[19][19] +
                  mat_A[12][20] * mat_B[20][19] +
                  mat_A[12][21] * mat_B[21][19] +
                  mat_A[12][22] * mat_B[22][19] +
                  mat_A[12][23] * mat_B[23][19] +
                  mat_A[12][24] * mat_B[24][19] +
                  mat_A[12][25] * mat_B[25][19] +
                  mat_A[12][26] * mat_B[26][19] +
                  mat_A[12][27] * mat_B[27][19] +
                  mat_A[12][28] * mat_B[28][19] +
                  mat_A[12][29] * mat_B[29][19] +
                  mat_A[12][30] * mat_B[30][19] +
                  mat_A[12][31] * mat_B[31][19];
    mat_C[12][20] <= 
                  mat_A[12][0] * mat_B[0][20] +
                  mat_A[12][1] * mat_B[1][20] +
                  mat_A[12][2] * mat_B[2][20] +
                  mat_A[12][3] * mat_B[3][20] +
                  mat_A[12][4] * mat_B[4][20] +
                  mat_A[12][5] * mat_B[5][20] +
                  mat_A[12][6] * mat_B[6][20] +
                  mat_A[12][7] * mat_B[7][20] +
                  mat_A[12][8] * mat_B[8][20] +
                  mat_A[12][9] * mat_B[9][20] +
                  mat_A[12][10] * mat_B[10][20] +
                  mat_A[12][11] * mat_B[11][20] +
                  mat_A[12][12] * mat_B[12][20] +
                  mat_A[12][13] * mat_B[13][20] +
                  mat_A[12][14] * mat_B[14][20] +
                  mat_A[12][15] * mat_B[15][20] +
                  mat_A[12][16] * mat_B[16][20] +
                  mat_A[12][17] * mat_B[17][20] +
                  mat_A[12][18] * mat_B[18][20] +
                  mat_A[12][19] * mat_B[19][20] +
                  mat_A[12][20] * mat_B[20][20] +
                  mat_A[12][21] * mat_B[21][20] +
                  mat_A[12][22] * mat_B[22][20] +
                  mat_A[12][23] * mat_B[23][20] +
                  mat_A[12][24] * mat_B[24][20] +
                  mat_A[12][25] * mat_B[25][20] +
                  mat_A[12][26] * mat_B[26][20] +
                  mat_A[12][27] * mat_B[27][20] +
                  mat_A[12][28] * mat_B[28][20] +
                  mat_A[12][29] * mat_B[29][20] +
                  mat_A[12][30] * mat_B[30][20] +
                  mat_A[12][31] * mat_B[31][20];
    mat_C[12][21] <= 
                  mat_A[12][0] * mat_B[0][21] +
                  mat_A[12][1] * mat_B[1][21] +
                  mat_A[12][2] * mat_B[2][21] +
                  mat_A[12][3] * mat_B[3][21] +
                  mat_A[12][4] * mat_B[4][21] +
                  mat_A[12][5] * mat_B[5][21] +
                  mat_A[12][6] * mat_B[6][21] +
                  mat_A[12][7] * mat_B[7][21] +
                  mat_A[12][8] * mat_B[8][21] +
                  mat_A[12][9] * mat_B[9][21] +
                  mat_A[12][10] * mat_B[10][21] +
                  mat_A[12][11] * mat_B[11][21] +
                  mat_A[12][12] * mat_B[12][21] +
                  mat_A[12][13] * mat_B[13][21] +
                  mat_A[12][14] * mat_B[14][21] +
                  mat_A[12][15] * mat_B[15][21] +
                  mat_A[12][16] * mat_B[16][21] +
                  mat_A[12][17] * mat_B[17][21] +
                  mat_A[12][18] * mat_B[18][21] +
                  mat_A[12][19] * mat_B[19][21] +
                  mat_A[12][20] * mat_B[20][21] +
                  mat_A[12][21] * mat_B[21][21] +
                  mat_A[12][22] * mat_B[22][21] +
                  mat_A[12][23] * mat_B[23][21] +
                  mat_A[12][24] * mat_B[24][21] +
                  mat_A[12][25] * mat_B[25][21] +
                  mat_A[12][26] * mat_B[26][21] +
                  mat_A[12][27] * mat_B[27][21] +
                  mat_A[12][28] * mat_B[28][21] +
                  mat_A[12][29] * mat_B[29][21] +
                  mat_A[12][30] * mat_B[30][21] +
                  mat_A[12][31] * mat_B[31][21];
    mat_C[12][22] <= 
                  mat_A[12][0] * mat_B[0][22] +
                  mat_A[12][1] * mat_B[1][22] +
                  mat_A[12][2] * mat_B[2][22] +
                  mat_A[12][3] * mat_B[3][22] +
                  mat_A[12][4] * mat_B[4][22] +
                  mat_A[12][5] * mat_B[5][22] +
                  mat_A[12][6] * mat_B[6][22] +
                  mat_A[12][7] * mat_B[7][22] +
                  mat_A[12][8] * mat_B[8][22] +
                  mat_A[12][9] * mat_B[9][22] +
                  mat_A[12][10] * mat_B[10][22] +
                  mat_A[12][11] * mat_B[11][22] +
                  mat_A[12][12] * mat_B[12][22] +
                  mat_A[12][13] * mat_B[13][22] +
                  mat_A[12][14] * mat_B[14][22] +
                  mat_A[12][15] * mat_B[15][22] +
                  mat_A[12][16] * mat_B[16][22] +
                  mat_A[12][17] * mat_B[17][22] +
                  mat_A[12][18] * mat_B[18][22] +
                  mat_A[12][19] * mat_B[19][22] +
                  mat_A[12][20] * mat_B[20][22] +
                  mat_A[12][21] * mat_B[21][22] +
                  mat_A[12][22] * mat_B[22][22] +
                  mat_A[12][23] * mat_B[23][22] +
                  mat_A[12][24] * mat_B[24][22] +
                  mat_A[12][25] * mat_B[25][22] +
                  mat_A[12][26] * mat_B[26][22] +
                  mat_A[12][27] * mat_B[27][22] +
                  mat_A[12][28] * mat_B[28][22] +
                  mat_A[12][29] * mat_B[29][22] +
                  mat_A[12][30] * mat_B[30][22] +
                  mat_A[12][31] * mat_B[31][22];
    mat_C[12][23] <= 
                  mat_A[12][0] * mat_B[0][23] +
                  mat_A[12][1] * mat_B[1][23] +
                  mat_A[12][2] * mat_B[2][23] +
                  mat_A[12][3] * mat_B[3][23] +
                  mat_A[12][4] * mat_B[4][23] +
                  mat_A[12][5] * mat_B[5][23] +
                  mat_A[12][6] * mat_B[6][23] +
                  mat_A[12][7] * mat_B[7][23] +
                  mat_A[12][8] * mat_B[8][23] +
                  mat_A[12][9] * mat_B[9][23] +
                  mat_A[12][10] * mat_B[10][23] +
                  mat_A[12][11] * mat_B[11][23] +
                  mat_A[12][12] * mat_B[12][23] +
                  mat_A[12][13] * mat_B[13][23] +
                  mat_A[12][14] * mat_B[14][23] +
                  mat_A[12][15] * mat_B[15][23] +
                  mat_A[12][16] * mat_B[16][23] +
                  mat_A[12][17] * mat_B[17][23] +
                  mat_A[12][18] * mat_B[18][23] +
                  mat_A[12][19] * mat_B[19][23] +
                  mat_A[12][20] * mat_B[20][23] +
                  mat_A[12][21] * mat_B[21][23] +
                  mat_A[12][22] * mat_B[22][23] +
                  mat_A[12][23] * mat_B[23][23] +
                  mat_A[12][24] * mat_B[24][23] +
                  mat_A[12][25] * mat_B[25][23] +
                  mat_A[12][26] * mat_B[26][23] +
                  mat_A[12][27] * mat_B[27][23] +
                  mat_A[12][28] * mat_B[28][23] +
                  mat_A[12][29] * mat_B[29][23] +
                  mat_A[12][30] * mat_B[30][23] +
                  mat_A[12][31] * mat_B[31][23];
    mat_C[12][24] <= 
                  mat_A[12][0] * mat_B[0][24] +
                  mat_A[12][1] * mat_B[1][24] +
                  mat_A[12][2] * mat_B[2][24] +
                  mat_A[12][3] * mat_B[3][24] +
                  mat_A[12][4] * mat_B[4][24] +
                  mat_A[12][5] * mat_B[5][24] +
                  mat_A[12][6] * mat_B[6][24] +
                  mat_A[12][7] * mat_B[7][24] +
                  mat_A[12][8] * mat_B[8][24] +
                  mat_A[12][9] * mat_B[9][24] +
                  mat_A[12][10] * mat_B[10][24] +
                  mat_A[12][11] * mat_B[11][24] +
                  mat_A[12][12] * mat_B[12][24] +
                  mat_A[12][13] * mat_B[13][24] +
                  mat_A[12][14] * mat_B[14][24] +
                  mat_A[12][15] * mat_B[15][24] +
                  mat_A[12][16] * mat_B[16][24] +
                  mat_A[12][17] * mat_B[17][24] +
                  mat_A[12][18] * mat_B[18][24] +
                  mat_A[12][19] * mat_B[19][24] +
                  mat_A[12][20] * mat_B[20][24] +
                  mat_A[12][21] * mat_B[21][24] +
                  mat_A[12][22] * mat_B[22][24] +
                  mat_A[12][23] * mat_B[23][24] +
                  mat_A[12][24] * mat_B[24][24] +
                  mat_A[12][25] * mat_B[25][24] +
                  mat_A[12][26] * mat_B[26][24] +
                  mat_A[12][27] * mat_B[27][24] +
                  mat_A[12][28] * mat_B[28][24] +
                  mat_A[12][29] * mat_B[29][24] +
                  mat_A[12][30] * mat_B[30][24] +
                  mat_A[12][31] * mat_B[31][24];
    mat_C[12][25] <= 
                  mat_A[12][0] * mat_B[0][25] +
                  mat_A[12][1] * mat_B[1][25] +
                  mat_A[12][2] * mat_B[2][25] +
                  mat_A[12][3] * mat_B[3][25] +
                  mat_A[12][4] * mat_B[4][25] +
                  mat_A[12][5] * mat_B[5][25] +
                  mat_A[12][6] * mat_B[6][25] +
                  mat_A[12][7] * mat_B[7][25] +
                  mat_A[12][8] * mat_B[8][25] +
                  mat_A[12][9] * mat_B[9][25] +
                  mat_A[12][10] * mat_B[10][25] +
                  mat_A[12][11] * mat_B[11][25] +
                  mat_A[12][12] * mat_B[12][25] +
                  mat_A[12][13] * mat_B[13][25] +
                  mat_A[12][14] * mat_B[14][25] +
                  mat_A[12][15] * mat_B[15][25] +
                  mat_A[12][16] * mat_B[16][25] +
                  mat_A[12][17] * mat_B[17][25] +
                  mat_A[12][18] * mat_B[18][25] +
                  mat_A[12][19] * mat_B[19][25] +
                  mat_A[12][20] * mat_B[20][25] +
                  mat_A[12][21] * mat_B[21][25] +
                  mat_A[12][22] * mat_B[22][25] +
                  mat_A[12][23] * mat_B[23][25] +
                  mat_A[12][24] * mat_B[24][25] +
                  mat_A[12][25] * mat_B[25][25] +
                  mat_A[12][26] * mat_B[26][25] +
                  mat_A[12][27] * mat_B[27][25] +
                  mat_A[12][28] * mat_B[28][25] +
                  mat_A[12][29] * mat_B[29][25] +
                  mat_A[12][30] * mat_B[30][25] +
                  mat_A[12][31] * mat_B[31][25];
    mat_C[12][26] <= 
                  mat_A[12][0] * mat_B[0][26] +
                  mat_A[12][1] * mat_B[1][26] +
                  mat_A[12][2] * mat_B[2][26] +
                  mat_A[12][3] * mat_B[3][26] +
                  mat_A[12][4] * mat_B[4][26] +
                  mat_A[12][5] * mat_B[5][26] +
                  mat_A[12][6] * mat_B[6][26] +
                  mat_A[12][7] * mat_B[7][26] +
                  mat_A[12][8] * mat_B[8][26] +
                  mat_A[12][9] * mat_B[9][26] +
                  mat_A[12][10] * mat_B[10][26] +
                  mat_A[12][11] * mat_B[11][26] +
                  mat_A[12][12] * mat_B[12][26] +
                  mat_A[12][13] * mat_B[13][26] +
                  mat_A[12][14] * mat_B[14][26] +
                  mat_A[12][15] * mat_B[15][26] +
                  mat_A[12][16] * mat_B[16][26] +
                  mat_A[12][17] * mat_B[17][26] +
                  mat_A[12][18] * mat_B[18][26] +
                  mat_A[12][19] * mat_B[19][26] +
                  mat_A[12][20] * mat_B[20][26] +
                  mat_A[12][21] * mat_B[21][26] +
                  mat_A[12][22] * mat_B[22][26] +
                  mat_A[12][23] * mat_B[23][26] +
                  mat_A[12][24] * mat_B[24][26] +
                  mat_A[12][25] * mat_B[25][26] +
                  mat_A[12][26] * mat_B[26][26] +
                  mat_A[12][27] * mat_B[27][26] +
                  mat_A[12][28] * mat_B[28][26] +
                  mat_A[12][29] * mat_B[29][26] +
                  mat_A[12][30] * mat_B[30][26] +
                  mat_A[12][31] * mat_B[31][26];
    mat_C[12][27] <= 
                  mat_A[12][0] * mat_B[0][27] +
                  mat_A[12][1] * mat_B[1][27] +
                  mat_A[12][2] * mat_B[2][27] +
                  mat_A[12][3] * mat_B[3][27] +
                  mat_A[12][4] * mat_B[4][27] +
                  mat_A[12][5] * mat_B[5][27] +
                  mat_A[12][6] * mat_B[6][27] +
                  mat_A[12][7] * mat_B[7][27] +
                  mat_A[12][8] * mat_B[8][27] +
                  mat_A[12][9] * mat_B[9][27] +
                  mat_A[12][10] * mat_B[10][27] +
                  mat_A[12][11] * mat_B[11][27] +
                  mat_A[12][12] * mat_B[12][27] +
                  mat_A[12][13] * mat_B[13][27] +
                  mat_A[12][14] * mat_B[14][27] +
                  mat_A[12][15] * mat_B[15][27] +
                  mat_A[12][16] * mat_B[16][27] +
                  mat_A[12][17] * mat_B[17][27] +
                  mat_A[12][18] * mat_B[18][27] +
                  mat_A[12][19] * mat_B[19][27] +
                  mat_A[12][20] * mat_B[20][27] +
                  mat_A[12][21] * mat_B[21][27] +
                  mat_A[12][22] * mat_B[22][27] +
                  mat_A[12][23] * mat_B[23][27] +
                  mat_A[12][24] * mat_B[24][27] +
                  mat_A[12][25] * mat_B[25][27] +
                  mat_A[12][26] * mat_B[26][27] +
                  mat_A[12][27] * mat_B[27][27] +
                  mat_A[12][28] * mat_B[28][27] +
                  mat_A[12][29] * mat_B[29][27] +
                  mat_A[12][30] * mat_B[30][27] +
                  mat_A[12][31] * mat_B[31][27];
    mat_C[12][28] <= 
                  mat_A[12][0] * mat_B[0][28] +
                  mat_A[12][1] * mat_B[1][28] +
                  mat_A[12][2] * mat_B[2][28] +
                  mat_A[12][3] * mat_B[3][28] +
                  mat_A[12][4] * mat_B[4][28] +
                  mat_A[12][5] * mat_B[5][28] +
                  mat_A[12][6] * mat_B[6][28] +
                  mat_A[12][7] * mat_B[7][28] +
                  mat_A[12][8] * mat_B[8][28] +
                  mat_A[12][9] * mat_B[9][28] +
                  mat_A[12][10] * mat_B[10][28] +
                  mat_A[12][11] * mat_B[11][28] +
                  mat_A[12][12] * mat_B[12][28] +
                  mat_A[12][13] * mat_B[13][28] +
                  mat_A[12][14] * mat_B[14][28] +
                  mat_A[12][15] * mat_B[15][28] +
                  mat_A[12][16] * mat_B[16][28] +
                  mat_A[12][17] * mat_B[17][28] +
                  mat_A[12][18] * mat_B[18][28] +
                  mat_A[12][19] * mat_B[19][28] +
                  mat_A[12][20] * mat_B[20][28] +
                  mat_A[12][21] * mat_B[21][28] +
                  mat_A[12][22] * mat_B[22][28] +
                  mat_A[12][23] * mat_B[23][28] +
                  mat_A[12][24] * mat_B[24][28] +
                  mat_A[12][25] * mat_B[25][28] +
                  mat_A[12][26] * mat_B[26][28] +
                  mat_A[12][27] * mat_B[27][28] +
                  mat_A[12][28] * mat_B[28][28] +
                  mat_A[12][29] * mat_B[29][28] +
                  mat_A[12][30] * mat_B[30][28] +
                  mat_A[12][31] * mat_B[31][28];
    mat_C[12][29] <= 
                  mat_A[12][0] * mat_B[0][29] +
                  mat_A[12][1] * mat_B[1][29] +
                  mat_A[12][2] * mat_B[2][29] +
                  mat_A[12][3] * mat_B[3][29] +
                  mat_A[12][4] * mat_B[4][29] +
                  mat_A[12][5] * mat_B[5][29] +
                  mat_A[12][6] * mat_B[6][29] +
                  mat_A[12][7] * mat_B[7][29] +
                  mat_A[12][8] * mat_B[8][29] +
                  mat_A[12][9] * mat_B[9][29] +
                  mat_A[12][10] * mat_B[10][29] +
                  mat_A[12][11] * mat_B[11][29] +
                  mat_A[12][12] * mat_B[12][29] +
                  mat_A[12][13] * mat_B[13][29] +
                  mat_A[12][14] * mat_B[14][29] +
                  mat_A[12][15] * mat_B[15][29] +
                  mat_A[12][16] * mat_B[16][29] +
                  mat_A[12][17] * mat_B[17][29] +
                  mat_A[12][18] * mat_B[18][29] +
                  mat_A[12][19] * mat_B[19][29] +
                  mat_A[12][20] * mat_B[20][29] +
                  mat_A[12][21] * mat_B[21][29] +
                  mat_A[12][22] * mat_B[22][29] +
                  mat_A[12][23] * mat_B[23][29] +
                  mat_A[12][24] * mat_B[24][29] +
                  mat_A[12][25] * mat_B[25][29] +
                  mat_A[12][26] * mat_B[26][29] +
                  mat_A[12][27] * mat_B[27][29] +
                  mat_A[12][28] * mat_B[28][29] +
                  mat_A[12][29] * mat_B[29][29] +
                  mat_A[12][30] * mat_B[30][29] +
                  mat_A[12][31] * mat_B[31][29];
    mat_C[12][30] <= 
                  mat_A[12][0] * mat_B[0][30] +
                  mat_A[12][1] * mat_B[1][30] +
                  mat_A[12][2] * mat_B[2][30] +
                  mat_A[12][3] * mat_B[3][30] +
                  mat_A[12][4] * mat_B[4][30] +
                  mat_A[12][5] * mat_B[5][30] +
                  mat_A[12][6] * mat_B[6][30] +
                  mat_A[12][7] * mat_B[7][30] +
                  mat_A[12][8] * mat_B[8][30] +
                  mat_A[12][9] * mat_B[9][30] +
                  mat_A[12][10] * mat_B[10][30] +
                  mat_A[12][11] * mat_B[11][30] +
                  mat_A[12][12] * mat_B[12][30] +
                  mat_A[12][13] * mat_B[13][30] +
                  mat_A[12][14] * mat_B[14][30] +
                  mat_A[12][15] * mat_B[15][30] +
                  mat_A[12][16] * mat_B[16][30] +
                  mat_A[12][17] * mat_B[17][30] +
                  mat_A[12][18] * mat_B[18][30] +
                  mat_A[12][19] * mat_B[19][30] +
                  mat_A[12][20] * mat_B[20][30] +
                  mat_A[12][21] * mat_B[21][30] +
                  mat_A[12][22] * mat_B[22][30] +
                  mat_A[12][23] * mat_B[23][30] +
                  mat_A[12][24] * mat_B[24][30] +
                  mat_A[12][25] * mat_B[25][30] +
                  mat_A[12][26] * mat_B[26][30] +
                  mat_A[12][27] * mat_B[27][30] +
                  mat_A[12][28] * mat_B[28][30] +
                  mat_A[12][29] * mat_B[29][30] +
                  mat_A[12][30] * mat_B[30][30] +
                  mat_A[12][31] * mat_B[31][30];
    mat_C[12][31] <= 
                  mat_A[12][0] * mat_B[0][31] +
                  mat_A[12][1] * mat_B[1][31] +
                  mat_A[12][2] * mat_B[2][31] +
                  mat_A[12][3] * mat_B[3][31] +
                  mat_A[12][4] * mat_B[4][31] +
                  mat_A[12][5] * mat_B[5][31] +
                  mat_A[12][6] * mat_B[6][31] +
                  mat_A[12][7] * mat_B[7][31] +
                  mat_A[12][8] * mat_B[8][31] +
                  mat_A[12][9] * mat_B[9][31] +
                  mat_A[12][10] * mat_B[10][31] +
                  mat_A[12][11] * mat_B[11][31] +
                  mat_A[12][12] * mat_B[12][31] +
                  mat_A[12][13] * mat_B[13][31] +
                  mat_A[12][14] * mat_B[14][31] +
                  mat_A[12][15] * mat_B[15][31] +
                  mat_A[12][16] * mat_B[16][31] +
                  mat_A[12][17] * mat_B[17][31] +
                  mat_A[12][18] * mat_B[18][31] +
                  mat_A[12][19] * mat_B[19][31] +
                  mat_A[12][20] * mat_B[20][31] +
                  mat_A[12][21] * mat_B[21][31] +
                  mat_A[12][22] * mat_B[22][31] +
                  mat_A[12][23] * mat_B[23][31] +
                  mat_A[12][24] * mat_B[24][31] +
                  mat_A[12][25] * mat_B[25][31] +
                  mat_A[12][26] * mat_B[26][31] +
                  mat_A[12][27] * mat_B[27][31] +
                  mat_A[12][28] * mat_B[28][31] +
                  mat_A[12][29] * mat_B[29][31] +
                  mat_A[12][30] * mat_B[30][31] +
                  mat_A[12][31] * mat_B[31][31];
    mat_C[13][0] <= 
                  mat_A[13][0] * mat_B[0][0] +
                  mat_A[13][1] * mat_B[1][0] +
                  mat_A[13][2] * mat_B[2][0] +
                  mat_A[13][3] * mat_B[3][0] +
                  mat_A[13][4] * mat_B[4][0] +
                  mat_A[13][5] * mat_B[5][0] +
                  mat_A[13][6] * mat_B[6][0] +
                  mat_A[13][7] * mat_B[7][0] +
                  mat_A[13][8] * mat_B[8][0] +
                  mat_A[13][9] * mat_B[9][0] +
                  mat_A[13][10] * mat_B[10][0] +
                  mat_A[13][11] * mat_B[11][0] +
                  mat_A[13][12] * mat_B[12][0] +
                  mat_A[13][13] * mat_B[13][0] +
                  mat_A[13][14] * mat_B[14][0] +
                  mat_A[13][15] * mat_B[15][0] +
                  mat_A[13][16] * mat_B[16][0] +
                  mat_A[13][17] * mat_B[17][0] +
                  mat_A[13][18] * mat_B[18][0] +
                  mat_A[13][19] * mat_B[19][0] +
                  mat_A[13][20] * mat_B[20][0] +
                  mat_A[13][21] * mat_B[21][0] +
                  mat_A[13][22] * mat_B[22][0] +
                  mat_A[13][23] * mat_B[23][0] +
                  mat_A[13][24] * mat_B[24][0] +
                  mat_A[13][25] * mat_B[25][0] +
                  mat_A[13][26] * mat_B[26][0] +
                  mat_A[13][27] * mat_B[27][0] +
                  mat_A[13][28] * mat_B[28][0] +
                  mat_A[13][29] * mat_B[29][0] +
                  mat_A[13][30] * mat_B[30][0] +
                  mat_A[13][31] * mat_B[31][0];
    mat_C[13][1] <= 
                  mat_A[13][0] * mat_B[0][1] +
                  mat_A[13][1] * mat_B[1][1] +
                  mat_A[13][2] * mat_B[2][1] +
                  mat_A[13][3] * mat_B[3][1] +
                  mat_A[13][4] * mat_B[4][1] +
                  mat_A[13][5] * mat_B[5][1] +
                  mat_A[13][6] * mat_B[6][1] +
                  mat_A[13][7] * mat_B[7][1] +
                  mat_A[13][8] * mat_B[8][1] +
                  mat_A[13][9] * mat_B[9][1] +
                  mat_A[13][10] * mat_B[10][1] +
                  mat_A[13][11] * mat_B[11][1] +
                  mat_A[13][12] * mat_B[12][1] +
                  mat_A[13][13] * mat_B[13][1] +
                  mat_A[13][14] * mat_B[14][1] +
                  mat_A[13][15] * mat_B[15][1] +
                  mat_A[13][16] * mat_B[16][1] +
                  mat_A[13][17] * mat_B[17][1] +
                  mat_A[13][18] * mat_B[18][1] +
                  mat_A[13][19] * mat_B[19][1] +
                  mat_A[13][20] * mat_B[20][1] +
                  mat_A[13][21] * mat_B[21][1] +
                  mat_A[13][22] * mat_B[22][1] +
                  mat_A[13][23] * mat_B[23][1] +
                  mat_A[13][24] * mat_B[24][1] +
                  mat_A[13][25] * mat_B[25][1] +
                  mat_A[13][26] * mat_B[26][1] +
                  mat_A[13][27] * mat_B[27][1] +
                  mat_A[13][28] * mat_B[28][1] +
                  mat_A[13][29] * mat_B[29][1] +
                  mat_A[13][30] * mat_B[30][1] +
                  mat_A[13][31] * mat_B[31][1];
    mat_C[13][2] <= 
                  mat_A[13][0] * mat_B[0][2] +
                  mat_A[13][1] * mat_B[1][2] +
                  mat_A[13][2] * mat_B[2][2] +
                  mat_A[13][3] * mat_B[3][2] +
                  mat_A[13][4] * mat_B[4][2] +
                  mat_A[13][5] * mat_B[5][2] +
                  mat_A[13][6] * mat_B[6][2] +
                  mat_A[13][7] * mat_B[7][2] +
                  mat_A[13][8] * mat_B[8][2] +
                  mat_A[13][9] * mat_B[9][2] +
                  mat_A[13][10] * mat_B[10][2] +
                  mat_A[13][11] * mat_B[11][2] +
                  mat_A[13][12] * mat_B[12][2] +
                  mat_A[13][13] * mat_B[13][2] +
                  mat_A[13][14] * mat_B[14][2] +
                  mat_A[13][15] * mat_B[15][2] +
                  mat_A[13][16] * mat_B[16][2] +
                  mat_A[13][17] * mat_B[17][2] +
                  mat_A[13][18] * mat_B[18][2] +
                  mat_A[13][19] * mat_B[19][2] +
                  mat_A[13][20] * mat_B[20][2] +
                  mat_A[13][21] * mat_B[21][2] +
                  mat_A[13][22] * mat_B[22][2] +
                  mat_A[13][23] * mat_B[23][2] +
                  mat_A[13][24] * mat_B[24][2] +
                  mat_A[13][25] * mat_B[25][2] +
                  mat_A[13][26] * mat_B[26][2] +
                  mat_A[13][27] * mat_B[27][2] +
                  mat_A[13][28] * mat_B[28][2] +
                  mat_A[13][29] * mat_B[29][2] +
                  mat_A[13][30] * mat_B[30][2] +
                  mat_A[13][31] * mat_B[31][2];
    mat_C[13][3] <= 
                  mat_A[13][0] * mat_B[0][3] +
                  mat_A[13][1] * mat_B[1][3] +
                  mat_A[13][2] * mat_B[2][3] +
                  mat_A[13][3] * mat_B[3][3] +
                  mat_A[13][4] * mat_B[4][3] +
                  mat_A[13][5] * mat_B[5][3] +
                  mat_A[13][6] * mat_B[6][3] +
                  mat_A[13][7] * mat_B[7][3] +
                  mat_A[13][8] * mat_B[8][3] +
                  mat_A[13][9] * mat_B[9][3] +
                  mat_A[13][10] * mat_B[10][3] +
                  mat_A[13][11] * mat_B[11][3] +
                  mat_A[13][12] * mat_B[12][3] +
                  mat_A[13][13] * mat_B[13][3] +
                  mat_A[13][14] * mat_B[14][3] +
                  mat_A[13][15] * mat_B[15][3] +
                  mat_A[13][16] * mat_B[16][3] +
                  mat_A[13][17] * mat_B[17][3] +
                  mat_A[13][18] * mat_B[18][3] +
                  mat_A[13][19] * mat_B[19][3] +
                  mat_A[13][20] * mat_B[20][3] +
                  mat_A[13][21] * mat_B[21][3] +
                  mat_A[13][22] * mat_B[22][3] +
                  mat_A[13][23] * mat_B[23][3] +
                  mat_A[13][24] * mat_B[24][3] +
                  mat_A[13][25] * mat_B[25][3] +
                  mat_A[13][26] * mat_B[26][3] +
                  mat_A[13][27] * mat_B[27][3] +
                  mat_A[13][28] * mat_B[28][3] +
                  mat_A[13][29] * mat_B[29][3] +
                  mat_A[13][30] * mat_B[30][3] +
                  mat_A[13][31] * mat_B[31][3];
    mat_C[13][4] <= 
                  mat_A[13][0] * mat_B[0][4] +
                  mat_A[13][1] * mat_B[1][4] +
                  mat_A[13][2] * mat_B[2][4] +
                  mat_A[13][3] * mat_B[3][4] +
                  mat_A[13][4] * mat_B[4][4] +
                  mat_A[13][5] * mat_B[5][4] +
                  mat_A[13][6] * mat_B[6][4] +
                  mat_A[13][7] * mat_B[7][4] +
                  mat_A[13][8] * mat_B[8][4] +
                  mat_A[13][9] * mat_B[9][4] +
                  mat_A[13][10] * mat_B[10][4] +
                  mat_A[13][11] * mat_B[11][4] +
                  mat_A[13][12] * mat_B[12][4] +
                  mat_A[13][13] * mat_B[13][4] +
                  mat_A[13][14] * mat_B[14][4] +
                  mat_A[13][15] * mat_B[15][4] +
                  mat_A[13][16] * mat_B[16][4] +
                  mat_A[13][17] * mat_B[17][4] +
                  mat_A[13][18] * mat_B[18][4] +
                  mat_A[13][19] * mat_B[19][4] +
                  mat_A[13][20] * mat_B[20][4] +
                  mat_A[13][21] * mat_B[21][4] +
                  mat_A[13][22] * mat_B[22][4] +
                  mat_A[13][23] * mat_B[23][4] +
                  mat_A[13][24] * mat_B[24][4] +
                  mat_A[13][25] * mat_B[25][4] +
                  mat_A[13][26] * mat_B[26][4] +
                  mat_A[13][27] * mat_B[27][4] +
                  mat_A[13][28] * mat_B[28][4] +
                  mat_A[13][29] * mat_B[29][4] +
                  mat_A[13][30] * mat_B[30][4] +
                  mat_A[13][31] * mat_B[31][4];
    mat_C[13][5] <= 
                  mat_A[13][0] * mat_B[0][5] +
                  mat_A[13][1] * mat_B[1][5] +
                  mat_A[13][2] * mat_B[2][5] +
                  mat_A[13][3] * mat_B[3][5] +
                  mat_A[13][4] * mat_B[4][5] +
                  mat_A[13][5] * mat_B[5][5] +
                  mat_A[13][6] * mat_B[6][5] +
                  mat_A[13][7] * mat_B[7][5] +
                  mat_A[13][8] * mat_B[8][5] +
                  mat_A[13][9] * mat_B[9][5] +
                  mat_A[13][10] * mat_B[10][5] +
                  mat_A[13][11] * mat_B[11][5] +
                  mat_A[13][12] * mat_B[12][5] +
                  mat_A[13][13] * mat_B[13][5] +
                  mat_A[13][14] * mat_B[14][5] +
                  mat_A[13][15] * mat_B[15][5] +
                  mat_A[13][16] * mat_B[16][5] +
                  mat_A[13][17] * mat_B[17][5] +
                  mat_A[13][18] * mat_B[18][5] +
                  mat_A[13][19] * mat_B[19][5] +
                  mat_A[13][20] * mat_B[20][5] +
                  mat_A[13][21] * mat_B[21][5] +
                  mat_A[13][22] * mat_B[22][5] +
                  mat_A[13][23] * mat_B[23][5] +
                  mat_A[13][24] * mat_B[24][5] +
                  mat_A[13][25] * mat_B[25][5] +
                  mat_A[13][26] * mat_B[26][5] +
                  mat_A[13][27] * mat_B[27][5] +
                  mat_A[13][28] * mat_B[28][5] +
                  mat_A[13][29] * mat_B[29][5] +
                  mat_A[13][30] * mat_B[30][5] +
                  mat_A[13][31] * mat_B[31][5];
    mat_C[13][6] <= 
                  mat_A[13][0] * mat_B[0][6] +
                  mat_A[13][1] * mat_B[1][6] +
                  mat_A[13][2] * mat_B[2][6] +
                  mat_A[13][3] * mat_B[3][6] +
                  mat_A[13][4] * mat_B[4][6] +
                  mat_A[13][5] * mat_B[5][6] +
                  mat_A[13][6] * mat_B[6][6] +
                  mat_A[13][7] * mat_B[7][6] +
                  mat_A[13][8] * mat_B[8][6] +
                  mat_A[13][9] * mat_B[9][6] +
                  mat_A[13][10] * mat_B[10][6] +
                  mat_A[13][11] * mat_B[11][6] +
                  mat_A[13][12] * mat_B[12][6] +
                  mat_A[13][13] * mat_B[13][6] +
                  mat_A[13][14] * mat_B[14][6] +
                  mat_A[13][15] * mat_B[15][6] +
                  mat_A[13][16] * mat_B[16][6] +
                  mat_A[13][17] * mat_B[17][6] +
                  mat_A[13][18] * mat_B[18][6] +
                  mat_A[13][19] * mat_B[19][6] +
                  mat_A[13][20] * mat_B[20][6] +
                  mat_A[13][21] * mat_B[21][6] +
                  mat_A[13][22] * mat_B[22][6] +
                  mat_A[13][23] * mat_B[23][6] +
                  mat_A[13][24] * mat_B[24][6] +
                  mat_A[13][25] * mat_B[25][6] +
                  mat_A[13][26] * mat_B[26][6] +
                  mat_A[13][27] * mat_B[27][6] +
                  mat_A[13][28] * mat_B[28][6] +
                  mat_A[13][29] * mat_B[29][6] +
                  mat_A[13][30] * mat_B[30][6] +
                  mat_A[13][31] * mat_B[31][6];
    mat_C[13][7] <= 
                  mat_A[13][0] * mat_B[0][7] +
                  mat_A[13][1] * mat_B[1][7] +
                  mat_A[13][2] * mat_B[2][7] +
                  mat_A[13][3] * mat_B[3][7] +
                  mat_A[13][4] * mat_B[4][7] +
                  mat_A[13][5] * mat_B[5][7] +
                  mat_A[13][6] * mat_B[6][7] +
                  mat_A[13][7] * mat_B[7][7] +
                  mat_A[13][8] * mat_B[8][7] +
                  mat_A[13][9] * mat_B[9][7] +
                  mat_A[13][10] * mat_B[10][7] +
                  mat_A[13][11] * mat_B[11][7] +
                  mat_A[13][12] * mat_B[12][7] +
                  mat_A[13][13] * mat_B[13][7] +
                  mat_A[13][14] * mat_B[14][7] +
                  mat_A[13][15] * mat_B[15][7] +
                  mat_A[13][16] * mat_B[16][7] +
                  mat_A[13][17] * mat_B[17][7] +
                  mat_A[13][18] * mat_B[18][7] +
                  mat_A[13][19] * mat_B[19][7] +
                  mat_A[13][20] * mat_B[20][7] +
                  mat_A[13][21] * mat_B[21][7] +
                  mat_A[13][22] * mat_B[22][7] +
                  mat_A[13][23] * mat_B[23][7] +
                  mat_A[13][24] * mat_B[24][7] +
                  mat_A[13][25] * mat_B[25][7] +
                  mat_A[13][26] * mat_B[26][7] +
                  mat_A[13][27] * mat_B[27][7] +
                  mat_A[13][28] * mat_B[28][7] +
                  mat_A[13][29] * mat_B[29][7] +
                  mat_A[13][30] * mat_B[30][7] +
                  mat_A[13][31] * mat_B[31][7];
    mat_C[13][8] <= 
                  mat_A[13][0] * mat_B[0][8] +
                  mat_A[13][1] * mat_B[1][8] +
                  mat_A[13][2] * mat_B[2][8] +
                  mat_A[13][3] * mat_B[3][8] +
                  mat_A[13][4] * mat_B[4][8] +
                  mat_A[13][5] * mat_B[5][8] +
                  mat_A[13][6] * mat_B[6][8] +
                  mat_A[13][7] * mat_B[7][8] +
                  mat_A[13][8] * mat_B[8][8] +
                  mat_A[13][9] * mat_B[9][8] +
                  mat_A[13][10] * mat_B[10][8] +
                  mat_A[13][11] * mat_B[11][8] +
                  mat_A[13][12] * mat_B[12][8] +
                  mat_A[13][13] * mat_B[13][8] +
                  mat_A[13][14] * mat_B[14][8] +
                  mat_A[13][15] * mat_B[15][8] +
                  mat_A[13][16] * mat_B[16][8] +
                  mat_A[13][17] * mat_B[17][8] +
                  mat_A[13][18] * mat_B[18][8] +
                  mat_A[13][19] * mat_B[19][8] +
                  mat_A[13][20] * mat_B[20][8] +
                  mat_A[13][21] * mat_B[21][8] +
                  mat_A[13][22] * mat_B[22][8] +
                  mat_A[13][23] * mat_B[23][8] +
                  mat_A[13][24] * mat_B[24][8] +
                  mat_A[13][25] * mat_B[25][8] +
                  mat_A[13][26] * mat_B[26][8] +
                  mat_A[13][27] * mat_B[27][8] +
                  mat_A[13][28] * mat_B[28][8] +
                  mat_A[13][29] * mat_B[29][8] +
                  mat_A[13][30] * mat_B[30][8] +
                  mat_A[13][31] * mat_B[31][8];
    mat_C[13][9] <= 
                  mat_A[13][0] * mat_B[0][9] +
                  mat_A[13][1] * mat_B[1][9] +
                  mat_A[13][2] * mat_B[2][9] +
                  mat_A[13][3] * mat_B[3][9] +
                  mat_A[13][4] * mat_B[4][9] +
                  mat_A[13][5] * mat_B[5][9] +
                  mat_A[13][6] * mat_B[6][9] +
                  mat_A[13][7] * mat_B[7][9] +
                  mat_A[13][8] * mat_B[8][9] +
                  mat_A[13][9] * mat_B[9][9] +
                  mat_A[13][10] * mat_B[10][9] +
                  mat_A[13][11] * mat_B[11][9] +
                  mat_A[13][12] * mat_B[12][9] +
                  mat_A[13][13] * mat_B[13][9] +
                  mat_A[13][14] * mat_B[14][9] +
                  mat_A[13][15] * mat_B[15][9] +
                  mat_A[13][16] * mat_B[16][9] +
                  mat_A[13][17] * mat_B[17][9] +
                  mat_A[13][18] * mat_B[18][9] +
                  mat_A[13][19] * mat_B[19][9] +
                  mat_A[13][20] * mat_B[20][9] +
                  mat_A[13][21] * mat_B[21][9] +
                  mat_A[13][22] * mat_B[22][9] +
                  mat_A[13][23] * mat_B[23][9] +
                  mat_A[13][24] * mat_B[24][9] +
                  mat_A[13][25] * mat_B[25][9] +
                  mat_A[13][26] * mat_B[26][9] +
                  mat_A[13][27] * mat_B[27][9] +
                  mat_A[13][28] * mat_B[28][9] +
                  mat_A[13][29] * mat_B[29][9] +
                  mat_A[13][30] * mat_B[30][9] +
                  mat_A[13][31] * mat_B[31][9];
    mat_C[13][10] <= 
                  mat_A[13][0] * mat_B[0][10] +
                  mat_A[13][1] * mat_B[1][10] +
                  mat_A[13][2] * mat_B[2][10] +
                  mat_A[13][3] * mat_B[3][10] +
                  mat_A[13][4] * mat_B[4][10] +
                  mat_A[13][5] * mat_B[5][10] +
                  mat_A[13][6] * mat_B[6][10] +
                  mat_A[13][7] * mat_B[7][10] +
                  mat_A[13][8] * mat_B[8][10] +
                  mat_A[13][9] * mat_B[9][10] +
                  mat_A[13][10] * mat_B[10][10] +
                  mat_A[13][11] * mat_B[11][10] +
                  mat_A[13][12] * mat_B[12][10] +
                  mat_A[13][13] * mat_B[13][10] +
                  mat_A[13][14] * mat_B[14][10] +
                  mat_A[13][15] * mat_B[15][10] +
                  mat_A[13][16] * mat_B[16][10] +
                  mat_A[13][17] * mat_B[17][10] +
                  mat_A[13][18] * mat_B[18][10] +
                  mat_A[13][19] * mat_B[19][10] +
                  mat_A[13][20] * mat_B[20][10] +
                  mat_A[13][21] * mat_B[21][10] +
                  mat_A[13][22] * mat_B[22][10] +
                  mat_A[13][23] * mat_B[23][10] +
                  mat_A[13][24] * mat_B[24][10] +
                  mat_A[13][25] * mat_B[25][10] +
                  mat_A[13][26] * mat_B[26][10] +
                  mat_A[13][27] * mat_B[27][10] +
                  mat_A[13][28] * mat_B[28][10] +
                  mat_A[13][29] * mat_B[29][10] +
                  mat_A[13][30] * mat_B[30][10] +
                  mat_A[13][31] * mat_B[31][10];
    mat_C[13][11] <= 
                  mat_A[13][0] * mat_B[0][11] +
                  mat_A[13][1] * mat_B[1][11] +
                  mat_A[13][2] * mat_B[2][11] +
                  mat_A[13][3] * mat_B[3][11] +
                  mat_A[13][4] * mat_B[4][11] +
                  mat_A[13][5] * mat_B[5][11] +
                  mat_A[13][6] * mat_B[6][11] +
                  mat_A[13][7] * mat_B[7][11] +
                  mat_A[13][8] * mat_B[8][11] +
                  mat_A[13][9] * mat_B[9][11] +
                  mat_A[13][10] * mat_B[10][11] +
                  mat_A[13][11] * mat_B[11][11] +
                  mat_A[13][12] * mat_B[12][11] +
                  mat_A[13][13] * mat_B[13][11] +
                  mat_A[13][14] * mat_B[14][11] +
                  mat_A[13][15] * mat_B[15][11] +
                  mat_A[13][16] * mat_B[16][11] +
                  mat_A[13][17] * mat_B[17][11] +
                  mat_A[13][18] * mat_B[18][11] +
                  mat_A[13][19] * mat_B[19][11] +
                  mat_A[13][20] * mat_B[20][11] +
                  mat_A[13][21] * mat_B[21][11] +
                  mat_A[13][22] * mat_B[22][11] +
                  mat_A[13][23] * mat_B[23][11] +
                  mat_A[13][24] * mat_B[24][11] +
                  mat_A[13][25] * mat_B[25][11] +
                  mat_A[13][26] * mat_B[26][11] +
                  mat_A[13][27] * mat_B[27][11] +
                  mat_A[13][28] * mat_B[28][11] +
                  mat_A[13][29] * mat_B[29][11] +
                  mat_A[13][30] * mat_B[30][11] +
                  mat_A[13][31] * mat_B[31][11];
    mat_C[13][12] <= 
                  mat_A[13][0] * mat_B[0][12] +
                  mat_A[13][1] * mat_B[1][12] +
                  mat_A[13][2] * mat_B[2][12] +
                  mat_A[13][3] * mat_B[3][12] +
                  mat_A[13][4] * mat_B[4][12] +
                  mat_A[13][5] * mat_B[5][12] +
                  mat_A[13][6] * mat_B[6][12] +
                  mat_A[13][7] * mat_B[7][12] +
                  mat_A[13][8] * mat_B[8][12] +
                  mat_A[13][9] * mat_B[9][12] +
                  mat_A[13][10] * mat_B[10][12] +
                  mat_A[13][11] * mat_B[11][12] +
                  mat_A[13][12] * mat_B[12][12] +
                  mat_A[13][13] * mat_B[13][12] +
                  mat_A[13][14] * mat_B[14][12] +
                  mat_A[13][15] * mat_B[15][12] +
                  mat_A[13][16] * mat_B[16][12] +
                  mat_A[13][17] * mat_B[17][12] +
                  mat_A[13][18] * mat_B[18][12] +
                  mat_A[13][19] * mat_B[19][12] +
                  mat_A[13][20] * mat_B[20][12] +
                  mat_A[13][21] * mat_B[21][12] +
                  mat_A[13][22] * mat_B[22][12] +
                  mat_A[13][23] * mat_B[23][12] +
                  mat_A[13][24] * mat_B[24][12] +
                  mat_A[13][25] * mat_B[25][12] +
                  mat_A[13][26] * mat_B[26][12] +
                  mat_A[13][27] * mat_B[27][12] +
                  mat_A[13][28] * mat_B[28][12] +
                  mat_A[13][29] * mat_B[29][12] +
                  mat_A[13][30] * mat_B[30][12] +
                  mat_A[13][31] * mat_B[31][12];
    mat_C[13][13] <= 
                  mat_A[13][0] * mat_B[0][13] +
                  mat_A[13][1] * mat_B[1][13] +
                  mat_A[13][2] * mat_B[2][13] +
                  mat_A[13][3] * mat_B[3][13] +
                  mat_A[13][4] * mat_B[4][13] +
                  mat_A[13][5] * mat_B[5][13] +
                  mat_A[13][6] * mat_B[6][13] +
                  mat_A[13][7] * mat_B[7][13] +
                  mat_A[13][8] * mat_B[8][13] +
                  mat_A[13][9] * mat_B[9][13] +
                  mat_A[13][10] * mat_B[10][13] +
                  mat_A[13][11] * mat_B[11][13] +
                  mat_A[13][12] * mat_B[12][13] +
                  mat_A[13][13] * mat_B[13][13] +
                  mat_A[13][14] * mat_B[14][13] +
                  mat_A[13][15] * mat_B[15][13] +
                  mat_A[13][16] * mat_B[16][13] +
                  mat_A[13][17] * mat_B[17][13] +
                  mat_A[13][18] * mat_B[18][13] +
                  mat_A[13][19] * mat_B[19][13] +
                  mat_A[13][20] * mat_B[20][13] +
                  mat_A[13][21] * mat_B[21][13] +
                  mat_A[13][22] * mat_B[22][13] +
                  mat_A[13][23] * mat_B[23][13] +
                  mat_A[13][24] * mat_B[24][13] +
                  mat_A[13][25] * mat_B[25][13] +
                  mat_A[13][26] * mat_B[26][13] +
                  mat_A[13][27] * mat_B[27][13] +
                  mat_A[13][28] * mat_B[28][13] +
                  mat_A[13][29] * mat_B[29][13] +
                  mat_A[13][30] * mat_B[30][13] +
                  mat_A[13][31] * mat_B[31][13];
    mat_C[13][14] <= 
                  mat_A[13][0] * mat_B[0][14] +
                  mat_A[13][1] * mat_B[1][14] +
                  mat_A[13][2] * mat_B[2][14] +
                  mat_A[13][3] * mat_B[3][14] +
                  mat_A[13][4] * mat_B[4][14] +
                  mat_A[13][5] * mat_B[5][14] +
                  mat_A[13][6] * mat_B[6][14] +
                  mat_A[13][7] * mat_B[7][14] +
                  mat_A[13][8] * mat_B[8][14] +
                  mat_A[13][9] * mat_B[9][14] +
                  mat_A[13][10] * mat_B[10][14] +
                  mat_A[13][11] * mat_B[11][14] +
                  mat_A[13][12] * mat_B[12][14] +
                  mat_A[13][13] * mat_B[13][14] +
                  mat_A[13][14] * mat_B[14][14] +
                  mat_A[13][15] * mat_B[15][14] +
                  mat_A[13][16] * mat_B[16][14] +
                  mat_A[13][17] * mat_B[17][14] +
                  mat_A[13][18] * mat_B[18][14] +
                  mat_A[13][19] * mat_B[19][14] +
                  mat_A[13][20] * mat_B[20][14] +
                  mat_A[13][21] * mat_B[21][14] +
                  mat_A[13][22] * mat_B[22][14] +
                  mat_A[13][23] * mat_B[23][14] +
                  mat_A[13][24] * mat_B[24][14] +
                  mat_A[13][25] * mat_B[25][14] +
                  mat_A[13][26] * mat_B[26][14] +
                  mat_A[13][27] * mat_B[27][14] +
                  mat_A[13][28] * mat_B[28][14] +
                  mat_A[13][29] * mat_B[29][14] +
                  mat_A[13][30] * mat_B[30][14] +
                  mat_A[13][31] * mat_B[31][14];
    mat_C[13][15] <= 
                  mat_A[13][0] * mat_B[0][15] +
                  mat_A[13][1] * mat_B[1][15] +
                  mat_A[13][2] * mat_B[2][15] +
                  mat_A[13][3] * mat_B[3][15] +
                  mat_A[13][4] * mat_B[4][15] +
                  mat_A[13][5] * mat_B[5][15] +
                  mat_A[13][6] * mat_B[6][15] +
                  mat_A[13][7] * mat_B[7][15] +
                  mat_A[13][8] * mat_B[8][15] +
                  mat_A[13][9] * mat_B[9][15] +
                  mat_A[13][10] * mat_B[10][15] +
                  mat_A[13][11] * mat_B[11][15] +
                  mat_A[13][12] * mat_B[12][15] +
                  mat_A[13][13] * mat_B[13][15] +
                  mat_A[13][14] * mat_B[14][15] +
                  mat_A[13][15] * mat_B[15][15] +
                  mat_A[13][16] * mat_B[16][15] +
                  mat_A[13][17] * mat_B[17][15] +
                  mat_A[13][18] * mat_B[18][15] +
                  mat_A[13][19] * mat_B[19][15] +
                  mat_A[13][20] * mat_B[20][15] +
                  mat_A[13][21] * mat_B[21][15] +
                  mat_A[13][22] * mat_B[22][15] +
                  mat_A[13][23] * mat_B[23][15] +
                  mat_A[13][24] * mat_B[24][15] +
                  mat_A[13][25] * mat_B[25][15] +
                  mat_A[13][26] * mat_B[26][15] +
                  mat_A[13][27] * mat_B[27][15] +
                  mat_A[13][28] * mat_B[28][15] +
                  mat_A[13][29] * mat_B[29][15] +
                  mat_A[13][30] * mat_B[30][15] +
                  mat_A[13][31] * mat_B[31][15];
    mat_C[13][16] <= 
                  mat_A[13][0] * mat_B[0][16] +
                  mat_A[13][1] * mat_B[1][16] +
                  mat_A[13][2] * mat_B[2][16] +
                  mat_A[13][3] * mat_B[3][16] +
                  mat_A[13][4] * mat_B[4][16] +
                  mat_A[13][5] * mat_B[5][16] +
                  mat_A[13][6] * mat_B[6][16] +
                  mat_A[13][7] * mat_B[7][16] +
                  mat_A[13][8] * mat_B[8][16] +
                  mat_A[13][9] * mat_B[9][16] +
                  mat_A[13][10] * mat_B[10][16] +
                  mat_A[13][11] * mat_B[11][16] +
                  mat_A[13][12] * mat_B[12][16] +
                  mat_A[13][13] * mat_B[13][16] +
                  mat_A[13][14] * mat_B[14][16] +
                  mat_A[13][15] * mat_B[15][16] +
                  mat_A[13][16] * mat_B[16][16] +
                  mat_A[13][17] * mat_B[17][16] +
                  mat_A[13][18] * mat_B[18][16] +
                  mat_A[13][19] * mat_B[19][16] +
                  mat_A[13][20] * mat_B[20][16] +
                  mat_A[13][21] * mat_B[21][16] +
                  mat_A[13][22] * mat_B[22][16] +
                  mat_A[13][23] * mat_B[23][16] +
                  mat_A[13][24] * mat_B[24][16] +
                  mat_A[13][25] * mat_B[25][16] +
                  mat_A[13][26] * mat_B[26][16] +
                  mat_A[13][27] * mat_B[27][16] +
                  mat_A[13][28] * mat_B[28][16] +
                  mat_A[13][29] * mat_B[29][16] +
                  mat_A[13][30] * mat_B[30][16] +
                  mat_A[13][31] * mat_B[31][16];
    mat_C[13][17] <= 
                  mat_A[13][0] * mat_B[0][17] +
                  mat_A[13][1] * mat_B[1][17] +
                  mat_A[13][2] * mat_B[2][17] +
                  mat_A[13][3] * mat_B[3][17] +
                  mat_A[13][4] * mat_B[4][17] +
                  mat_A[13][5] * mat_B[5][17] +
                  mat_A[13][6] * mat_B[6][17] +
                  mat_A[13][7] * mat_B[7][17] +
                  mat_A[13][8] * mat_B[8][17] +
                  mat_A[13][9] * mat_B[9][17] +
                  mat_A[13][10] * mat_B[10][17] +
                  mat_A[13][11] * mat_B[11][17] +
                  mat_A[13][12] * mat_B[12][17] +
                  mat_A[13][13] * mat_B[13][17] +
                  mat_A[13][14] * mat_B[14][17] +
                  mat_A[13][15] * mat_B[15][17] +
                  mat_A[13][16] * mat_B[16][17] +
                  mat_A[13][17] * mat_B[17][17] +
                  mat_A[13][18] * mat_B[18][17] +
                  mat_A[13][19] * mat_B[19][17] +
                  mat_A[13][20] * mat_B[20][17] +
                  mat_A[13][21] * mat_B[21][17] +
                  mat_A[13][22] * mat_B[22][17] +
                  mat_A[13][23] * mat_B[23][17] +
                  mat_A[13][24] * mat_B[24][17] +
                  mat_A[13][25] * mat_B[25][17] +
                  mat_A[13][26] * mat_B[26][17] +
                  mat_A[13][27] * mat_B[27][17] +
                  mat_A[13][28] * mat_B[28][17] +
                  mat_A[13][29] * mat_B[29][17] +
                  mat_A[13][30] * mat_B[30][17] +
                  mat_A[13][31] * mat_B[31][17];
    mat_C[13][18] <= 
                  mat_A[13][0] * mat_B[0][18] +
                  mat_A[13][1] * mat_B[1][18] +
                  mat_A[13][2] * mat_B[2][18] +
                  mat_A[13][3] * mat_B[3][18] +
                  mat_A[13][4] * mat_B[4][18] +
                  mat_A[13][5] * mat_B[5][18] +
                  mat_A[13][6] * mat_B[6][18] +
                  mat_A[13][7] * mat_B[7][18] +
                  mat_A[13][8] * mat_B[8][18] +
                  mat_A[13][9] * mat_B[9][18] +
                  mat_A[13][10] * mat_B[10][18] +
                  mat_A[13][11] * mat_B[11][18] +
                  mat_A[13][12] * mat_B[12][18] +
                  mat_A[13][13] * mat_B[13][18] +
                  mat_A[13][14] * mat_B[14][18] +
                  mat_A[13][15] * mat_B[15][18] +
                  mat_A[13][16] * mat_B[16][18] +
                  mat_A[13][17] * mat_B[17][18] +
                  mat_A[13][18] * mat_B[18][18] +
                  mat_A[13][19] * mat_B[19][18] +
                  mat_A[13][20] * mat_B[20][18] +
                  mat_A[13][21] * mat_B[21][18] +
                  mat_A[13][22] * mat_B[22][18] +
                  mat_A[13][23] * mat_B[23][18] +
                  mat_A[13][24] * mat_B[24][18] +
                  mat_A[13][25] * mat_B[25][18] +
                  mat_A[13][26] * mat_B[26][18] +
                  mat_A[13][27] * mat_B[27][18] +
                  mat_A[13][28] * mat_B[28][18] +
                  mat_A[13][29] * mat_B[29][18] +
                  mat_A[13][30] * mat_B[30][18] +
                  mat_A[13][31] * mat_B[31][18];
    mat_C[13][19] <= 
                  mat_A[13][0] * mat_B[0][19] +
                  mat_A[13][1] * mat_B[1][19] +
                  mat_A[13][2] * mat_B[2][19] +
                  mat_A[13][3] * mat_B[3][19] +
                  mat_A[13][4] * mat_B[4][19] +
                  mat_A[13][5] * mat_B[5][19] +
                  mat_A[13][6] * mat_B[6][19] +
                  mat_A[13][7] * mat_B[7][19] +
                  mat_A[13][8] * mat_B[8][19] +
                  mat_A[13][9] * mat_B[9][19] +
                  mat_A[13][10] * mat_B[10][19] +
                  mat_A[13][11] * mat_B[11][19] +
                  mat_A[13][12] * mat_B[12][19] +
                  mat_A[13][13] * mat_B[13][19] +
                  mat_A[13][14] * mat_B[14][19] +
                  mat_A[13][15] * mat_B[15][19] +
                  mat_A[13][16] * mat_B[16][19] +
                  mat_A[13][17] * mat_B[17][19] +
                  mat_A[13][18] * mat_B[18][19] +
                  mat_A[13][19] * mat_B[19][19] +
                  mat_A[13][20] * mat_B[20][19] +
                  mat_A[13][21] * mat_B[21][19] +
                  mat_A[13][22] * mat_B[22][19] +
                  mat_A[13][23] * mat_B[23][19] +
                  mat_A[13][24] * mat_B[24][19] +
                  mat_A[13][25] * mat_B[25][19] +
                  mat_A[13][26] * mat_B[26][19] +
                  mat_A[13][27] * mat_B[27][19] +
                  mat_A[13][28] * mat_B[28][19] +
                  mat_A[13][29] * mat_B[29][19] +
                  mat_A[13][30] * mat_B[30][19] +
                  mat_A[13][31] * mat_B[31][19];
    mat_C[13][20] <= 
                  mat_A[13][0] * mat_B[0][20] +
                  mat_A[13][1] * mat_B[1][20] +
                  mat_A[13][2] * mat_B[2][20] +
                  mat_A[13][3] * mat_B[3][20] +
                  mat_A[13][4] * mat_B[4][20] +
                  mat_A[13][5] * mat_B[5][20] +
                  mat_A[13][6] * mat_B[6][20] +
                  mat_A[13][7] * mat_B[7][20] +
                  mat_A[13][8] * mat_B[8][20] +
                  mat_A[13][9] * mat_B[9][20] +
                  mat_A[13][10] * mat_B[10][20] +
                  mat_A[13][11] * mat_B[11][20] +
                  mat_A[13][12] * mat_B[12][20] +
                  mat_A[13][13] * mat_B[13][20] +
                  mat_A[13][14] * mat_B[14][20] +
                  mat_A[13][15] * mat_B[15][20] +
                  mat_A[13][16] * mat_B[16][20] +
                  mat_A[13][17] * mat_B[17][20] +
                  mat_A[13][18] * mat_B[18][20] +
                  mat_A[13][19] * mat_B[19][20] +
                  mat_A[13][20] * mat_B[20][20] +
                  mat_A[13][21] * mat_B[21][20] +
                  mat_A[13][22] * mat_B[22][20] +
                  mat_A[13][23] * mat_B[23][20] +
                  mat_A[13][24] * mat_B[24][20] +
                  mat_A[13][25] * mat_B[25][20] +
                  mat_A[13][26] * mat_B[26][20] +
                  mat_A[13][27] * mat_B[27][20] +
                  mat_A[13][28] * mat_B[28][20] +
                  mat_A[13][29] * mat_B[29][20] +
                  mat_A[13][30] * mat_B[30][20] +
                  mat_A[13][31] * mat_B[31][20];
    mat_C[13][21] <= 
                  mat_A[13][0] * mat_B[0][21] +
                  mat_A[13][1] * mat_B[1][21] +
                  mat_A[13][2] * mat_B[2][21] +
                  mat_A[13][3] * mat_B[3][21] +
                  mat_A[13][4] * mat_B[4][21] +
                  mat_A[13][5] * mat_B[5][21] +
                  mat_A[13][6] * mat_B[6][21] +
                  mat_A[13][7] * mat_B[7][21] +
                  mat_A[13][8] * mat_B[8][21] +
                  mat_A[13][9] * mat_B[9][21] +
                  mat_A[13][10] * mat_B[10][21] +
                  mat_A[13][11] * mat_B[11][21] +
                  mat_A[13][12] * mat_B[12][21] +
                  mat_A[13][13] * mat_B[13][21] +
                  mat_A[13][14] * mat_B[14][21] +
                  mat_A[13][15] * mat_B[15][21] +
                  mat_A[13][16] * mat_B[16][21] +
                  mat_A[13][17] * mat_B[17][21] +
                  mat_A[13][18] * mat_B[18][21] +
                  mat_A[13][19] * mat_B[19][21] +
                  mat_A[13][20] * mat_B[20][21] +
                  mat_A[13][21] * mat_B[21][21] +
                  mat_A[13][22] * mat_B[22][21] +
                  mat_A[13][23] * mat_B[23][21] +
                  mat_A[13][24] * mat_B[24][21] +
                  mat_A[13][25] * mat_B[25][21] +
                  mat_A[13][26] * mat_B[26][21] +
                  mat_A[13][27] * mat_B[27][21] +
                  mat_A[13][28] * mat_B[28][21] +
                  mat_A[13][29] * mat_B[29][21] +
                  mat_A[13][30] * mat_B[30][21] +
                  mat_A[13][31] * mat_B[31][21];
    mat_C[13][22] <= 
                  mat_A[13][0] * mat_B[0][22] +
                  mat_A[13][1] * mat_B[1][22] +
                  mat_A[13][2] * mat_B[2][22] +
                  mat_A[13][3] * mat_B[3][22] +
                  mat_A[13][4] * mat_B[4][22] +
                  mat_A[13][5] * mat_B[5][22] +
                  mat_A[13][6] * mat_B[6][22] +
                  mat_A[13][7] * mat_B[7][22] +
                  mat_A[13][8] * mat_B[8][22] +
                  mat_A[13][9] * mat_B[9][22] +
                  mat_A[13][10] * mat_B[10][22] +
                  mat_A[13][11] * mat_B[11][22] +
                  mat_A[13][12] * mat_B[12][22] +
                  mat_A[13][13] * mat_B[13][22] +
                  mat_A[13][14] * mat_B[14][22] +
                  mat_A[13][15] * mat_B[15][22] +
                  mat_A[13][16] * mat_B[16][22] +
                  mat_A[13][17] * mat_B[17][22] +
                  mat_A[13][18] * mat_B[18][22] +
                  mat_A[13][19] * mat_B[19][22] +
                  mat_A[13][20] * mat_B[20][22] +
                  mat_A[13][21] * mat_B[21][22] +
                  mat_A[13][22] * mat_B[22][22] +
                  mat_A[13][23] * mat_B[23][22] +
                  mat_A[13][24] * mat_B[24][22] +
                  mat_A[13][25] * mat_B[25][22] +
                  mat_A[13][26] * mat_B[26][22] +
                  mat_A[13][27] * mat_B[27][22] +
                  mat_A[13][28] * mat_B[28][22] +
                  mat_A[13][29] * mat_B[29][22] +
                  mat_A[13][30] * mat_B[30][22] +
                  mat_A[13][31] * mat_B[31][22];
    mat_C[13][23] <= 
                  mat_A[13][0] * mat_B[0][23] +
                  mat_A[13][1] * mat_B[1][23] +
                  mat_A[13][2] * mat_B[2][23] +
                  mat_A[13][3] * mat_B[3][23] +
                  mat_A[13][4] * mat_B[4][23] +
                  mat_A[13][5] * mat_B[5][23] +
                  mat_A[13][6] * mat_B[6][23] +
                  mat_A[13][7] * mat_B[7][23] +
                  mat_A[13][8] * mat_B[8][23] +
                  mat_A[13][9] * mat_B[9][23] +
                  mat_A[13][10] * mat_B[10][23] +
                  mat_A[13][11] * mat_B[11][23] +
                  mat_A[13][12] * mat_B[12][23] +
                  mat_A[13][13] * mat_B[13][23] +
                  mat_A[13][14] * mat_B[14][23] +
                  mat_A[13][15] * mat_B[15][23] +
                  mat_A[13][16] * mat_B[16][23] +
                  mat_A[13][17] * mat_B[17][23] +
                  mat_A[13][18] * mat_B[18][23] +
                  mat_A[13][19] * mat_B[19][23] +
                  mat_A[13][20] * mat_B[20][23] +
                  mat_A[13][21] * mat_B[21][23] +
                  mat_A[13][22] * mat_B[22][23] +
                  mat_A[13][23] * mat_B[23][23] +
                  mat_A[13][24] * mat_B[24][23] +
                  mat_A[13][25] * mat_B[25][23] +
                  mat_A[13][26] * mat_B[26][23] +
                  mat_A[13][27] * mat_B[27][23] +
                  mat_A[13][28] * mat_B[28][23] +
                  mat_A[13][29] * mat_B[29][23] +
                  mat_A[13][30] * mat_B[30][23] +
                  mat_A[13][31] * mat_B[31][23];
    mat_C[13][24] <= 
                  mat_A[13][0] * mat_B[0][24] +
                  mat_A[13][1] * mat_B[1][24] +
                  mat_A[13][2] * mat_B[2][24] +
                  mat_A[13][3] * mat_B[3][24] +
                  mat_A[13][4] * mat_B[4][24] +
                  mat_A[13][5] * mat_B[5][24] +
                  mat_A[13][6] * mat_B[6][24] +
                  mat_A[13][7] * mat_B[7][24] +
                  mat_A[13][8] * mat_B[8][24] +
                  mat_A[13][9] * mat_B[9][24] +
                  mat_A[13][10] * mat_B[10][24] +
                  mat_A[13][11] * mat_B[11][24] +
                  mat_A[13][12] * mat_B[12][24] +
                  mat_A[13][13] * mat_B[13][24] +
                  mat_A[13][14] * mat_B[14][24] +
                  mat_A[13][15] * mat_B[15][24] +
                  mat_A[13][16] * mat_B[16][24] +
                  mat_A[13][17] * mat_B[17][24] +
                  mat_A[13][18] * mat_B[18][24] +
                  mat_A[13][19] * mat_B[19][24] +
                  mat_A[13][20] * mat_B[20][24] +
                  mat_A[13][21] * mat_B[21][24] +
                  mat_A[13][22] * mat_B[22][24] +
                  mat_A[13][23] * mat_B[23][24] +
                  mat_A[13][24] * mat_B[24][24] +
                  mat_A[13][25] * mat_B[25][24] +
                  mat_A[13][26] * mat_B[26][24] +
                  mat_A[13][27] * mat_B[27][24] +
                  mat_A[13][28] * mat_B[28][24] +
                  mat_A[13][29] * mat_B[29][24] +
                  mat_A[13][30] * mat_B[30][24] +
                  mat_A[13][31] * mat_B[31][24];
    mat_C[13][25] <= 
                  mat_A[13][0] * mat_B[0][25] +
                  mat_A[13][1] * mat_B[1][25] +
                  mat_A[13][2] * mat_B[2][25] +
                  mat_A[13][3] * mat_B[3][25] +
                  mat_A[13][4] * mat_B[4][25] +
                  mat_A[13][5] * mat_B[5][25] +
                  mat_A[13][6] * mat_B[6][25] +
                  mat_A[13][7] * mat_B[7][25] +
                  mat_A[13][8] * mat_B[8][25] +
                  mat_A[13][9] * mat_B[9][25] +
                  mat_A[13][10] * mat_B[10][25] +
                  mat_A[13][11] * mat_B[11][25] +
                  mat_A[13][12] * mat_B[12][25] +
                  mat_A[13][13] * mat_B[13][25] +
                  mat_A[13][14] * mat_B[14][25] +
                  mat_A[13][15] * mat_B[15][25] +
                  mat_A[13][16] * mat_B[16][25] +
                  mat_A[13][17] * mat_B[17][25] +
                  mat_A[13][18] * mat_B[18][25] +
                  mat_A[13][19] * mat_B[19][25] +
                  mat_A[13][20] * mat_B[20][25] +
                  mat_A[13][21] * mat_B[21][25] +
                  mat_A[13][22] * mat_B[22][25] +
                  mat_A[13][23] * mat_B[23][25] +
                  mat_A[13][24] * mat_B[24][25] +
                  mat_A[13][25] * mat_B[25][25] +
                  mat_A[13][26] * mat_B[26][25] +
                  mat_A[13][27] * mat_B[27][25] +
                  mat_A[13][28] * mat_B[28][25] +
                  mat_A[13][29] * mat_B[29][25] +
                  mat_A[13][30] * mat_B[30][25] +
                  mat_A[13][31] * mat_B[31][25];
    mat_C[13][26] <= 
                  mat_A[13][0] * mat_B[0][26] +
                  mat_A[13][1] * mat_B[1][26] +
                  mat_A[13][2] * mat_B[2][26] +
                  mat_A[13][3] * mat_B[3][26] +
                  mat_A[13][4] * mat_B[4][26] +
                  mat_A[13][5] * mat_B[5][26] +
                  mat_A[13][6] * mat_B[6][26] +
                  mat_A[13][7] * mat_B[7][26] +
                  mat_A[13][8] * mat_B[8][26] +
                  mat_A[13][9] * mat_B[9][26] +
                  mat_A[13][10] * mat_B[10][26] +
                  mat_A[13][11] * mat_B[11][26] +
                  mat_A[13][12] * mat_B[12][26] +
                  mat_A[13][13] * mat_B[13][26] +
                  mat_A[13][14] * mat_B[14][26] +
                  mat_A[13][15] * mat_B[15][26] +
                  mat_A[13][16] * mat_B[16][26] +
                  mat_A[13][17] * mat_B[17][26] +
                  mat_A[13][18] * mat_B[18][26] +
                  mat_A[13][19] * mat_B[19][26] +
                  mat_A[13][20] * mat_B[20][26] +
                  mat_A[13][21] * mat_B[21][26] +
                  mat_A[13][22] * mat_B[22][26] +
                  mat_A[13][23] * mat_B[23][26] +
                  mat_A[13][24] * mat_B[24][26] +
                  mat_A[13][25] * mat_B[25][26] +
                  mat_A[13][26] * mat_B[26][26] +
                  mat_A[13][27] * mat_B[27][26] +
                  mat_A[13][28] * mat_B[28][26] +
                  mat_A[13][29] * mat_B[29][26] +
                  mat_A[13][30] * mat_B[30][26] +
                  mat_A[13][31] * mat_B[31][26];
    mat_C[13][27] <= 
                  mat_A[13][0] * mat_B[0][27] +
                  mat_A[13][1] * mat_B[1][27] +
                  mat_A[13][2] * mat_B[2][27] +
                  mat_A[13][3] * mat_B[3][27] +
                  mat_A[13][4] * mat_B[4][27] +
                  mat_A[13][5] * mat_B[5][27] +
                  mat_A[13][6] * mat_B[6][27] +
                  mat_A[13][7] * mat_B[7][27] +
                  mat_A[13][8] * mat_B[8][27] +
                  mat_A[13][9] * mat_B[9][27] +
                  mat_A[13][10] * mat_B[10][27] +
                  mat_A[13][11] * mat_B[11][27] +
                  mat_A[13][12] * mat_B[12][27] +
                  mat_A[13][13] * mat_B[13][27] +
                  mat_A[13][14] * mat_B[14][27] +
                  mat_A[13][15] * mat_B[15][27] +
                  mat_A[13][16] * mat_B[16][27] +
                  mat_A[13][17] * mat_B[17][27] +
                  mat_A[13][18] * mat_B[18][27] +
                  mat_A[13][19] * mat_B[19][27] +
                  mat_A[13][20] * mat_B[20][27] +
                  mat_A[13][21] * mat_B[21][27] +
                  mat_A[13][22] * mat_B[22][27] +
                  mat_A[13][23] * mat_B[23][27] +
                  mat_A[13][24] * mat_B[24][27] +
                  mat_A[13][25] * mat_B[25][27] +
                  mat_A[13][26] * mat_B[26][27] +
                  mat_A[13][27] * mat_B[27][27] +
                  mat_A[13][28] * mat_B[28][27] +
                  mat_A[13][29] * mat_B[29][27] +
                  mat_A[13][30] * mat_B[30][27] +
                  mat_A[13][31] * mat_B[31][27];
    mat_C[13][28] <= 
                  mat_A[13][0] * mat_B[0][28] +
                  mat_A[13][1] * mat_B[1][28] +
                  mat_A[13][2] * mat_B[2][28] +
                  mat_A[13][3] * mat_B[3][28] +
                  mat_A[13][4] * mat_B[4][28] +
                  mat_A[13][5] * mat_B[5][28] +
                  mat_A[13][6] * mat_B[6][28] +
                  mat_A[13][7] * mat_B[7][28] +
                  mat_A[13][8] * mat_B[8][28] +
                  mat_A[13][9] * mat_B[9][28] +
                  mat_A[13][10] * mat_B[10][28] +
                  mat_A[13][11] * mat_B[11][28] +
                  mat_A[13][12] * mat_B[12][28] +
                  mat_A[13][13] * mat_B[13][28] +
                  mat_A[13][14] * mat_B[14][28] +
                  mat_A[13][15] * mat_B[15][28] +
                  mat_A[13][16] * mat_B[16][28] +
                  mat_A[13][17] * mat_B[17][28] +
                  mat_A[13][18] * mat_B[18][28] +
                  mat_A[13][19] * mat_B[19][28] +
                  mat_A[13][20] * mat_B[20][28] +
                  mat_A[13][21] * mat_B[21][28] +
                  mat_A[13][22] * mat_B[22][28] +
                  mat_A[13][23] * mat_B[23][28] +
                  mat_A[13][24] * mat_B[24][28] +
                  mat_A[13][25] * mat_B[25][28] +
                  mat_A[13][26] * mat_B[26][28] +
                  mat_A[13][27] * mat_B[27][28] +
                  mat_A[13][28] * mat_B[28][28] +
                  mat_A[13][29] * mat_B[29][28] +
                  mat_A[13][30] * mat_B[30][28] +
                  mat_A[13][31] * mat_B[31][28];
    mat_C[13][29] <= 
                  mat_A[13][0] * mat_B[0][29] +
                  mat_A[13][1] * mat_B[1][29] +
                  mat_A[13][2] * mat_B[2][29] +
                  mat_A[13][3] * mat_B[3][29] +
                  mat_A[13][4] * mat_B[4][29] +
                  mat_A[13][5] * mat_B[5][29] +
                  mat_A[13][6] * mat_B[6][29] +
                  mat_A[13][7] * mat_B[7][29] +
                  mat_A[13][8] * mat_B[8][29] +
                  mat_A[13][9] * mat_B[9][29] +
                  mat_A[13][10] * mat_B[10][29] +
                  mat_A[13][11] * mat_B[11][29] +
                  mat_A[13][12] * mat_B[12][29] +
                  mat_A[13][13] * mat_B[13][29] +
                  mat_A[13][14] * mat_B[14][29] +
                  mat_A[13][15] * mat_B[15][29] +
                  mat_A[13][16] * mat_B[16][29] +
                  mat_A[13][17] * mat_B[17][29] +
                  mat_A[13][18] * mat_B[18][29] +
                  mat_A[13][19] * mat_B[19][29] +
                  mat_A[13][20] * mat_B[20][29] +
                  mat_A[13][21] * mat_B[21][29] +
                  mat_A[13][22] * mat_B[22][29] +
                  mat_A[13][23] * mat_B[23][29] +
                  mat_A[13][24] * mat_B[24][29] +
                  mat_A[13][25] * mat_B[25][29] +
                  mat_A[13][26] * mat_B[26][29] +
                  mat_A[13][27] * mat_B[27][29] +
                  mat_A[13][28] * mat_B[28][29] +
                  mat_A[13][29] * mat_B[29][29] +
                  mat_A[13][30] * mat_B[30][29] +
                  mat_A[13][31] * mat_B[31][29];
    mat_C[13][30] <= 
                  mat_A[13][0] * mat_B[0][30] +
                  mat_A[13][1] * mat_B[1][30] +
                  mat_A[13][2] * mat_B[2][30] +
                  mat_A[13][3] * mat_B[3][30] +
                  mat_A[13][4] * mat_B[4][30] +
                  mat_A[13][5] * mat_B[5][30] +
                  mat_A[13][6] * mat_B[6][30] +
                  mat_A[13][7] * mat_B[7][30] +
                  mat_A[13][8] * mat_B[8][30] +
                  mat_A[13][9] * mat_B[9][30] +
                  mat_A[13][10] * mat_B[10][30] +
                  mat_A[13][11] * mat_B[11][30] +
                  mat_A[13][12] * mat_B[12][30] +
                  mat_A[13][13] * mat_B[13][30] +
                  mat_A[13][14] * mat_B[14][30] +
                  mat_A[13][15] * mat_B[15][30] +
                  mat_A[13][16] * mat_B[16][30] +
                  mat_A[13][17] * mat_B[17][30] +
                  mat_A[13][18] * mat_B[18][30] +
                  mat_A[13][19] * mat_B[19][30] +
                  mat_A[13][20] * mat_B[20][30] +
                  mat_A[13][21] * mat_B[21][30] +
                  mat_A[13][22] * mat_B[22][30] +
                  mat_A[13][23] * mat_B[23][30] +
                  mat_A[13][24] * mat_B[24][30] +
                  mat_A[13][25] * mat_B[25][30] +
                  mat_A[13][26] * mat_B[26][30] +
                  mat_A[13][27] * mat_B[27][30] +
                  mat_A[13][28] * mat_B[28][30] +
                  mat_A[13][29] * mat_B[29][30] +
                  mat_A[13][30] * mat_B[30][30] +
                  mat_A[13][31] * mat_B[31][30];
    mat_C[13][31] <= 
                  mat_A[13][0] * mat_B[0][31] +
                  mat_A[13][1] * mat_B[1][31] +
                  mat_A[13][2] * mat_B[2][31] +
                  mat_A[13][3] * mat_B[3][31] +
                  mat_A[13][4] * mat_B[4][31] +
                  mat_A[13][5] * mat_B[5][31] +
                  mat_A[13][6] * mat_B[6][31] +
                  mat_A[13][7] * mat_B[7][31] +
                  mat_A[13][8] * mat_B[8][31] +
                  mat_A[13][9] * mat_B[9][31] +
                  mat_A[13][10] * mat_B[10][31] +
                  mat_A[13][11] * mat_B[11][31] +
                  mat_A[13][12] * mat_B[12][31] +
                  mat_A[13][13] * mat_B[13][31] +
                  mat_A[13][14] * mat_B[14][31] +
                  mat_A[13][15] * mat_B[15][31] +
                  mat_A[13][16] * mat_B[16][31] +
                  mat_A[13][17] * mat_B[17][31] +
                  mat_A[13][18] * mat_B[18][31] +
                  mat_A[13][19] * mat_B[19][31] +
                  mat_A[13][20] * mat_B[20][31] +
                  mat_A[13][21] * mat_B[21][31] +
                  mat_A[13][22] * mat_B[22][31] +
                  mat_A[13][23] * mat_B[23][31] +
                  mat_A[13][24] * mat_B[24][31] +
                  mat_A[13][25] * mat_B[25][31] +
                  mat_A[13][26] * mat_B[26][31] +
                  mat_A[13][27] * mat_B[27][31] +
                  mat_A[13][28] * mat_B[28][31] +
                  mat_A[13][29] * mat_B[29][31] +
                  mat_A[13][30] * mat_B[30][31] +
                  mat_A[13][31] * mat_B[31][31];
    mat_C[14][0] <= 
                  mat_A[14][0] * mat_B[0][0] +
                  mat_A[14][1] * mat_B[1][0] +
                  mat_A[14][2] * mat_B[2][0] +
                  mat_A[14][3] * mat_B[3][0] +
                  mat_A[14][4] * mat_B[4][0] +
                  mat_A[14][5] * mat_B[5][0] +
                  mat_A[14][6] * mat_B[6][0] +
                  mat_A[14][7] * mat_B[7][0] +
                  mat_A[14][8] * mat_B[8][0] +
                  mat_A[14][9] * mat_B[9][0] +
                  mat_A[14][10] * mat_B[10][0] +
                  mat_A[14][11] * mat_B[11][0] +
                  mat_A[14][12] * mat_B[12][0] +
                  mat_A[14][13] * mat_B[13][0] +
                  mat_A[14][14] * mat_B[14][0] +
                  mat_A[14][15] * mat_B[15][0] +
                  mat_A[14][16] * mat_B[16][0] +
                  mat_A[14][17] * mat_B[17][0] +
                  mat_A[14][18] * mat_B[18][0] +
                  mat_A[14][19] * mat_B[19][0] +
                  mat_A[14][20] * mat_B[20][0] +
                  mat_A[14][21] * mat_B[21][0] +
                  mat_A[14][22] * mat_B[22][0] +
                  mat_A[14][23] * mat_B[23][0] +
                  mat_A[14][24] * mat_B[24][0] +
                  mat_A[14][25] * mat_B[25][0] +
                  mat_A[14][26] * mat_B[26][0] +
                  mat_A[14][27] * mat_B[27][0] +
                  mat_A[14][28] * mat_B[28][0] +
                  mat_A[14][29] * mat_B[29][0] +
                  mat_A[14][30] * mat_B[30][0] +
                  mat_A[14][31] * mat_B[31][0];
    mat_C[14][1] <= 
                  mat_A[14][0] * mat_B[0][1] +
                  mat_A[14][1] * mat_B[1][1] +
                  mat_A[14][2] * mat_B[2][1] +
                  mat_A[14][3] * mat_B[3][1] +
                  mat_A[14][4] * mat_B[4][1] +
                  mat_A[14][5] * mat_B[5][1] +
                  mat_A[14][6] * mat_B[6][1] +
                  mat_A[14][7] * mat_B[7][1] +
                  mat_A[14][8] * mat_B[8][1] +
                  mat_A[14][9] * mat_B[9][1] +
                  mat_A[14][10] * mat_B[10][1] +
                  mat_A[14][11] * mat_B[11][1] +
                  mat_A[14][12] * mat_B[12][1] +
                  mat_A[14][13] * mat_B[13][1] +
                  mat_A[14][14] * mat_B[14][1] +
                  mat_A[14][15] * mat_B[15][1] +
                  mat_A[14][16] * mat_B[16][1] +
                  mat_A[14][17] * mat_B[17][1] +
                  mat_A[14][18] * mat_B[18][1] +
                  mat_A[14][19] * mat_B[19][1] +
                  mat_A[14][20] * mat_B[20][1] +
                  mat_A[14][21] * mat_B[21][1] +
                  mat_A[14][22] * mat_B[22][1] +
                  mat_A[14][23] * mat_B[23][1] +
                  mat_A[14][24] * mat_B[24][1] +
                  mat_A[14][25] * mat_B[25][1] +
                  mat_A[14][26] * mat_B[26][1] +
                  mat_A[14][27] * mat_B[27][1] +
                  mat_A[14][28] * mat_B[28][1] +
                  mat_A[14][29] * mat_B[29][1] +
                  mat_A[14][30] * mat_B[30][1] +
                  mat_A[14][31] * mat_B[31][1];
    mat_C[14][2] <= 
                  mat_A[14][0] * mat_B[0][2] +
                  mat_A[14][1] * mat_B[1][2] +
                  mat_A[14][2] * mat_B[2][2] +
                  mat_A[14][3] * mat_B[3][2] +
                  mat_A[14][4] * mat_B[4][2] +
                  mat_A[14][5] * mat_B[5][2] +
                  mat_A[14][6] * mat_B[6][2] +
                  mat_A[14][7] * mat_B[7][2] +
                  mat_A[14][8] * mat_B[8][2] +
                  mat_A[14][9] * mat_B[9][2] +
                  mat_A[14][10] * mat_B[10][2] +
                  mat_A[14][11] * mat_B[11][2] +
                  mat_A[14][12] * mat_B[12][2] +
                  mat_A[14][13] * mat_B[13][2] +
                  mat_A[14][14] * mat_B[14][2] +
                  mat_A[14][15] * mat_B[15][2] +
                  mat_A[14][16] * mat_B[16][2] +
                  mat_A[14][17] * mat_B[17][2] +
                  mat_A[14][18] * mat_B[18][2] +
                  mat_A[14][19] * mat_B[19][2] +
                  mat_A[14][20] * mat_B[20][2] +
                  mat_A[14][21] * mat_B[21][2] +
                  mat_A[14][22] * mat_B[22][2] +
                  mat_A[14][23] * mat_B[23][2] +
                  mat_A[14][24] * mat_B[24][2] +
                  mat_A[14][25] * mat_B[25][2] +
                  mat_A[14][26] * mat_B[26][2] +
                  mat_A[14][27] * mat_B[27][2] +
                  mat_A[14][28] * mat_B[28][2] +
                  mat_A[14][29] * mat_B[29][2] +
                  mat_A[14][30] * mat_B[30][2] +
                  mat_A[14][31] * mat_B[31][2];
    mat_C[14][3] <= 
                  mat_A[14][0] * mat_B[0][3] +
                  mat_A[14][1] * mat_B[1][3] +
                  mat_A[14][2] * mat_B[2][3] +
                  mat_A[14][3] * mat_B[3][3] +
                  mat_A[14][4] * mat_B[4][3] +
                  mat_A[14][5] * mat_B[5][3] +
                  mat_A[14][6] * mat_B[6][3] +
                  mat_A[14][7] * mat_B[7][3] +
                  mat_A[14][8] * mat_B[8][3] +
                  mat_A[14][9] * mat_B[9][3] +
                  mat_A[14][10] * mat_B[10][3] +
                  mat_A[14][11] * mat_B[11][3] +
                  mat_A[14][12] * mat_B[12][3] +
                  mat_A[14][13] * mat_B[13][3] +
                  mat_A[14][14] * mat_B[14][3] +
                  mat_A[14][15] * mat_B[15][3] +
                  mat_A[14][16] * mat_B[16][3] +
                  mat_A[14][17] * mat_B[17][3] +
                  mat_A[14][18] * mat_B[18][3] +
                  mat_A[14][19] * mat_B[19][3] +
                  mat_A[14][20] * mat_B[20][3] +
                  mat_A[14][21] * mat_B[21][3] +
                  mat_A[14][22] * mat_B[22][3] +
                  mat_A[14][23] * mat_B[23][3] +
                  mat_A[14][24] * mat_B[24][3] +
                  mat_A[14][25] * mat_B[25][3] +
                  mat_A[14][26] * mat_B[26][3] +
                  mat_A[14][27] * mat_B[27][3] +
                  mat_A[14][28] * mat_B[28][3] +
                  mat_A[14][29] * mat_B[29][3] +
                  mat_A[14][30] * mat_B[30][3] +
                  mat_A[14][31] * mat_B[31][3];
    mat_C[14][4] <= 
                  mat_A[14][0] * mat_B[0][4] +
                  mat_A[14][1] * mat_B[1][4] +
                  mat_A[14][2] * mat_B[2][4] +
                  mat_A[14][3] * mat_B[3][4] +
                  mat_A[14][4] * mat_B[4][4] +
                  mat_A[14][5] * mat_B[5][4] +
                  mat_A[14][6] * mat_B[6][4] +
                  mat_A[14][7] * mat_B[7][4] +
                  mat_A[14][8] * mat_B[8][4] +
                  mat_A[14][9] * mat_B[9][4] +
                  mat_A[14][10] * mat_B[10][4] +
                  mat_A[14][11] * mat_B[11][4] +
                  mat_A[14][12] * mat_B[12][4] +
                  mat_A[14][13] * mat_B[13][4] +
                  mat_A[14][14] * mat_B[14][4] +
                  mat_A[14][15] * mat_B[15][4] +
                  mat_A[14][16] * mat_B[16][4] +
                  mat_A[14][17] * mat_B[17][4] +
                  mat_A[14][18] * mat_B[18][4] +
                  mat_A[14][19] * mat_B[19][4] +
                  mat_A[14][20] * mat_B[20][4] +
                  mat_A[14][21] * mat_B[21][4] +
                  mat_A[14][22] * mat_B[22][4] +
                  mat_A[14][23] * mat_B[23][4] +
                  mat_A[14][24] * mat_B[24][4] +
                  mat_A[14][25] * mat_B[25][4] +
                  mat_A[14][26] * mat_B[26][4] +
                  mat_A[14][27] * mat_B[27][4] +
                  mat_A[14][28] * mat_B[28][4] +
                  mat_A[14][29] * mat_B[29][4] +
                  mat_A[14][30] * mat_B[30][4] +
                  mat_A[14][31] * mat_B[31][4];
    mat_C[14][5] <= 
                  mat_A[14][0] * mat_B[0][5] +
                  mat_A[14][1] * mat_B[1][5] +
                  mat_A[14][2] * mat_B[2][5] +
                  mat_A[14][3] * mat_B[3][5] +
                  mat_A[14][4] * mat_B[4][5] +
                  mat_A[14][5] * mat_B[5][5] +
                  mat_A[14][6] * mat_B[6][5] +
                  mat_A[14][7] * mat_B[7][5] +
                  mat_A[14][8] * mat_B[8][5] +
                  mat_A[14][9] * mat_B[9][5] +
                  mat_A[14][10] * mat_B[10][5] +
                  mat_A[14][11] * mat_B[11][5] +
                  mat_A[14][12] * mat_B[12][5] +
                  mat_A[14][13] * mat_B[13][5] +
                  mat_A[14][14] * mat_B[14][5] +
                  mat_A[14][15] * mat_B[15][5] +
                  mat_A[14][16] * mat_B[16][5] +
                  mat_A[14][17] * mat_B[17][5] +
                  mat_A[14][18] * mat_B[18][5] +
                  mat_A[14][19] * mat_B[19][5] +
                  mat_A[14][20] * mat_B[20][5] +
                  mat_A[14][21] * mat_B[21][5] +
                  mat_A[14][22] * mat_B[22][5] +
                  mat_A[14][23] * mat_B[23][5] +
                  mat_A[14][24] * mat_B[24][5] +
                  mat_A[14][25] * mat_B[25][5] +
                  mat_A[14][26] * mat_B[26][5] +
                  mat_A[14][27] * mat_B[27][5] +
                  mat_A[14][28] * mat_B[28][5] +
                  mat_A[14][29] * mat_B[29][5] +
                  mat_A[14][30] * mat_B[30][5] +
                  mat_A[14][31] * mat_B[31][5];
    mat_C[14][6] <= 
                  mat_A[14][0] * mat_B[0][6] +
                  mat_A[14][1] * mat_B[1][6] +
                  mat_A[14][2] * mat_B[2][6] +
                  mat_A[14][3] * mat_B[3][6] +
                  mat_A[14][4] * mat_B[4][6] +
                  mat_A[14][5] * mat_B[5][6] +
                  mat_A[14][6] * mat_B[6][6] +
                  mat_A[14][7] * mat_B[7][6] +
                  mat_A[14][8] * mat_B[8][6] +
                  mat_A[14][9] * mat_B[9][6] +
                  mat_A[14][10] * mat_B[10][6] +
                  mat_A[14][11] * mat_B[11][6] +
                  mat_A[14][12] * mat_B[12][6] +
                  mat_A[14][13] * mat_B[13][6] +
                  mat_A[14][14] * mat_B[14][6] +
                  mat_A[14][15] * mat_B[15][6] +
                  mat_A[14][16] * mat_B[16][6] +
                  mat_A[14][17] * mat_B[17][6] +
                  mat_A[14][18] * mat_B[18][6] +
                  mat_A[14][19] * mat_B[19][6] +
                  mat_A[14][20] * mat_B[20][6] +
                  mat_A[14][21] * mat_B[21][6] +
                  mat_A[14][22] * mat_B[22][6] +
                  mat_A[14][23] * mat_B[23][6] +
                  mat_A[14][24] * mat_B[24][6] +
                  mat_A[14][25] * mat_B[25][6] +
                  mat_A[14][26] * mat_B[26][6] +
                  mat_A[14][27] * mat_B[27][6] +
                  mat_A[14][28] * mat_B[28][6] +
                  mat_A[14][29] * mat_B[29][6] +
                  mat_A[14][30] * mat_B[30][6] +
                  mat_A[14][31] * mat_B[31][6];
    mat_C[14][7] <= 
                  mat_A[14][0] * mat_B[0][7] +
                  mat_A[14][1] * mat_B[1][7] +
                  mat_A[14][2] * mat_B[2][7] +
                  mat_A[14][3] * mat_B[3][7] +
                  mat_A[14][4] * mat_B[4][7] +
                  mat_A[14][5] * mat_B[5][7] +
                  mat_A[14][6] * mat_B[6][7] +
                  mat_A[14][7] * mat_B[7][7] +
                  mat_A[14][8] * mat_B[8][7] +
                  mat_A[14][9] * mat_B[9][7] +
                  mat_A[14][10] * mat_B[10][7] +
                  mat_A[14][11] * mat_B[11][7] +
                  mat_A[14][12] * mat_B[12][7] +
                  mat_A[14][13] * mat_B[13][7] +
                  mat_A[14][14] * mat_B[14][7] +
                  mat_A[14][15] * mat_B[15][7] +
                  mat_A[14][16] * mat_B[16][7] +
                  mat_A[14][17] * mat_B[17][7] +
                  mat_A[14][18] * mat_B[18][7] +
                  mat_A[14][19] * mat_B[19][7] +
                  mat_A[14][20] * mat_B[20][7] +
                  mat_A[14][21] * mat_B[21][7] +
                  mat_A[14][22] * mat_B[22][7] +
                  mat_A[14][23] * mat_B[23][7] +
                  mat_A[14][24] * mat_B[24][7] +
                  mat_A[14][25] * mat_B[25][7] +
                  mat_A[14][26] * mat_B[26][7] +
                  mat_A[14][27] * mat_B[27][7] +
                  mat_A[14][28] * mat_B[28][7] +
                  mat_A[14][29] * mat_B[29][7] +
                  mat_A[14][30] * mat_B[30][7] +
                  mat_A[14][31] * mat_B[31][7];
    mat_C[14][8] <= 
                  mat_A[14][0] * mat_B[0][8] +
                  mat_A[14][1] * mat_B[1][8] +
                  mat_A[14][2] * mat_B[2][8] +
                  mat_A[14][3] * mat_B[3][8] +
                  mat_A[14][4] * mat_B[4][8] +
                  mat_A[14][5] * mat_B[5][8] +
                  mat_A[14][6] * mat_B[6][8] +
                  mat_A[14][7] * mat_B[7][8] +
                  mat_A[14][8] * mat_B[8][8] +
                  mat_A[14][9] * mat_B[9][8] +
                  mat_A[14][10] * mat_B[10][8] +
                  mat_A[14][11] * mat_B[11][8] +
                  mat_A[14][12] * mat_B[12][8] +
                  mat_A[14][13] * mat_B[13][8] +
                  mat_A[14][14] * mat_B[14][8] +
                  mat_A[14][15] * mat_B[15][8] +
                  mat_A[14][16] * mat_B[16][8] +
                  mat_A[14][17] * mat_B[17][8] +
                  mat_A[14][18] * mat_B[18][8] +
                  mat_A[14][19] * mat_B[19][8] +
                  mat_A[14][20] * mat_B[20][8] +
                  mat_A[14][21] * mat_B[21][8] +
                  mat_A[14][22] * mat_B[22][8] +
                  mat_A[14][23] * mat_B[23][8] +
                  mat_A[14][24] * mat_B[24][8] +
                  mat_A[14][25] * mat_B[25][8] +
                  mat_A[14][26] * mat_B[26][8] +
                  mat_A[14][27] * mat_B[27][8] +
                  mat_A[14][28] * mat_B[28][8] +
                  mat_A[14][29] * mat_B[29][8] +
                  mat_A[14][30] * mat_B[30][8] +
                  mat_A[14][31] * mat_B[31][8];
    mat_C[14][9] <= 
                  mat_A[14][0] * mat_B[0][9] +
                  mat_A[14][1] * mat_B[1][9] +
                  mat_A[14][2] * mat_B[2][9] +
                  mat_A[14][3] * mat_B[3][9] +
                  mat_A[14][4] * mat_B[4][9] +
                  mat_A[14][5] * mat_B[5][9] +
                  mat_A[14][6] * mat_B[6][9] +
                  mat_A[14][7] * mat_B[7][9] +
                  mat_A[14][8] * mat_B[8][9] +
                  mat_A[14][9] * mat_B[9][9] +
                  mat_A[14][10] * mat_B[10][9] +
                  mat_A[14][11] * mat_B[11][9] +
                  mat_A[14][12] * mat_B[12][9] +
                  mat_A[14][13] * mat_B[13][9] +
                  mat_A[14][14] * mat_B[14][9] +
                  mat_A[14][15] * mat_B[15][9] +
                  mat_A[14][16] * mat_B[16][9] +
                  mat_A[14][17] * mat_B[17][9] +
                  mat_A[14][18] * mat_B[18][9] +
                  mat_A[14][19] * mat_B[19][9] +
                  mat_A[14][20] * mat_B[20][9] +
                  mat_A[14][21] * mat_B[21][9] +
                  mat_A[14][22] * mat_B[22][9] +
                  mat_A[14][23] * mat_B[23][9] +
                  mat_A[14][24] * mat_B[24][9] +
                  mat_A[14][25] * mat_B[25][9] +
                  mat_A[14][26] * mat_B[26][9] +
                  mat_A[14][27] * mat_B[27][9] +
                  mat_A[14][28] * mat_B[28][9] +
                  mat_A[14][29] * mat_B[29][9] +
                  mat_A[14][30] * mat_B[30][9] +
                  mat_A[14][31] * mat_B[31][9];
    mat_C[14][10] <= 
                  mat_A[14][0] * mat_B[0][10] +
                  mat_A[14][1] * mat_B[1][10] +
                  mat_A[14][2] * mat_B[2][10] +
                  mat_A[14][3] * mat_B[3][10] +
                  mat_A[14][4] * mat_B[4][10] +
                  mat_A[14][5] * mat_B[5][10] +
                  mat_A[14][6] * mat_B[6][10] +
                  mat_A[14][7] * mat_B[7][10] +
                  mat_A[14][8] * mat_B[8][10] +
                  mat_A[14][9] * mat_B[9][10] +
                  mat_A[14][10] * mat_B[10][10] +
                  mat_A[14][11] * mat_B[11][10] +
                  mat_A[14][12] * mat_B[12][10] +
                  mat_A[14][13] * mat_B[13][10] +
                  mat_A[14][14] * mat_B[14][10] +
                  mat_A[14][15] * mat_B[15][10] +
                  mat_A[14][16] * mat_B[16][10] +
                  mat_A[14][17] * mat_B[17][10] +
                  mat_A[14][18] * mat_B[18][10] +
                  mat_A[14][19] * mat_B[19][10] +
                  mat_A[14][20] * mat_B[20][10] +
                  mat_A[14][21] * mat_B[21][10] +
                  mat_A[14][22] * mat_B[22][10] +
                  mat_A[14][23] * mat_B[23][10] +
                  mat_A[14][24] * mat_B[24][10] +
                  mat_A[14][25] * mat_B[25][10] +
                  mat_A[14][26] * mat_B[26][10] +
                  mat_A[14][27] * mat_B[27][10] +
                  mat_A[14][28] * mat_B[28][10] +
                  mat_A[14][29] * mat_B[29][10] +
                  mat_A[14][30] * mat_B[30][10] +
                  mat_A[14][31] * mat_B[31][10];
    mat_C[14][11] <= 
                  mat_A[14][0] * mat_B[0][11] +
                  mat_A[14][1] * mat_B[1][11] +
                  mat_A[14][2] * mat_B[2][11] +
                  mat_A[14][3] * mat_B[3][11] +
                  mat_A[14][4] * mat_B[4][11] +
                  mat_A[14][5] * mat_B[5][11] +
                  mat_A[14][6] * mat_B[6][11] +
                  mat_A[14][7] * mat_B[7][11] +
                  mat_A[14][8] * mat_B[8][11] +
                  mat_A[14][9] * mat_B[9][11] +
                  mat_A[14][10] * mat_B[10][11] +
                  mat_A[14][11] * mat_B[11][11] +
                  mat_A[14][12] * mat_B[12][11] +
                  mat_A[14][13] * mat_B[13][11] +
                  mat_A[14][14] * mat_B[14][11] +
                  mat_A[14][15] * mat_B[15][11] +
                  mat_A[14][16] * mat_B[16][11] +
                  mat_A[14][17] * mat_B[17][11] +
                  mat_A[14][18] * mat_B[18][11] +
                  mat_A[14][19] * mat_B[19][11] +
                  mat_A[14][20] * mat_B[20][11] +
                  mat_A[14][21] * mat_B[21][11] +
                  mat_A[14][22] * mat_B[22][11] +
                  mat_A[14][23] * mat_B[23][11] +
                  mat_A[14][24] * mat_B[24][11] +
                  mat_A[14][25] * mat_B[25][11] +
                  mat_A[14][26] * mat_B[26][11] +
                  mat_A[14][27] * mat_B[27][11] +
                  mat_A[14][28] * mat_B[28][11] +
                  mat_A[14][29] * mat_B[29][11] +
                  mat_A[14][30] * mat_B[30][11] +
                  mat_A[14][31] * mat_B[31][11];
    mat_C[14][12] <= 
                  mat_A[14][0] * mat_B[0][12] +
                  mat_A[14][1] * mat_B[1][12] +
                  mat_A[14][2] * mat_B[2][12] +
                  mat_A[14][3] * mat_B[3][12] +
                  mat_A[14][4] * mat_B[4][12] +
                  mat_A[14][5] * mat_B[5][12] +
                  mat_A[14][6] * mat_B[6][12] +
                  mat_A[14][7] * mat_B[7][12] +
                  mat_A[14][8] * mat_B[8][12] +
                  mat_A[14][9] * mat_B[9][12] +
                  mat_A[14][10] * mat_B[10][12] +
                  mat_A[14][11] * mat_B[11][12] +
                  mat_A[14][12] * mat_B[12][12] +
                  mat_A[14][13] * mat_B[13][12] +
                  mat_A[14][14] * mat_B[14][12] +
                  mat_A[14][15] * mat_B[15][12] +
                  mat_A[14][16] * mat_B[16][12] +
                  mat_A[14][17] * mat_B[17][12] +
                  mat_A[14][18] * mat_B[18][12] +
                  mat_A[14][19] * mat_B[19][12] +
                  mat_A[14][20] * mat_B[20][12] +
                  mat_A[14][21] * mat_B[21][12] +
                  mat_A[14][22] * mat_B[22][12] +
                  mat_A[14][23] * mat_B[23][12] +
                  mat_A[14][24] * mat_B[24][12] +
                  mat_A[14][25] * mat_B[25][12] +
                  mat_A[14][26] * mat_B[26][12] +
                  mat_A[14][27] * mat_B[27][12] +
                  mat_A[14][28] * mat_B[28][12] +
                  mat_A[14][29] * mat_B[29][12] +
                  mat_A[14][30] * mat_B[30][12] +
                  mat_A[14][31] * mat_B[31][12];
    mat_C[14][13] <= 
                  mat_A[14][0] * mat_B[0][13] +
                  mat_A[14][1] * mat_B[1][13] +
                  mat_A[14][2] * mat_B[2][13] +
                  mat_A[14][3] * mat_B[3][13] +
                  mat_A[14][4] * mat_B[4][13] +
                  mat_A[14][5] * mat_B[5][13] +
                  mat_A[14][6] * mat_B[6][13] +
                  mat_A[14][7] * mat_B[7][13] +
                  mat_A[14][8] * mat_B[8][13] +
                  mat_A[14][9] * mat_B[9][13] +
                  mat_A[14][10] * mat_B[10][13] +
                  mat_A[14][11] * mat_B[11][13] +
                  mat_A[14][12] * mat_B[12][13] +
                  mat_A[14][13] * mat_B[13][13] +
                  mat_A[14][14] * mat_B[14][13] +
                  mat_A[14][15] * mat_B[15][13] +
                  mat_A[14][16] * mat_B[16][13] +
                  mat_A[14][17] * mat_B[17][13] +
                  mat_A[14][18] * mat_B[18][13] +
                  mat_A[14][19] * mat_B[19][13] +
                  mat_A[14][20] * mat_B[20][13] +
                  mat_A[14][21] * mat_B[21][13] +
                  mat_A[14][22] * mat_B[22][13] +
                  mat_A[14][23] * mat_B[23][13] +
                  mat_A[14][24] * mat_B[24][13] +
                  mat_A[14][25] * mat_B[25][13] +
                  mat_A[14][26] * mat_B[26][13] +
                  mat_A[14][27] * mat_B[27][13] +
                  mat_A[14][28] * mat_B[28][13] +
                  mat_A[14][29] * mat_B[29][13] +
                  mat_A[14][30] * mat_B[30][13] +
                  mat_A[14][31] * mat_B[31][13];
    mat_C[14][14] <= 
                  mat_A[14][0] * mat_B[0][14] +
                  mat_A[14][1] * mat_B[1][14] +
                  mat_A[14][2] * mat_B[2][14] +
                  mat_A[14][3] * mat_B[3][14] +
                  mat_A[14][4] * mat_B[4][14] +
                  mat_A[14][5] * mat_B[5][14] +
                  mat_A[14][6] * mat_B[6][14] +
                  mat_A[14][7] * mat_B[7][14] +
                  mat_A[14][8] * mat_B[8][14] +
                  mat_A[14][9] * mat_B[9][14] +
                  mat_A[14][10] * mat_B[10][14] +
                  mat_A[14][11] * mat_B[11][14] +
                  mat_A[14][12] * mat_B[12][14] +
                  mat_A[14][13] * mat_B[13][14] +
                  mat_A[14][14] * mat_B[14][14] +
                  mat_A[14][15] * mat_B[15][14] +
                  mat_A[14][16] * mat_B[16][14] +
                  mat_A[14][17] * mat_B[17][14] +
                  mat_A[14][18] * mat_B[18][14] +
                  mat_A[14][19] * mat_B[19][14] +
                  mat_A[14][20] * mat_B[20][14] +
                  mat_A[14][21] * mat_B[21][14] +
                  mat_A[14][22] * mat_B[22][14] +
                  mat_A[14][23] * mat_B[23][14] +
                  mat_A[14][24] * mat_B[24][14] +
                  mat_A[14][25] * mat_B[25][14] +
                  mat_A[14][26] * mat_B[26][14] +
                  mat_A[14][27] * mat_B[27][14] +
                  mat_A[14][28] * mat_B[28][14] +
                  mat_A[14][29] * mat_B[29][14] +
                  mat_A[14][30] * mat_B[30][14] +
                  mat_A[14][31] * mat_B[31][14];
    mat_C[14][15] <= 
                  mat_A[14][0] * mat_B[0][15] +
                  mat_A[14][1] * mat_B[1][15] +
                  mat_A[14][2] * mat_B[2][15] +
                  mat_A[14][3] * mat_B[3][15] +
                  mat_A[14][4] * mat_B[4][15] +
                  mat_A[14][5] * mat_B[5][15] +
                  mat_A[14][6] * mat_B[6][15] +
                  mat_A[14][7] * mat_B[7][15] +
                  mat_A[14][8] * mat_B[8][15] +
                  mat_A[14][9] * mat_B[9][15] +
                  mat_A[14][10] * mat_B[10][15] +
                  mat_A[14][11] * mat_B[11][15] +
                  mat_A[14][12] * mat_B[12][15] +
                  mat_A[14][13] * mat_B[13][15] +
                  mat_A[14][14] * mat_B[14][15] +
                  mat_A[14][15] * mat_B[15][15] +
                  mat_A[14][16] * mat_B[16][15] +
                  mat_A[14][17] * mat_B[17][15] +
                  mat_A[14][18] * mat_B[18][15] +
                  mat_A[14][19] * mat_B[19][15] +
                  mat_A[14][20] * mat_B[20][15] +
                  mat_A[14][21] * mat_B[21][15] +
                  mat_A[14][22] * mat_B[22][15] +
                  mat_A[14][23] * mat_B[23][15] +
                  mat_A[14][24] * mat_B[24][15] +
                  mat_A[14][25] * mat_B[25][15] +
                  mat_A[14][26] * mat_B[26][15] +
                  mat_A[14][27] * mat_B[27][15] +
                  mat_A[14][28] * mat_B[28][15] +
                  mat_A[14][29] * mat_B[29][15] +
                  mat_A[14][30] * mat_B[30][15] +
                  mat_A[14][31] * mat_B[31][15];
    mat_C[14][16] <= 
                  mat_A[14][0] * mat_B[0][16] +
                  mat_A[14][1] * mat_B[1][16] +
                  mat_A[14][2] * mat_B[2][16] +
                  mat_A[14][3] * mat_B[3][16] +
                  mat_A[14][4] * mat_B[4][16] +
                  mat_A[14][5] * mat_B[5][16] +
                  mat_A[14][6] * mat_B[6][16] +
                  mat_A[14][7] * mat_B[7][16] +
                  mat_A[14][8] * mat_B[8][16] +
                  mat_A[14][9] * mat_B[9][16] +
                  mat_A[14][10] * mat_B[10][16] +
                  mat_A[14][11] * mat_B[11][16] +
                  mat_A[14][12] * mat_B[12][16] +
                  mat_A[14][13] * mat_B[13][16] +
                  mat_A[14][14] * mat_B[14][16] +
                  mat_A[14][15] * mat_B[15][16] +
                  mat_A[14][16] * mat_B[16][16] +
                  mat_A[14][17] * mat_B[17][16] +
                  mat_A[14][18] * mat_B[18][16] +
                  mat_A[14][19] * mat_B[19][16] +
                  mat_A[14][20] * mat_B[20][16] +
                  mat_A[14][21] * mat_B[21][16] +
                  mat_A[14][22] * mat_B[22][16] +
                  mat_A[14][23] * mat_B[23][16] +
                  mat_A[14][24] * mat_B[24][16] +
                  mat_A[14][25] * mat_B[25][16] +
                  mat_A[14][26] * mat_B[26][16] +
                  mat_A[14][27] * mat_B[27][16] +
                  mat_A[14][28] * mat_B[28][16] +
                  mat_A[14][29] * mat_B[29][16] +
                  mat_A[14][30] * mat_B[30][16] +
                  mat_A[14][31] * mat_B[31][16];
    mat_C[14][17] <= 
                  mat_A[14][0] * mat_B[0][17] +
                  mat_A[14][1] * mat_B[1][17] +
                  mat_A[14][2] * mat_B[2][17] +
                  mat_A[14][3] * mat_B[3][17] +
                  mat_A[14][4] * mat_B[4][17] +
                  mat_A[14][5] * mat_B[5][17] +
                  mat_A[14][6] * mat_B[6][17] +
                  mat_A[14][7] * mat_B[7][17] +
                  mat_A[14][8] * mat_B[8][17] +
                  mat_A[14][9] * mat_B[9][17] +
                  mat_A[14][10] * mat_B[10][17] +
                  mat_A[14][11] * mat_B[11][17] +
                  mat_A[14][12] * mat_B[12][17] +
                  mat_A[14][13] * mat_B[13][17] +
                  mat_A[14][14] * mat_B[14][17] +
                  mat_A[14][15] * mat_B[15][17] +
                  mat_A[14][16] * mat_B[16][17] +
                  mat_A[14][17] * mat_B[17][17] +
                  mat_A[14][18] * mat_B[18][17] +
                  mat_A[14][19] * mat_B[19][17] +
                  mat_A[14][20] * mat_B[20][17] +
                  mat_A[14][21] * mat_B[21][17] +
                  mat_A[14][22] * mat_B[22][17] +
                  mat_A[14][23] * mat_B[23][17] +
                  mat_A[14][24] * mat_B[24][17] +
                  mat_A[14][25] * mat_B[25][17] +
                  mat_A[14][26] * mat_B[26][17] +
                  mat_A[14][27] * mat_B[27][17] +
                  mat_A[14][28] * mat_B[28][17] +
                  mat_A[14][29] * mat_B[29][17] +
                  mat_A[14][30] * mat_B[30][17] +
                  mat_A[14][31] * mat_B[31][17];
    mat_C[14][18] <= 
                  mat_A[14][0] * mat_B[0][18] +
                  mat_A[14][1] * mat_B[1][18] +
                  mat_A[14][2] * mat_B[2][18] +
                  mat_A[14][3] * mat_B[3][18] +
                  mat_A[14][4] * mat_B[4][18] +
                  mat_A[14][5] * mat_B[5][18] +
                  mat_A[14][6] * mat_B[6][18] +
                  mat_A[14][7] * mat_B[7][18] +
                  mat_A[14][8] * mat_B[8][18] +
                  mat_A[14][9] * mat_B[9][18] +
                  mat_A[14][10] * mat_B[10][18] +
                  mat_A[14][11] * mat_B[11][18] +
                  mat_A[14][12] * mat_B[12][18] +
                  mat_A[14][13] * mat_B[13][18] +
                  mat_A[14][14] * mat_B[14][18] +
                  mat_A[14][15] * mat_B[15][18] +
                  mat_A[14][16] * mat_B[16][18] +
                  mat_A[14][17] * mat_B[17][18] +
                  mat_A[14][18] * mat_B[18][18] +
                  mat_A[14][19] * mat_B[19][18] +
                  mat_A[14][20] * mat_B[20][18] +
                  mat_A[14][21] * mat_B[21][18] +
                  mat_A[14][22] * mat_B[22][18] +
                  mat_A[14][23] * mat_B[23][18] +
                  mat_A[14][24] * mat_B[24][18] +
                  mat_A[14][25] * mat_B[25][18] +
                  mat_A[14][26] * mat_B[26][18] +
                  mat_A[14][27] * mat_B[27][18] +
                  mat_A[14][28] * mat_B[28][18] +
                  mat_A[14][29] * mat_B[29][18] +
                  mat_A[14][30] * mat_B[30][18] +
                  mat_A[14][31] * mat_B[31][18];
    mat_C[14][19] <= 
                  mat_A[14][0] * mat_B[0][19] +
                  mat_A[14][1] * mat_B[1][19] +
                  mat_A[14][2] * mat_B[2][19] +
                  mat_A[14][3] * mat_B[3][19] +
                  mat_A[14][4] * mat_B[4][19] +
                  mat_A[14][5] * mat_B[5][19] +
                  mat_A[14][6] * mat_B[6][19] +
                  mat_A[14][7] * mat_B[7][19] +
                  mat_A[14][8] * mat_B[8][19] +
                  mat_A[14][9] * mat_B[9][19] +
                  mat_A[14][10] * mat_B[10][19] +
                  mat_A[14][11] * mat_B[11][19] +
                  mat_A[14][12] * mat_B[12][19] +
                  mat_A[14][13] * mat_B[13][19] +
                  mat_A[14][14] * mat_B[14][19] +
                  mat_A[14][15] * mat_B[15][19] +
                  mat_A[14][16] * mat_B[16][19] +
                  mat_A[14][17] * mat_B[17][19] +
                  mat_A[14][18] * mat_B[18][19] +
                  mat_A[14][19] * mat_B[19][19] +
                  mat_A[14][20] * mat_B[20][19] +
                  mat_A[14][21] * mat_B[21][19] +
                  mat_A[14][22] * mat_B[22][19] +
                  mat_A[14][23] * mat_B[23][19] +
                  mat_A[14][24] * mat_B[24][19] +
                  mat_A[14][25] * mat_B[25][19] +
                  mat_A[14][26] * mat_B[26][19] +
                  mat_A[14][27] * mat_B[27][19] +
                  mat_A[14][28] * mat_B[28][19] +
                  mat_A[14][29] * mat_B[29][19] +
                  mat_A[14][30] * mat_B[30][19] +
                  mat_A[14][31] * mat_B[31][19];
    mat_C[14][20] <= 
                  mat_A[14][0] * mat_B[0][20] +
                  mat_A[14][1] * mat_B[1][20] +
                  mat_A[14][2] * mat_B[2][20] +
                  mat_A[14][3] * mat_B[3][20] +
                  mat_A[14][4] * mat_B[4][20] +
                  mat_A[14][5] * mat_B[5][20] +
                  mat_A[14][6] * mat_B[6][20] +
                  mat_A[14][7] * mat_B[7][20] +
                  mat_A[14][8] * mat_B[8][20] +
                  mat_A[14][9] * mat_B[9][20] +
                  mat_A[14][10] * mat_B[10][20] +
                  mat_A[14][11] * mat_B[11][20] +
                  mat_A[14][12] * mat_B[12][20] +
                  mat_A[14][13] * mat_B[13][20] +
                  mat_A[14][14] * mat_B[14][20] +
                  mat_A[14][15] * mat_B[15][20] +
                  mat_A[14][16] * mat_B[16][20] +
                  mat_A[14][17] * mat_B[17][20] +
                  mat_A[14][18] * mat_B[18][20] +
                  mat_A[14][19] * mat_B[19][20] +
                  mat_A[14][20] * mat_B[20][20] +
                  mat_A[14][21] * mat_B[21][20] +
                  mat_A[14][22] * mat_B[22][20] +
                  mat_A[14][23] * mat_B[23][20] +
                  mat_A[14][24] * mat_B[24][20] +
                  mat_A[14][25] * mat_B[25][20] +
                  mat_A[14][26] * mat_B[26][20] +
                  mat_A[14][27] * mat_B[27][20] +
                  mat_A[14][28] * mat_B[28][20] +
                  mat_A[14][29] * mat_B[29][20] +
                  mat_A[14][30] * mat_B[30][20] +
                  mat_A[14][31] * mat_B[31][20];
    mat_C[14][21] <= 
                  mat_A[14][0] * mat_B[0][21] +
                  mat_A[14][1] * mat_B[1][21] +
                  mat_A[14][2] * mat_B[2][21] +
                  mat_A[14][3] * mat_B[3][21] +
                  mat_A[14][4] * mat_B[4][21] +
                  mat_A[14][5] * mat_B[5][21] +
                  mat_A[14][6] * mat_B[6][21] +
                  mat_A[14][7] * mat_B[7][21] +
                  mat_A[14][8] * mat_B[8][21] +
                  mat_A[14][9] * mat_B[9][21] +
                  mat_A[14][10] * mat_B[10][21] +
                  mat_A[14][11] * mat_B[11][21] +
                  mat_A[14][12] * mat_B[12][21] +
                  mat_A[14][13] * mat_B[13][21] +
                  mat_A[14][14] * mat_B[14][21] +
                  mat_A[14][15] * mat_B[15][21] +
                  mat_A[14][16] * mat_B[16][21] +
                  mat_A[14][17] * mat_B[17][21] +
                  mat_A[14][18] * mat_B[18][21] +
                  mat_A[14][19] * mat_B[19][21] +
                  mat_A[14][20] * mat_B[20][21] +
                  mat_A[14][21] * mat_B[21][21] +
                  mat_A[14][22] * mat_B[22][21] +
                  mat_A[14][23] * mat_B[23][21] +
                  mat_A[14][24] * mat_B[24][21] +
                  mat_A[14][25] * mat_B[25][21] +
                  mat_A[14][26] * mat_B[26][21] +
                  mat_A[14][27] * mat_B[27][21] +
                  mat_A[14][28] * mat_B[28][21] +
                  mat_A[14][29] * mat_B[29][21] +
                  mat_A[14][30] * mat_B[30][21] +
                  mat_A[14][31] * mat_B[31][21];
    mat_C[14][22] <= 
                  mat_A[14][0] * mat_B[0][22] +
                  mat_A[14][1] * mat_B[1][22] +
                  mat_A[14][2] * mat_B[2][22] +
                  mat_A[14][3] * mat_B[3][22] +
                  mat_A[14][4] * mat_B[4][22] +
                  mat_A[14][5] * mat_B[5][22] +
                  mat_A[14][6] * mat_B[6][22] +
                  mat_A[14][7] * mat_B[7][22] +
                  mat_A[14][8] * mat_B[8][22] +
                  mat_A[14][9] * mat_B[9][22] +
                  mat_A[14][10] * mat_B[10][22] +
                  mat_A[14][11] * mat_B[11][22] +
                  mat_A[14][12] * mat_B[12][22] +
                  mat_A[14][13] * mat_B[13][22] +
                  mat_A[14][14] * mat_B[14][22] +
                  mat_A[14][15] * mat_B[15][22] +
                  mat_A[14][16] * mat_B[16][22] +
                  mat_A[14][17] * mat_B[17][22] +
                  mat_A[14][18] * mat_B[18][22] +
                  mat_A[14][19] * mat_B[19][22] +
                  mat_A[14][20] * mat_B[20][22] +
                  mat_A[14][21] * mat_B[21][22] +
                  mat_A[14][22] * mat_B[22][22] +
                  mat_A[14][23] * mat_B[23][22] +
                  mat_A[14][24] * mat_B[24][22] +
                  mat_A[14][25] * mat_B[25][22] +
                  mat_A[14][26] * mat_B[26][22] +
                  mat_A[14][27] * mat_B[27][22] +
                  mat_A[14][28] * mat_B[28][22] +
                  mat_A[14][29] * mat_B[29][22] +
                  mat_A[14][30] * mat_B[30][22] +
                  mat_A[14][31] * mat_B[31][22];
    mat_C[14][23] <= 
                  mat_A[14][0] * mat_B[0][23] +
                  mat_A[14][1] * mat_B[1][23] +
                  mat_A[14][2] * mat_B[2][23] +
                  mat_A[14][3] * mat_B[3][23] +
                  mat_A[14][4] * mat_B[4][23] +
                  mat_A[14][5] * mat_B[5][23] +
                  mat_A[14][6] * mat_B[6][23] +
                  mat_A[14][7] * mat_B[7][23] +
                  mat_A[14][8] * mat_B[8][23] +
                  mat_A[14][9] * mat_B[9][23] +
                  mat_A[14][10] * mat_B[10][23] +
                  mat_A[14][11] * mat_B[11][23] +
                  mat_A[14][12] * mat_B[12][23] +
                  mat_A[14][13] * mat_B[13][23] +
                  mat_A[14][14] * mat_B[14][23] +
                  mat_A[14][15] * mat_B[15][23] +
                  mat_A[14][16] * mat_B[16][23] +
                  mat_A[14][17] * mat_B[17][23] +
                  mat_A[14][18] * mat_B[18][23] +
                  mat_A[14][19] * mat_B[19][23] +
                  mat_A[14][20] * mat_B[20][23] +
                  mat_A[14][21] * mat_B[21][23] +
                  mat_A[14][22] * mat_B[22][23] +
                  mat_A[14][23] * mat_B[23][23] +
                  mat_A[14][24] * mat_B[24][23] +
                  mat_A[14][25] * mat_B[25][23] +
                  mat_A[14][26] * mat_B[26][23] +
                  mat_A[14][27] * mat_B[27][23] +
                  mat_A[14][28] * mat_B[28][23] +
                  mat_A[14][29] * mat_B[29][23] +
                  mat_A[14][30] * mat_B[30][23] +
                  mat_A[14][31] * mat_B[31][23];
    mat_C[14][24] <= 
                  mat_A[14][0] * mat_B[0][24] +
                  mat_A[14][1] * mat_B[1][24] +
                  mat_A[14][2] * mat_B[2][24] +
                  mat_A[14][3] * mat_B[3][24] +
                  mat_A[14][4] * mat_B[4][24] +
                  mat_A[14][5] * mat_B[5][24] +
                  mat_A[14][6] * mat_B[6][24] +
                  mat_A[14][7] * mat_B[7][24] +
                  mat_A[14][8] * mat_B[8][24] +
                  mat_A[14][9] * mat_B[9][24] +
                  mat_A[14][10] * mat_B[10][24] +
                  mat_A[14][11] * mat_B[11][24] +
                  mat_A[14][12] * mat_B[12][24] +
                  mat_A[14][13] * mat_B[13][24] +
                  mat_A[14][14] * mat_B[14][24] +
                  mat_A[14][15] * mat_B[15][24] +
                  mat_A[14][16] * mat_B[16][24] +
                  mat_A[14][17] * mat_B[17][24] +
                  mat_A[14][18] * mat_B[18][24] +
                  mat_A[14][19] * mat_B[19][24] +
                  mat_A[14][20] * mat_B[20][24] +
                  mat_A[14][21] * mat_B[21][24] +
                  mat_A[14][22] * mat_B[22][24] +
                  mat_A[14][23] * mat_B[23][24] +
                  mat_A[14][24] * mat_B[24][24] +
                  mat_A[14][25] * mat_B[25][24] +
                  mat_A[14][26] * mat_B[26][24] +
                  mat_A[14][27] * mat_B[27][24] +
                  mat_A[14][28] * mat_B[28][24] +
                  mat_A[14][29] * mat_B[29][24] +
                  mat_A[14][30] * mat_B[30][24] +
                  mat_A[14][31] * mat_B[31][24];
    mat_C[14][25] <= 
                  mat_A[14][0] * mat_B[0][25] +
                  mat_A[14][1] * mat_B[1][25] +
                  mat_A[14][2] * mat_B[2][25] +
                  mat_A[14][3] * mat_B[3][25] +
                  mat_A[14][4] * mat_B[4][25] +
                  mat_A[14][5] * mat_B[5][25] +
                  mat_A[14][6] * mat_B[6][25] +
                  mat_A[14][7] * mat_B[7][25] +
                  mat_A[14][8] * mat_B[8][25] +
                  mat_A[14][9] * mat_B[9][25] +
                  mat_A[14][10] * mat_B[10][25] +
                  mat_A[14][11] * mat_B[11][25] +
                  mat_A[14][12] * mat_B[12][25] +
                  mat_A[14][13] * mat_B[13][25] +
                  mat_A[14][14] * mat_B[14][25] +
                  mat_A[14][15] * mat_B[15][25] +
                  mat_A[14][16] * mat_B[16][25] +
                  mat_A[14][17] * mat_B[17][25] +
                  mat_A[14][18] * mat_B[18][25] +
                  mat_A[14][19] * mat_B[19][25] +
                  mat_A[14][20] * mat_B[20][25] +
                  mat_A[14][21] * mat_B[21][25] +
                  mat_A[14][22] * mat_B[22][25] +
                  mat_A[14][23] * mat_B[23][25] +
                  mat_A[14][24] * mat_B[24][25] +
                  mat_A[14][25] * mat_B[25][25] +
                  mat_A[14][26] * mat_B[26][25] +
                  mat_A[14][27] * mat_B[27][25] +
                  mat_A[14][28] * mat_B[28][25] +
                  mat_A[14][29] * mat_B[29][25] +
                  mat_A[14][30] * mat_B[30][25] +
                  mat_A[14][31] * mat_B[31][25];
    mat_C[14][26] <= 
                  mat_A[14][0] * mat_B[0][26] +
                  mat_A[14][1] * mat_B[1][26] +
                  mat_A[14][2] * mat_B[2][26] +
                  mat_A[14][3] * mat_B[3][26] +
                  mat_A[14][4] * mat_B[4][26] +
                  mat_A[14][5] * mat_B[5][26] +
                  mat_A[14][6] * mat_B[6][26] +
                  mat_A[14][7] * mat_B[7][26] +
                  mat_A[14][8] * mat_B[8][26] +
                  mat_A[14][9] * mat_B[9][26] +
                  mat_A[14][10] * mat_B[10][26] +
                  mat_A[14][11] * mat_B[11][26] +
                  mat_A[14][12] * mat_B[12][26] +
                  mat_A[14][13] * mat_B[13][26] +
                  mat_A[14][14] * mat_B[14][26] +
                  mat_A[14][15] * mat_B[15][26] +
                  mat_A[14][16] * mat_B[16][26] +
                  mat_A[14][17] * mat_B[17][26] +
                  mat_A[14][18] * mat_B[18][26] +
                  mat_A[14][19] * mat_B[19][26] +
                  mat_A[14][20] * mat_B[20][26] +
                  mat_A[14][21] * mat_B[21][26] +
                  mat_A[14][22] * mat_B[22][26] +
                  mat_A[14][23] * mat_B[23][26] +
                  mat_A[14][24] * mat_B[24][26] +
                  mat_A[14][25] * mat_B[25][26] +
                  mat_A[14][26] * mat_B[26][26] +
                  mat_A[14][27] * mat_B[27][26] +
                  mat_A[14][28] * mat_B[28][26] +
                  mat_A[14][29] * mat_B[29][26] +
                  mat_A[14][30] * mat_B[30][26] +
                  mat_A[14][31] * mat_B[31][26];
    mat_C[14][27] <= 
                  mat_A[14][0] * mat_B[0][27] +
                  mat_A[14][1] * mat_B[1][27] +
                  mat_A[14][2] * mat_B[2][27] +
                  mat_A[14][3] * mat_B[3][27] +
                  mat_A[14][4] * mat_B[4][27] +
                  mat_A[14][5] * mat_B[5][27] +
                  mat_A[14][6] * mat_B[6][27] +
                  mat_A[14][7] * mat_B[7][27] +
                  mat_A[14][8] * mat_B[8][27] +
                  mat_A[14][9] * mat_B[9][27] +
                  mat_A[14][10] * mat_B[10][27] +
                  mat_A[14][11] * mat_B[11][27] +
                  mat_A[14][12] * mat_B[12][27] +
                  mat_A[14][13] * mat_B[13][27] +
                  mat_A[14][14] * mat_B[14][27] +
                  mat_A[14][15] * mat_B[15][27] +
                  mat_A[14][16] * mat_B[16][27] +
                  mat_A[14][17] * mat_B[17][27] +
                  mat_A[14][18] * mat_B[18][27] +
                  mat_A[14][19] * mat_B[19][27] +
                  mat_A[14][20] * mat_B[20][27] +
                  mat_A[14][21] * mat_B[21][27] +
                  mat_A[14][22] * mat_B[22][27] +
                  mat_A[14][23] * mat_B[23][27] +
                  mat_A[14][24] * mat_B[24][27] +
                  mat_A[14][25] * mat_B[25][27] +
                  mat_A[14][26] * mat_B[26][27] +
                  mat_A[14][27] * mat_B[27][27] +
                  mat_A[14][28] * mat_B[28][27] +
                  mat_A[14][29] * mat_B[29][27] +
                  mat_A[14][30] * mat_B[30][27] +
                  mat_A[14][31] * mat_B[31][27];
    mat_C[14][28] <= 
                  mat_A[14][0] * mat_B[0][28] +
                  mat_A[14][1] * mat_B[1][28] +
                  mat_A[14][2] * mat_B[2][28] +
                  mat_A[14][3] * mat_B[3][28] +
                  mat_A[14][4] * mat_B[4][28] +
                  mat_A[14][5] * mat_B[5][28] +
                  mat_A[14][6] * mat_B[6][28] +
                  mat_A[14][7] * mat_B[7][28] +
                  mat_A[14][8] * mat_B[8][28] +
                  mat_A[14][9] * mat_B[9][28] +
                  mat_A[14][10] * mat_B[10][28] +
                  mat_A[14][11] * mat_B[11][28] +
                  mat_A[14][12] * mat_B[12][28] +
                  mat_A[14][13] * mat_B[13][28] +
                  mat_A[14][14] * mat_B[14][28] +
                  mat_A[14][15] * mat_B[15][28] +
                  mat_A[14][16] * mat_B[16][28] +
                  mat_A[14][17] * mat_B[17][28] +
                  mat_A[14][18] * mat_B[18][28] +
                  mat_A[14][19] * mat_B[19][28] +
                  mat_A[14][20] * mat_B[20][28] +
                  mat_A[14][21] * mat_B[21][28] +
                  mat_A[14][22] * mat_B[22][28] +
                  mat_A[14][23] * mat_B[23][28] +
                  mat_A[14][24] * mat_B[24][28] +
                  mat_A[14][25] * mat_B[25][28] +
                  mat_A[14][26] * mat_B[26][28] +
                  mat_A[14][27] * mat_B[27][28] +
                  mat_A[14][28] * mat_B[28][28] +
                  mat_A[14][29] * mat_B[29][28] +
                  mat_A[14][30] * mat_B[30][28] +
                  mat_A[14][31] * mat_B[31][28];
    mat_C[14][29] <= 
                  mat_A[14][0] * mat_B[0][29] +
                  mat_A[14][1] * mat_B[1][29] +
                  mat_A[14][2] * mat_B[2][29] +
                  mat_A[14][3] * mat_B[3][29] +
                  mat_A[14][4] * mat_B[4][29] +
                  mat_A[14][5] * mat_B[5][29] +
                  mat_A[14][6] * mat_B[6][29] +
                  mat_A[14][7] * mat_B[7][29] +
                  mat_A[14][8] * mat_B[8][29] +
                  mat_A[14][9] * mat_B[9][29] +
                  mat_A[14][10] * mat_B[10][29] +
                  mat_A[14][11] * mat_B[11][29] +
                  mat_A[14][12] * mat_B[12][29] +
                  mat_A[14][13] * mat_B[13][29] +
                  mat_A[14][14] * mat_B[14][29] +
                  mat_A[14][15] * mat_B[15][29] +
                  mat_A[14][16] * mat_B[16][29] +
                  mat_A[14][17] * mat_B[17][29] +
                  mat_A[14][18] * mat_B[18][29] +
                  mat_A[14][19] * mat_B[19][29] +
                  mat_A[14][20] * mat_B[20][29] +
                  mat_A[14][21] * mat_B[21][29] +
                  mat_A[14][22] * mat_B[22][29] +
                  mat_A[14][23] * mat_B[23][29] +
                  mat_A[14][24] * mat_B[24][29] +
                  mat_A[14][25] * mat_B[25][29] +
                  mat_A[14][26] * mat_B[26][29] +
                  mat_A[14][27] * mat_B[27][29] +
                  mat_A[14][28] * mat_B[28][29] +
                  mat_A[14][29] * mat_B[29][29] +
                  mat_A[14][30] * mat_B[30][29] +
                  mat_A[14][31] * mat_B[31][29];
    mat_C[14][30] <= 
                  mat_A[14][0] * mat_B[0][30] +
                  mat_A[14][1] * mat_B[1][30] +
                  mat_A[14][2] * mat_B[2][30] +
                  mat_A[14][3] * mat_B[3][30] +
                  mat_A[14][4] * mat_B[4][30] +
                  mat_A[14][5] * mat_B[5][30] +
                  mat_A[14][6] * mat_B[6][30] +
                  mat_A[14][7] * mat_B[7][30] +
                  mat_A[14][8] * mat_B[8][30] +
                  mat_A[14][9] * mat_B[9][30] +
                  mat_A[14][10] * mat_B[10][30] +
                  mat_A[14][11] * mat_B[11][30] +
                  mat_A[14][12] * mat_B[12][30] +
                  mat_A[14][13] * mat_B[13][30] +
                  mat_A[14][14] * mat_B[14][30] +
                  mat_A[14][15] * mat_B[15][30] +
                  mat_A[14][16] * mat_B[16][30] +
                  mat_A[14][17] * mat_B[17][30] +
                  mat_A[14][18] * mat_B[18][30] +
                  mat_A[14][19] * mat_B[19][30] +
                  mat_A[14][20] * mat_B[20][30] +
                  mat_A[14][21] * mat_B[21][30] +
                  mat_A[14][22] * mat_B[22][30] +
                  mat_A[14][23] * mat_B[23][30] +
                  mat_A[14][24] * mat_B[24][30] +
                  mat_A[14][25] * mat_B[25][30] +
                  mat_A[14][26] * mat_B[26][30] +
                  mat_A[14][27] * mat_B[27][30] +
                  mat_A[14][28] * mat_B[28][30] +
                  mat_A[14][29] * mat_B[29][30] +
                  mat_A[14][30] * mat_B[30][30] +
                  mat_A[14][31] * mat_B[31][30];
    mat_C[14][31] <= 
                  mat_A[14][0] * mat_B[0][31] +
                  mat_A[14][1] * mat_B[1][31] +
                  mat_A[14][2] * mat_B[2][31] +
                  mat_A[14][3] * mat_B[3][31] +
                  mat_A[14][4] * mat_B[4][31] +
                  mat_A[14][5] * mat_B[5][31] +
                  mat_A[14][6] * mat_B[6][31] +
                  mat_A[14][7] * mat_B[7][31] +
                  mat_A[14][8] * mat_B[8][31] +
                  mat_A[14][9] * mat_B[9][31] +
                  mat_A[14][10] * mat_B[10][31] +
                  mat_A[14][11] * mat_B[11][31] +
                  mat_A[14][12] * mat_B[12][31] +
                  mat_A[14][13] * mat_B[13][31] +
                  mat_A[14][14] * mat_B[14][31] +
                  mat_A[14][15] * mat_B[15][31] +
                  mat_A[14][16] * mat_B[16][31] +
                  mat_A[14][17] * mat_B[17][31] +
                  mat_A[14][18] * mat_B[18][31] +
                  mat_A[14][19] * mat_B[19][31] +
                  mat_A[14][20] * mat_B[20][31] +
                  mat_A[14][21] * mat_B[21][31] +
                  mat_A[14][22] * mat_B[22][31] +
                  mat_A[14][23] * mat_B[23][31] +
                  mat_A[14][24] * mat_B[24][31] +
                  mat_A[14][25] * mat_B[25][31] +
                  mat_A[14][26] * mat_B[26][31] +
                  mat_A[14][27] * mat_B[27][31] +
                  mat_A[14][28] * mat_B[28][31] +
                  mat_A[14][29] * mat_B[29][31] +
                  mat_A[14][30] * mat_B[30][31] +
                  mat_A[14][31] * mat_B[31][31];
    mat_C[15][0] <= 
                  mat_A[15][0] * mat_B[0][0] +
                  mat_A[15][1] * mat_B[1][0] +
                  mat_A[15][2] * mat_B[2][0] +
                  mat_A[15][3] * mat_B[3][0] +
                  mat_A[15][4] * mat_B[4][0] +
                  mat_A[15][5] * mat_B[5][0] +
                  mat_A[15][6] * mat_B[6][0] +
                  mat_A[15][7] * mat_B[7][0] +
                  mat_A[15][8] * mat_B[8][0] +
                  mat_A[15][9] * mat_B[9][0] +
                  mat_A[15][10] * mat_B[10][0] +
                  mat_A[15][11] * mat_B[11][0] +
                  mat_A[15][12] * mat_B[12][0] +
                  mat_A[15][13] * mat_B[13][0] +
                  mat_A[15][14] * mat_B[14][0] +
                  mat_A[15][15] * mat_B[15][0] +
                  mat_A[15][16] * mat_B[16][0] +
                  mat_A[15][17] * mat_B[17][0] +
                  mat_A[15][18] * mat_B[18][0] +
                  mat_A[15][19] * mat_B[19][0] +
                  mat_A[15][20] * mat_B[20][0] +
                  mat_A[15][21] * mat_B[21][0] +
                  mat_A[15][22] * mat_B[22][0] +
                  mat_A[15][23] * mat_B[23][0] +
                  mat_A[15][24] * mat_B[24][0] +
                  mat_A[15][25] * mat_B[25][0] +
                  mat_A[15][26] * mat_B[26][0] +
                  mat_A[15][27] * mat_B[27][0] +
                  mat_A[15][28] * mat_B[28][0] +
                  mat_A[15][29] * mat_B[29][0] +
                  mat_A[15][30] * mat_B[30][0] +
                  mat_A[15][31] * mat_B[31][0];
    mat_C[15][1] <= 
                  mat_A[15][0] * mat_B[0][1] +
                  mat_A[15][1] * mat_B[1][1] +
                  mat_A[15][2] * mat_B[2][1] +
                  mat_A[15][3] * mat_B[3][1] +
                  mat_A[15][4] * mat_B[4][1] +
                  mat_A[15][5] * mat_B[5][1] +
                  mat_A[15][6] * mat_B[6][1] +
                  mat_A[15][7] * mat_B[7][1] +
                  mat_A[15][8] * mat_B[8][1] +
                  mat_A[15][9] * mat_B[9][1] +
                  mat_A[15][10] * mat_B[10][1] +
                  mat_A[15][11] * mat_B[11][1] +
                  mat_A[15][12] * mat_B[12][1] +
                  mat_A[15][13] * mat_B[13][1] +
                  mat_A[15][14] * mat_B[14][1] +
                  mat_A[15][15] * mat_B[15][1] +
                  mat_A[15][16] * mat_B[16][1] +
                  mat_A[15][17] * mat_B[17][1] +
                  mat_A[15][18] * mat_B[18][1] +
                  mat_A[15][19] * mat_B[19][1] +
                  mat_A[15][20] * mat_B[20][1] +
                  mat_A[15][21] * mat_B[21][1] +
                  mat_A[15][22] * mat_B[22][1] +
                  mat_A[15][23] * mat_B[23][1] +
                  mat_A[15][24] * mat_B[24][1] +
                  mat_A[15][25] * mat_B[25][1] +
                  mat_A[15][26] * mat_B[26][1] +
                  mat_A[15][27] * mat_B[27][1] +
                  mat_A[15][28] * mat_B[28][1] +
                  mat_A[15][29] * mat_B[29][1] +
                  mat_A[15][30] * mat_B[30][1] +
                  mat_A[15][31] * mat_B[31][1];
    mat_C[15][2] <= 
                  mat_A[15][0] * mat_B[0][2] +
                  mat_A[15][1] * mat_B[1][2] +
                  mat_A[15][2] * mat_B[2][2] +
                  mat_A[15][3] * mat_B[3][2] +
                  mat_A[15][4] * mat_B[4][2] +
                  mat_A[15][5] * mat_B[5][2] +
                  mat_A[15][6] * mat_B[6][2] +
                  mat_A[15][7] * mat_B[7][2] +
                  mat_A[15][8] * mat_B[8][2] +
                  mat_A[15][9] * mat_B[9][2] +
                  mat_A[15][10] * mat_B[10][2] +
                  mat_A[15][11] * mat_B[11][2] +
                  mat_A[15][12] * mat_B[12][2] +
                  mat_A[15][13] * mat_B[13][2] +
                  mat_A[15][14] * mat_B[14][2] +
                  mat_A[15][15] * mat_B[15][2] +
                  mat_A[15][16] * mat_B[16][2] +
                  mat_A[15][17] * mat_B[17][2] +
                  mat_A[15][18] * mat_B[18][2] +
                  mat_A[15][19] * mat_B[19][2] +
                  mat_A[15][20] * mat_B[20][2] +
                  mat_A[15][21] * mat_B[21][2] +
                  mat_A[15][22] * mat_B[22][2] +
                  mat_A[15][23] * mat_B[23][2] +
                  mat_A[15][24] * mat_B[24][2] +
                  mat_A[15][25] * mat_B[25][2] +
                  mat_A[15][26] * mat_B[26][2] +
                  mat_A[15][27] * mat_B[27][2] +
                  mat_A[15][28] * mat_B[28][2] +
                  mat_A[15][29] * mat_B[29][2] +
                  mat_A[15][30] * mat_B[30][2] +
                  mat_A[15][31] * mat_B[31][2];
    mat_C[15][3] <= 
                  mat_A[15][0] * mat_B[0][3] +
                  mat_A[15][1] * mat_B[1][3] +
                  mat_A[15][2] * mat_B[2][3] +
                  mat_A[15][3] * mat_B[3][3] +
                  mat_A[15][4] * mat_B[4][3] +
                  mat_A[15][5] * mat_B[5][3] +
                  mat_A[15][6] * mat_B[6][3] +
                  mat_A[15][7] * mat_B[7][3] +
                  mat_A[15][8] * mat_B[8][3] +
                  mat_A[15][9] * mat_B[9][3] +
                  mat_A[15][10] * mat_B[10][3] +
                  mat_A[15][11] * mat_B[11][3] +
                  mat_A[15][12] * mat_B[12][3] +
                  mat_A[15][13] * mat_B[13][3] +
                  mat_A[15][14] * mat_B[14][3] +
                  mat_A[15][15] * mat_B[15][3] +
                  mat_A[15][16] * mat_B[16][3] +
                  mat_A[15][17] * mat_B[17][3] +
                  mat_A[15][18] * mat_B[18][3] +
                  mat_A[15][19] * mat_B[19][3] +
                  mat_A[15][20] * mat_B[20][3] +
                  mat_A[15][21] * mat_B[21][3] +
                  mat_A[15][22] * mat_B[22][3] +
                  mat_A[15][23] * mat_B[23][3] +
                  mat_A[15][24] * mat_B[24][3] +
                  mat_A[15][25] * mat_B[25][3] +
                  mat_A[15][26] * mat_B[26][3] +
                  mat_A[15][27] * mat_B[27][3] +
                  mat_A[15][28] * mat_B[28][3] +
                  mat_A[15][29] * mat_B[29][3] +
                  mat_A[15][30] * mat_B[30][3] +
                  mat_A[15][31] * mat_B[31][3];
    mat_C[15][4] <= 
                  mat_A[15][0] * mat_B[0][4] +
                  mat_A[15][1] * mat_B[1][4] +
                  mat_A[15][2] * mat_B[2][4] +
                  mat_A[15][3] * mat_B[3][4] +
                  mat_A[15][4] * mat_B[4][4] +
                  mat_A[15][5] * mat_B[5][4] +
                  mat_A[15][6] * mat_B[6][4] +
                  mat_A[15][7] * mat_B[7][4] +
                  mat_A[15][8] * mat_B[8][4] +
                  mat_A[15][9] * mat_B[9][4] +
                  mat_A[15][10] * mat_B[10][4] +
                  mat_A[15][11] * mat_B[11][4] +
                  mat_A[15][12] * mat_B[12][4] +
                  mat_A[15][13] * mat_B[13][4] +
                  mat_A[15][14] * mat_B[14][4] +
                  mat_A[15][15] * mat_B[15][4] +
                  mat_A[15][16] * mat_B[16][4] +
                  mat_A[15][17] * mat_B[17][4] +
                  mat_A[15][18] * mat_B[18][4] +
                  mat_A[15][19] * mat_B[19][4] +
                  mat_A[15][20] * mat_B[20][4] +
                  mat_A[15][21] * mat_B[21][4] +
                  mat_A[15][22] * mat_B[22][4] +
                  mat_A[15][23] * mat_B[23][4] +
                  mat_A[15][24] * mat_B[24][4] +
                  mat_A[15][25] * mat_B[25][4] +
                  mat_A[15][26] * mat_B[26][4] +
                  mat_A[15][27] * mat_B[27][4] +
                  mat_A[15][28] * mat_B[28][4] +
                  mat_A[15][29] * mat_B[29][4] +
                  mat_A[15][30] * mat_B[30][4] +
                  mat_A[15][31] * mat_B[31][4];
    mat_C[15][5] <= 
                  mat_A[15][0] * mat_B[0][5] +
                  mat_A[15][1] * mat_B[1][5] +
                  mat_A[15][2] * mat_B[2][5] +
                  mat_A[15][3] * mat_B[3][5] +
                  mat_A[15][4] * mat_B[4][5] +
                  mat_A[15][5] * mat_B[5][5] +
                  mat_A[15][6] * mat_B[6][5] +
                  mat_A[15][7] * mat_B[7][5] +
                  mat_A[15][8] * mat_B[8][5] +
                  mat_A[15][9] * mat_B[9][5] +
                  mat_A[15][10] * mat_B[10][5] +
                  mat_A[15][11] * mat_B[11][5] +
                  mat_A[15][12] * mat_B[12][5] +
                  mat_A[15][13] * mat_B[13][5] +
                  mat_A[15][14] * mat_B[14][5] +
                  mat_A[15][15] * mat_B[15][5] +
                  mat_A[15][16] * mat_B[16][5] +
                  mat_A[15][17] * mat_B[17][5] +
                  mat_A[15][18] * mat_B[18][5] +
                  mat_A[15][19] * mat_B[19][5] +
                  mat_A[15][20] * mat_B[20][5] +
                  mat_A[15][21] * mat_B[21][5] +
                  mat_A[15][22] * mat_B[22][5] +
                  mat_A[15][23] * mat_B[23][5] +
                  mat_A[15][24] * mat_B[24][5] +
                  mat_A[15][25] * mat_B[25][5] +
                  mat_A[15][26] * mat_B[26][5] +
                  mat_A[15][27] * mat_B[27][5] +
                  mat_A[15][28] * mat_B[28][5] +
                  mat_A[15][29] * mat_B[29][5] +
                  mat_A[15][30] * mat_B[30][5] +
                  mat_A[15][31] * mat_B[31][5];
    mat_C[15][6] <= 
                  mat_A[15][0] * mat_B[0][6] +
                  mat_A[15][1] * mat_B[1][6] +
                  mat_A[15][2] * mat_B[2][6] +
                  mat_A[15][3] * mat_B[3][6] +
                  mat_A[15][4] * mat_B[4][6] +
                  mat_A[15][5] * mat_B[5][6] +
                  mat_A[15][6] * mat_B[6][6] +
                  mat_A[15][7] * mat_B[7][6] +
                  mat_A[15][8] * mat_B[8][6] +
                  mat_A[15][9] * mat_B[9][6] +
                  mat_A[15][10] * mat_B[10][6] +
                  mat_A[15][11] * mat_B[11][6] +
                  mat_A[15][12] * mat_B[12][6] +
                  mat_A[15][13] * mat_B[13][6] +
                  mat_A[15][14] * mat_B[14][6] +
                  mat_A[15][15] * mat_B[15][6] +
                  mat_A[15][16] * mat_B[16][6] +
                  mat_A[15][17] * mat_B[17][6] +
                  mat_A[15][18] * mat_B[18][6] +
                  mat_A[15][19] * mat_B[19][6] +
                  mat_A[15][20] * mat_B[20][6] +
                  mat_A[15][21] * mat_B[21][6] +
                  mat_A[15][22] * mat_B[22][6] +
                  mat_A[15][23] * mat_B[23][6] +
                  mat_A[15][24] * mat_B[24][6] +
                  mat_A[15][25] * mat_B[25][6] +
                  mat_A[15][26] * mat_B[26][6] +
                  mat_A[15][27] * mat_B[27][6] +
                  mat_A[15][28] * mat_B[28][6] +
                  mat_A[15][29] * mat_B[29][6] +
                  mat_A[15][30] * mat_B[30][6] +
                  mat_A[15][31] * mat_B[31][6];
    mat_C[15][7] <= 
                  mat_A[15][0] * mat_B[0][7] +
                  mat_A[15][1] * mat_B[1][7] +
                  mat_A[15][2] * mat_B[2][7] +
                  mat_A[15][3] * mat_B[3][7] +
                  mat_A[15][4] * mat_B[4][7] +
                  mat_A[15][5] * mat_B[5][7] +
                  mat_A[15][6] * mat_B[6][7] +
                  mat_A[15][7] * mat_B[7][7] +
                  mat_A[15][8] * mat_B[8][7] +
                  mat_A[15][9] * mat_B[9][7] +
                  mat_A[15][10] * mat_B[10][7] +
                  mat_A[15][11] * mat_B[11][7] +
                  mat_A[15][12] * mat_B[12][7] +
                  mat_A[15][13] * mat_B[13][7] +
                  mat_A[15][14] * mat_B[14][7] +
                  mat_A[15][15] * mat_B[15][7] +
                  mat_A[15][16] * mat_B[16][7] +
                  mat_A[15][17] * mat_B[17][7] +
                  mat_A[15][18] * mat_B[18][7] +
                  mat_A[15][19] * mat_B[19][7] +
                  mat_A[15][20] * mat_B[20][7] +
                  mat_A[15][21] * mat_B[21][7] +
                  mat_A[15][22] * mat_B[22][7] +
                  mat_A[15][23] * mat_B[23][7] +
                  mat_A[15][24] * mat_B[24][7] +
                  mat_A[15][25] * mat_B[25][7] +
                  mat_A[15][26] * mat_B[26][7] +
                  mat_A[15][27] * mat_B[27][7] +
                  mat_A[15][28] * mat_B[28][7] +
                  mat_A[15][29] * mat_B[29][7] +
                  mat_A[15][30] * mat_B[30][7] +
                  mat_A[15][31] * mat_B[31][7];
    mat_C[15][8] <= 
                  mat_A[15][0] * mat_B[0][8] +
                  mat_A[15][1] * mat_B[1][8] +
                  mat_A[15][2] * mat_B[2][8] +
                  mat_A[15][3] * mat_B[3][8] +
                  mat_A[15][4] * mat_B[4][8] +
                  mat_A[15][5] * mat_B[5][8] +
                  mat_A[15][6] * mat_B[6][8] +
                  mat_A[15][7] * mat_B[7][8] +
                  mat_A[15][8] * mat_B[8][8] +
                  mat_A[15][9] * mat_B[9][8] +
                  mat_A[15][10] * mat_B[10][8] +
                  mat_A[15][11] * mat_B[11][8] +
                  mat_A[15][12] * mat_B[12][8] +
                  mat_A[15][13] * mat_B[13][8] +
                  mat_A[15][14] * mat_B[14][8] +
                  mat_A[15][15] * mat_B[15][8] +
                  mat_A[15][16] * mat_B[16][8] +
                  mat_A[15][17] * mat_B[17][8] +
                  mat_A[15][18] * mat_B[18][8] +
                  mat_A[15][19] * mat_B[19][8] +
                  mat_A[15][20] * mat_B[20][8] +
                  mat_A[15][21] * mat_B[21][8] +
                  mat_A[15][22] * mat_B[22][8] +
                  mat_A[15][23] * mat_B[23][8] +
                  mat_A[15][24] * mat_B[24][8] +
                  mat_A[15][25] * mat_B[25][8] +
                  mat_A[15][26] * mat_B[26][8] +
                  mat_A[15][27] * mat_B[27][8] +
                  mat_A[15][28] * mat_B[28][8] +
                  mat_A[15][29] * mat_B[29][8] +
                  mat_A[15][30] * mat_B[30][8] +
                  mat_A[15][31] * mat_B[31][8];
    mat_C[15][9] <= 
                  mat_A[15][0] * mat_B[0][9] +
                  mat_A[15][1] * mat_B[1][9] +
                  mat_A[15][2] * mat_B[2][9] +
                  mat_A[15][3] * mat_B[3][9] +
                  mat_A[15][4] * mat_B[4][9] +
                  mat_A[15][5] * mat_B[5][9] +
                  mat_A[15][6] * mat_B[6][9] +
                  mat_A[15][7] * mat_B[7][9] +
                  mat_A[15][8] * mat_B[8][9] +
                  mat_A[15][9] * mat_B[9][9] +
                  mat_A[15][10] * mat_B[10][9] +
                  mat_A[15][11] * mat_B[11][9] +
                  mat_A[15][12] * mat_B[12][9] +
                  mat_A[15][13] * mat_B[13][9] +
                  mat_A[15][14] * mat_B[14][9] +
                  mat_A[15][15] * mat_B[15][9] +
                  mat_A[15][16] * mat_B[16][9] +
                  mat_A[15][17] * mat_B[17][9] +
                  mat_A[15][18] * mat_B[18][9] +
                  mat_A[15][19] * mat_B[19][9] +
                  mat_A[15][20] * mat_B[20][9] +
                  mat_A[15][21] * mat_B[21][9] +
                  mat_A[15][22] * mat_B[22][9] +
                  mat_A[15][23] * mat_B[23][9] +
                  mat_A[15][24] * mat_B[24][9] +
                  mat_A[15][25] * mat_B[25][9] +
                  mat_A[15][26] * mat_B[26][9] +
                  mat_A[15][27] * mat_B[27][9] +
                  mat_A[15][28] * mat_B[28][9] +
                  mat_A[15][29] * mat_B[29][9] +
                  mat_A[15][30] * mat_B[30][9] +
                  mat_A[15][31] * mat_B[31][9];
    mat_C[15][10] <= 
                  mat_A[15][0] * mat_B[0][10] +
                  mat_A[15][1] * mat_B[1][10] +
                  mat_A[15][2] * mat_B[2][10] +
                  mat_A[15][3] * mat_B[3][10] +
                  mat_A[15][4] * mat_B[4][10] +
                  mat_A[15][5] * mat_B[5][10] +
                  mat_A[15][6] * mat_B[6][10] +
                  mat_A[15][7] * mat_B[7][10] +
                  mat_A[15][8] * mat_B[8][10] +
                  mat_A[15][9] * mat_B[9][10] +
                  mat_A[15][10] * mat_B[10][10] +
                  mat_A[15][11] * mat_B[11][10] +
                  mat_A[15][12] * mat_B[12][10] +
                  mat_A[15][13] * mat_B[13][10] +
                  mat_A[15][14] * mat_B[14][10] +
                  mat_A[15][15] * mat_B[15][10] +
                  mat_A[15][16] * mat_B[16][10] +
                  mat_A[15][17] * mat_B[17][10] +
                  mat_A[15][18] * mat_B[18][10] +
                  mat_A[15][19] * mat_B[19][10] +
                  mat_A[15][20] * mat_B[20][10] +
                  mat_A[15][21] * mat_B[21][10] +
                  mat_A[15][22] * mat_B[22][10] +
                  mat_A[15][23] * mat_B[23][10] +
                  mat_A[15][24] * mat_B[24][10] +
                  mat_A[15][25] * mat_B[25][10] +
                  mat_A[15][26] * mat_B[26][10] +
                  mat_A[15][27] * mat_B[27][10] +
                  mat_A[15][28] * mat_B[28][10] +
                  mat_A[15][29] * mat_B[29][10] +
                  mat_A[15][30] * mat_B[30][10] +
                  mat_A[15][31] * mat_B[31][10];
    mat_C[15][11] <= 
                  mat_A[15][0] * mat_B[0][11] +
                  mat_A[15][1] * mat_B[1][11] +
                  mat_A[15][2] * mat_B[2][11] +
                  mat_A[15][3] * mat_B[3][11] +
                  mat_A[15][4] * mat_B[4][11] +
                  mat_A[15][5] * mat_B[5][11] +
                  mat_A[15][6] * mat_B[6][11] +
                  mat_A[15][7] * mat_B[7][11] +
                  mat_A[15][8] * mat_B[8][11] +
                  mat_A[15][9] * mat_B[9][11] +
                  mat_A[15][10] * mat_B[10][11] +
                  mat_A[15][11] * mat_B[11][11] +
                  mat_A[15][12] * mat_B[12][11] +
                  mat_A[15][13] * mat_B[13][11] +
                  mat_A[15][14] * mat_B[14][11] +
                  mat_A[15][15] * mat_B[15][11] +
                  mat_A[15][16] * mat_B[16][11] +
                  mat_A[15][17] * mat_B[17][11] +
                  mat_A[15][18] * mat_B[18][11] +
                  mat_A[15][19] * mat_B[19][11] +
                  mat_A[15][20] * mat_B[20][11] +
                  mat_A[15][21] * mat_B[21][11] +
                  mat_A[15][22] * mat_B[22][11] +
                  mat_A[15][23] * mat_B[23][11] +
                  mat_A[15][24] * mat_B[24][11] +
                  mat_A[15][25] * mat_B[25][11] +
                  mat_A[15][26] * mat_B[26][11] +
                  mat_A[15][27] * mat_B[27][11] +
                  mat_A[15][28] * mat_B[28][11] +
                  mat_A[15][29] * mat_B[29][11] +
                  mat_A[15][30] * mat_B[30][11] +
                  mat_A[15][31] * mat_B[31][11];
    mat_C[15][12] <= 
                  mat_A[15][0] * mat_B[0][12] +
                  mat_A[15][1] * mat_B[1][12] +
                  mat_A[15][2] * mat_B[2][12] +
                  mat_A[15][3] * mat_B[3][12] +
                  mat_A[15][4] * mat_B[4][12] +
                  mat_A[15][5] * mat_B[5][12] +
                  mat_A[15][6] * mat_B[6][12] +
                  mat_A[15][7] * mat_B[7][12] +
                  mat_A[15][8] * mat_B[8][12] +
                  mat_A[15][9] * mat_B[9][12] +
                  mat_A[15][10] * mat_B[10][12] +
                  mat_A[15][11] * mat_B[11][12] +
                  mat_A[15][12] * mat_B[12][12] +
                  mat_A[15][13] * mat_B[13][12] +
                  mat_A[15][14] * mat_B[14][12] +
                  mat_A[15][15] * mat_B[15][12] +
                  mat_A[15][16] * mat_B[16][12] +
                  mat_A[15][17] * mat_B[17][12] +
                  mat_A[15][18] * mat_B[18][12] +
                  mat_A[15][19] * mat_B[19][12] +
                  mat_A[15][20] * mat_B[20][12] +
                  mat_A[15][21] * mat_B[21][12] +
                  mat_A[15][22] * mat_B[22][12] +
                  mat_A[15][23] * mat_B[23][12] +
                  mat_A[15][24] * mat_B[24][12] +
                  mat_A[15][25] * mat_B[25][12] +
                  mat_A[15][26] * mat_B[26][12] +
                  mat_A[15][27] * mat_B[27][12] +
                  mat_A[15][28] * mat_B[28][12] +
                  mat_A[15][29] * mat_B[29][12] +
                  mat_A[15][30] * mat_B[30][12] +
                  mat_A[15][31] * mat_B[31][12];
    mat_C[15][13] <= 
                  mat_A[15][0] * mat_B[0][13] +
                  mat_A[15][1] * mat_B[1][13] +
                  mat_A[15][2] * mat_B[2][13] +
                  mat_A[15][3] * mat_B[3][13] +
                  mat_A[15][4] * mat_B[4][13] +
                  mat_A[15][5] * mat_B[5][13] +
                  mat_A[15][6] * mat_B[6][13] +
                  mat_A[15][7] * mat_B[7][13] +
                  mat_A[15][8] * mat_B[8][13] +
                  mat_A[15][9] * mat_B[9][13] +
                  mat_A[15][10] * mat_B[10][13] +
                  mat_A[15][11] * mat_B[11][13] +
                  mat_A[15][12] * mat_B[12][13] +
                  mat_A[15][13] * mat_B[13][13] +
                  mat_A[15][14] * mat_B[14][13] +
                  mat_A[15][15] * mat_B[15][13] +
                  mat_A[15][16] * mat_B[16][13] +
                  mat_A[15][17] * mat_B[17][13] +
                  mat_A[15][18] * mat_B[18][13] +
                  mat_A[15][19] * mat_B[19][13] +
                  mat_A[15][20] * mat_B[20][13] +
                  mat_A[15][21] * mat_B[21][13] +
                  mat_A[15][22] * mat_B[22][13] +
                  mat_A[15][23] * mat_B[23][13] +
                  mat_A[15][24] * mat_B[24][13] +
                  mat_A[15][25] * mat_B[25][13] +
                  mat_A[15][26] * mat_B[26][13] +
                  mat_A[15][27] * mat_B[27][13] +
                  mat_A[15][28] * mat_B[28][13] +
                  mat_A[15][29] * mat_B[29][13] +
                  mat_A[15][30] * mat_B[30][13] +
                  mat_A[15][31] * mat_B[31][13];
    mat_C[15][14] <= 
                  mat_A[15][0] * mat_B[0][14] +
                  mat_A[15][1] * mat_B[1][14] +
                  mat_A[15][2] * mat_B[2][14] +
                  mat_A[15][3] * mat_B[3][14] +
                  mat_A[15][4] * mat_B[4][14] +
                  mat_A[15][5] * mat_B[5][14] +
                  mat_A[15][6] * mat_B[6][14] +
                  mat_A[15][7] * mat_B[7][14] +
                  mat_A[15][8] * mat_B[8][14] +
                  mat_A[15][9] * mat_B[9][14] +
                  mat_A[15][10] * mat_B[10][14] +
                  mat_A[15][11] * mat_B[11][14] +
                  mat_A[15][12] * mat_B[12][14] +
                  mat_A[15][13] * mat_B[13][14] +
                  mat_A[15][14] * mat_B[14][14] +
                  mat_A[15][15] * mat_B[15][14] +
                  mat_A[15][16] * mat_B[16][14] +
                  mat_A[15][17] * mat_B[17][14] +
                  mat_A[15][18] * mat_B[18][14] +
                  mat_A[15][19] * mat_B[19][14] +
                  mat_A[15][20] * mat_B[20][14] +
                  mat_A[15][21] * mat_B[21][14] +
                  mat_A[15][22] * mat_B[22][14] +
                  mat_A[15][23] * mat_B[23][14] +
                  mat_A[15][24] * mat_B[24][14] +
                  mat_A[15][25] * mat_B[25][14] +
                  mat_A[15][26] * mat_B[26][14] +
                  mat_A[15][27] * mat_B[27][14] +
                  mat_A[15][28] * mat_B[28][14] +
                  mat_A[15][29] * mat_B[29][14] +
                  mat_A[15][30] * mat_B[30][14] +
                  mat_A[15][31] * mat_B[31][14];
    mat_C[15][15] <= 
                  mat_A[15][0] * mat_B[0][15] +
                  mat_A[15][1] * mat_B[1][15] +
                  mat_A[15][2] * mat_B[2][15] +
                  mat_A[15][3] * mat_B[3][15] +
                  mat_A[15][4] * mat_B[4][15] +
                  mat_A[15][5] * mat_B[5][15] +
                  mat_A[15][6] * mat_B[6][15] +
                  mat_A[15][7] * mat_B[7][15] +
                  mat_A[15][8] * mat_B[8][15] +
                  mat_A[15][9] * mat_B[9][15] +
                  mat_A[15][10] * mat_B[10][15] +
                  mat_A[15][11] * mat_B[11][15] +
                  mat_A[15][12] * mat_B[12][15] +
                  mat_A[15][13] * mat_B[13][15] +
                  mat_A[15][14] * mat_B[14][15] +
                  mat_A[15][15] * mat_B[15][15] +
                  mat_A[15][16] * mat_B[16][15] +
                  mat_A[15][17] * mat_B[17][15] +
                  mat_A[15][18] * mat_B[18][15] +
                  mat_A[15][19] * mat_B[19][15] +
                  mat_A[15][20] * mat_B[20][15] +
                  mat_A[15][21] * mat_B[21][15] +
                  mat_A[15][22] * mat_B[22][15] +
                  mat_A[15][23] * mat_B[23][15] +
                  mat_A[15][24] * mat_B[24][15] +
                  mat_A[15][25] * mat_B[25][15] +
                  mat_A[15][26] * mat_B[26][15] +
                  mat_A[15][27] * mat_B[27][15] +
                  mat_A[15][28] * mat_B[28][15] +
                  mat_A[15][29] * mat_B[29][15] +
                  mat_A[15][30] * mat_B[30][15] +
                  mat_A[15][31] * mat_B[31][15];
    mat_C[15][16] <= 
                  mat_A[15][0] * mat_B[0][16] +
                  mat_A[15][1] * mat_B[1][16] +
                  mat_A[15][2] * mat_B[2][16] +
                  mat_A[15][3] * mat_B[3][16] +
                  mat_A[15][4] * mat_B[4][16] +
                  mat_A[15][5] * mat_B[5][16] +
                  mat_A[15][6] * mat_B[6][16] +
                  mat_A[15][7] * mat_B[7][16] +
                  mat_A[15][8] * mat_B[8][16] +
                  mat_A[15][9] * mat_B[9][16] +
                  mat_A[15][10] * mat_B[10][16] +
                  mat_A[15][11] * mat_B[11][16] +
                  mat_A[15][12] * mat_B[12][16] +
                  mat_A[15][13] * mat_B[13][16] +
                  mat_A[15][14] * mat_B[14][16] +
                  mat_A[15][15] * mat_B[15][16] +
                  mat_A[15][16] * mat_B[16][16] +
                  mat_A[15][17] * mat_B[17][16] +
                  mat_A[15][18] * mat_B[18][16] +
                  mat_A[15][19] * mat_B[19][16] +
                  mat_A[15][20] * mat_B[20][16] +
                  mat_A[15][21] * mat_B[21][16] +
                  mat_A[15][22] * mat_B[22][16] +
                  mat_A[15][23] * mat_B[23][16] +
                  mat_A[15][24] * mat_B[24][16] +
                  mat_A[15][25] * mat_B[25][16] +
                  mat_A[15][26] * mat_B[26][16] +
                  mat_A[15][27] * mat_B[27][16] +
                  mat_A[15][28] * mat_B[28][16] +
                  mat_A[15][29] * mat_B[29][16] +
                  mat_A[15][30] * mat_B[30][16] +
                  mat_A[15][31] * mat_B[31][16];
    mat_C[15][17] <= 
                  mat_A[15][0] * mat_B[0][17] +
                  mat_A[15][1] * mat_B[1][17] +
                  mat_A[15][2] * mat_B[2][17] +
                  mat_A[15][3] * mat_B[3][17] +
                  mat_A[15][4] * mat_B[4][17] +
                  mat_A[15][5] * mat_B[5][17] +
                  mat_A[15][6] * mat_B[6][17] +
                  mat_A[15][7] * mat_B[7][17] +
                  mat_A[15][8] * mat_B[8][17] +
                  mat_A[15][9] * mat_B[9][17] +
                  mat_A[15][10] * mat_B[10][17] +
                  mat_A[15][11] * mat_B[11][17] +
                  mat_A[15][12] * mat_B[12][17] +
                  mat_A[15][13] * mat_B[13][17] +
                  mat_A[15][14] * mat_B[14][17] +
                  mat_A[15][15] * mat_B[15][17] +
                  mat_A[15][16] * mat_B[16][17] +
                  mat_A[15][17] * mat_B[17][17] +
                  mat_A[15][18] * mat_B[18][17] +
                  mat_A[15][19] * mat_B[19][17] +
                  mat_A[15][20] * mat_B[20][17] +
                  mat_A[15][21] * mat_B[21][17] +
                  mat_A[15][22] * mat_B[22][17] +
                  mat_A[15][23] * mat_B[23][17] +
                  mat_A[15][24] * mat_B[24][17] +
                  mat_A[15][25] * mat_B[25][17] +
                  mat_A[15][26] * mat_B[26][17] +
                  mat_A[15][27] * mat_B[27][17] +
                  mat_A[15][28] * mat_B[28][17] +
                  mat_A[15][29] * mat_B[29][17] +
                  mat_A[15][30] * mat_B[30][17] +
                  mat_A[15][31] * mat_B[31][17];
    mat_C[15][18] <= 
                  mat_A[15][0] * mat_B[0][18] +
                  mat_A[15][1] * mat_B[1][18] +
                  mat_A[15][2] * mat_B[2][18] +
                  mat_A[15][3] * mat_B[3][18] +
                  mat_A[15][4] * mat_B[4][18] +
                  mat_A[15][5] * mat_B[5][18] +
                  mat_A[15][6] * mat_B[6][18] +
                  mat_A[15][7] * mat_B[7][18] +
                  mat_A[15][8] * mat_B[8][18] +
                  mat_A[15][9] * mat_B[9][18] +
                  mat_A[15][10] * mat_B[10][18] +
                  mat_A[15][11] * mat_B[11][18] +
                  mat_A[15][12] * mat_B[12][18] +
                  mat_A[15][13] * mat_B[13][18] +
                  mat_A[15][14] * mat_B[14][18] +
                  mat_A[15][15] * mat_B[15][18] +
                  mat_A[15][16] * mat_B[16][18] +
                  mat_A[15][17] * mat_B[17][18] +
                  mat_A[15][18] * mat_B[18][18] +
                  mat_A[15][19] * mat_B[19][18] +
                  mat_A[15][20] * mat_B[20][18] +
                  mat_A[15][21] * mat_B[21][18] +
                  mat_A[15][22] * mat_B[22][18] +
                  mat_A[15][23] * mat_B[23][18] +
                  mat_A[15][24] * mat_B[24][18] +
                  mat_A[15][25] * mat_B[25][18] +
                  mat_A[15][26] * mat_B[26][18] +
                  mat_A[15][27] * mat_B[27][18] +
                  mat_A[15][28] * mat_B[28][18] +
                  mat_A[15][29] * mat_B[29][18] +
                  mat_A[15][30] * mat_B[30][18] +
                  mat_A[15][31] * mat_B[31][18];
    mat_C[15][19] <= 
                  mat_A[15][0] * mat_B[0][19] +
                  mat_A[15][1] * mat_B[1][19] +
                  mat_A[15][2] * mat_B[2][19] +
                  mat_A[15][3] * mat_B[3][19] +
                  mat_A[15][4] * mat_B[4][19] +
                  mat_A[15][5] * mat_B[5][19] +
                  mat_A[15][6] * mat_B[6][19] +
                  mat_A[15][7] * mat_B[7][19] +
                  mat_A[15][8] * mat_B[8][19] +
                  mat_A[15][9] * mat_B[9][19] +
                  mat_A[15][10] * mat_B[10][19] +
                  mat_A[15][11] * mat_B[11][19] +
                  mat_A[15][12] * mat_B[12][19] +
                  mat_A[15][13] * mat_B[13][19] +
                  mat_A[15][14] * mat_B[14][19] +
                  mat_A[15][15] * mat_B[15][19] +
                  mat_A[15][16] * mat_B[16][19] +
                  mat_A[15][17] * mat_B[17][19] +
                  mat_A[15][18] * mat_B[18][19] +
                  mat_A[15][19] * mat_B[19][19] +
                  mat_A[15][20] * mat_B[20][19] +
                  mat_A[15][21] * mat_B[21][19] +
                  mat_A[15][22] * mat_B[22][19] +
                  mat_A[15][23] * mat_B[23][19] +
                  mat_A[15][24] * mat_B[24][19] +
                  mat_A[15][25] * mat_B[25][19] +
                  mat_A[15][26] * mat_B[26][19] +
                  mat_A[15][27] * mat_B[27][19] +
                  mat_A[15][28] * mat_B[28][19] +
                  mat_A[15][29] * mat_B[29][19] +
                  mat_A[15][30] * mat_B[30][19] +
                  mat_A[15][31] * mat_B[31][19];
    mat_C[15][20] <= 
                  mat_A[15][0] * mat_B[0][20] +
                  mat_A[15][1] * mat_B[1][20] +
                  mat_A[15][2] * mat_B[2][20] +
                  mat_A[15][3] * mat_B[3][20] +
                  mat_A[15][4] * mat_B[4][20] +
                  mat_A[15][5] * mat_B[5][20] +
                  mat_A[15][6] * mat_B[6][20] +
                  mat_A[15][7] * mat_B[7][20] +
                  mat_A[15][8] * mat_B[8][20] +
                  mat_A[15][9] * mat_B[9][20] +
                  mat_A[15][10] * mat_B[10][20] +
                  mat_A[15][11] * mat_B[11][20] +
                  mat_A[15][12] * mat_B[12][20] +
                  mat_A[15][13] * mat_B[13][20] +
                  mat_A[15][14] * mat_B[14][20] +
                  mat_A[15][15] * mat_B[15][20] +
                  mat_A[15][16] * mat_B[16][20] +
                  mat_A[15][17] * mat_B[17][20] +
                  mat_A[15][18] * mat_B[18][20] +
                  mat_A[15][19] * mat_B[19][20] +
                  mat_A[15][20] * mat_B[20][20] +
                  mat_A[15][21] * mat_B[21][20] +
                  mat_A[15][22] * mat_B[22][20] +
                  mat_A[15][23] * mat_B[23][20] +
                  mat_A[15][24] * mat_B[24][20] +
                  mat_A[15][25] * mat_B[25][20] +
                  mat_A[15][26] * mat_B[26][20] +
                  mat_A[15][27] * mat_B[27][20] +
                  mat_A[15][28] * mat_B[28][20] +
                  mat_A[15][29] * mat_B[29][20] +
                  mat_A[15][30] * mat_B[30][20] +
                  mat_A[15][31] * mat_B[31][20];
    mat_C[15][21] <= 
                  mat_A[15][0] * mat_B[0][21] +
                  mat_A[15][1] * mat_B[1][21] +
                  mat_A[15][2] * mat_B[2][21] +
                  mat_A[15][3] * mat_B[3][21] +
                  mat_A[15][4] * mat_B[4][21] +
                  mat_A[15][5] * mat_B[5][21] +
                  mat_A[15][6] * mat_B[6][21] +
                  mat_A[15][7] * mat_B[7][21] +
                  mat_A[15][8] * mat_B[8][21] +
                  mat_A[15][9] * mat_B[9][21] +
                  mat_A[15][10] * mat_B[10][21] +
                  mat_A[15][11] * mat_B[11][21] +
                  mat_A[15][12] * mat_B[12][21] +
                  mat_A[15][13] * mat_B[13][21] +
                  mat_A[15][14] * mat_B[14][21] +
                  mat_A[15][15] * mat_B[15][21] +
                  mat_A[15][16] * mat_B[16][21] +
                  mat_A[15][17] * mat_B[17][21] +
                  mat_A[15][18] * mat_B[18][21] +
                  mat_A[15][19] * mat_B[19][21] +
                  mat_A[15][20] * mat_B[20][21] +
                  mat_A[15][21] * mat_B[21][21] +
                  mat_A[15][22] * mat_B[22][21] +
                  mat_A[15][23] * mat_B[23][21] +
                  mat_A[15][24] * mat_B[24][21] +
                  mat_A[15][25] * mat_B[25][21] +
                  mat_A[15][26] * mat_B[26][21] +
                  mat_A[15][27] * mat_B[27][21] +
                  mat_A[15][28] * mat_B[28][21] +
                  mat_A[15][29] * mat_B[29][21] +
                  mat_A[15][30] * mat_B[30][21] +
                  mat_A[15][31] * mat_B[31][21];
    mat_C[15][22] <= 
                  mat_A[15][0] * mat_B[0][22] +
                  mat_A[15][1] * mat_B[1][22] +
                  mat_A[15][2] * mat_B[2][22] +
                  mat_A[15][3] * mat_B[3][22] +
                  mat_A[15][4] * mat_B[4][22] +
                  mat_A[15][5] * mat_B[5][22] +
                  mat_A[15][6] * mat_B[6][22] +
                  mat_A[15][7] * mat_B[7][22] +
                  mat_A[15][8] * mat_B[8][22] +
                  mat_A[15][9] * mat_B[9][22] +
                  mat_A[15][10] * mat_B[10][22] +
                  mat_A[15][11] * mat_B[11][22] +
                  mat_A[15][12] * mat_B[12][22] +
                  mat_A[15][13] * mat_B[13][22] +
                  mat_A[15][14] * mat_B[14][22] +
                  mat_A[15][15] * mat_B[15][22] +
                  mat_A[15][16] * mat_B[16][22] +
                  mat_A[15][17] * mat_B[17][22] +
                  mat_A[15][18] * mat_B[18][22] +
                  mat_A[15][19] * mat_B[19][22] +
                  mat_A[15][20] * mat_B[20][22] +
                  mat_A[15][21] * mat_B[21][22] +
                  mat_A[15][22] * mat_B[22][22] +
                  mat_A[15][23] * mat_B[23][22] +
                  mat_A[15][24] * mat_B[24][22] +
                  mat_A[15][25] * mat_B[25][22] +
                  mat_A[15][26] * mat_B[26][22] +
                  mat_A[15][27] * mat_B[27][22] +
                  mat_A[15][28] * mat_B[28][22] +
                  mat_A[15][29] * mat_B[29][22] +
                  mat_A[15][30] * mat_B[30][22] +
                  mat_A[15][31] * mat_B[31][22];
    mat_C[15][23] <= 
                  mat_A[15][0] * mat_B[0][23] +
                  mat_A[15][1] * mat_B[1][23] +
                  mat_A[15][2] * mat_B[2][23] +
                  mat_A[15][3] * mat_B[3][23] +
                  mat_A[15][4] * mat_B[4][23] +
                  mat_A[15][5] * mat_B[5][23] +
                  mat_A[15][6] * mat_B[6][23] +
                  mat_A[15][7] * mat_B[7][23] +
                  mat_A[15][8] * mat_B[8][23] +
                  mat_A[15][9] * mat_B[9][23] +
                  mat_A[15][10] * mat_B[10][23] +
                  mat_A[15][11] * mat_B[11][23] +
                  mat_A[15][12] * mat_B[12][23] +
                  mat_A[15][13] * mat_B[13][23] +
                  mat_A[15][14] * mat_B[14][23] +
                  mat_A[15][15] * mat_B[15][23] +
                  mat_A[15][16] * mat_B[16][23] +
                  mat_A[15][17] * mat_B[17][23] +
                  mat_A[15][18] * mat_B[18][23] +
                  mat_A[15][19] * mat_B[19][23] +
                  mat_A[15][20] * mat_B[20][23] +
                  mat_A[15][21] * mat_B[21][23] +
                  mat_A[15][22] * mat_B[22][23] +
                  mat_A[15][23] * mat_B[23][23] +
                  mat_A[15][24] * mat_B[24][23] +
                  mat_A[15][25] * mat_B[25][23] +
                  mat_A[15][26] * mat_B[26][23] +
                  mat_A[15][27] * mat_B[27][23] +
                  mat_A[15][28] * mat_B[28][23] +
                  mat_A[15][29] * mat_B[29][23] +
                  mat_A[15][30] * mat_B[30][23] +
                  mat_A[15][31] * mat_B[31][23];
    mat_C[15][24] <= 
                  mat_A[15][0] * mat_B[0][24] +
                  mat_A[15][1] * mat_B[1][24] +
                  mat_A[15][2] * mat_B[2][24] +
                  mat_A[15][3] * mat_B[3][24] +
                  mat_A[15][4] * mat_B[4][24] +
                  mat_A[15][5] * mat_B[5][24] +
                  mat_A[15][6] * mat_B[6][24] +
                  mat_A[15][7] * mat_B[7][24] +
                  mat_A[15][8] * mat_B[8][24] +
                  mat_A[15][9] * mat_B[9][24] +
                  mat_A[15][10] * mat_B[10][24] +
                  mat_A[15][11] * mat_B[11][24] +
                  mat_A[15][12] * mat_B[12][24] +
                  mat_A[15][13] * mat_B[13][24] +
                  mat_A[15][14] * mat_B[14][24] +
                  mat_A[15][15] * mat_B[15][24] +
                  mat_A[15][16] * mat_B[16][24] +
                  mat_A[15][17] * mat_B[17][24] +
                  mat_A[15][18] * mat_B[18][24] +
                  mat_A[15][19] * mat_B[19][24] +
                  mat_A[15][20] * mat_B[20][24] +
                  mat_A[15][21] * mat_B[21][24] +
                  mat_A[15][22] * mat_B[22][24] +
                  mat_A[15][23] * mat_B[23][24] +
                  mat_A[15][24] * mat_B[24][24] +
                  mat_A[15][25] * mat_B[25][24] +
                  mat_A[15][26] * mat_B[26][24] +
                  mat_A[15][27] * mat_B[27][24] +
                  mat_A[15][28] * mat_B[28][24] +
                  mat_A[15][29] * mat_B[29][24] +
                  mat_A[15][30] * mat_B[30][24] +
                  mat_A[15][31] * mat_B[31][24];
    mat_C[15][25] <= 
                  mat_A[15][0] * mat_B[0][25] +
                  mat_A[15][1] * mat_B[1][25] +
                  mat_A[15][2] * mat_B[2][25] +
                  mat_A[15][3] * mat_B[3][25] +
                  mat_A[15][4] * mat_B[4][25] +
                  mat_A[15][5] * mat_B[5][25] +
                  mat_A[15][6] * mat_B[6][25] +
                  mat_A[15][7] * mat_B[7][25] +
                  mat_A[15][8] * mat_B[8][25] +
                  mat_A[15][9] * mat_B[9][25] +
                  mat_A[15][10] * mat_B[10][25] +
                  mat_A[15][11] * mat_B[11][25] +
                  mat_A[15][12] * mat_B[12][25] +
                  mat_A[15][13] * mat_B[13][25] +
                  mat_A[15][14] * mat_B[14][25] +
                  mat_A[15][15] * mat_B[15][25] +
                  mat_A[15][16] * mat_B[16][25] +
                  mat_A[15][17] * mat_B[17][25] +
                  mat_A[15][18] * mat_B[18][25] +
                  mat_A[15][19] * mat_B[19][25] +
                  mat_A[15][20] * mat_B[20][25] +
                  mat_A[15][21] * mat_B[21][25] +
                  mat_A[15][22] * mat_B[22][25] +
                  mat_A[15][23] * mat_B[23][25] +
                  mat_A[15][24] * mat_B[24][25] +
                  mat_A[15][25] * mat_B[25][25] +
                  mat_A[15][26] * mat_B[26][25] +
                  mat_A[15][27] * mat_B[27][25] +
                  mat_A[15][28] * mat_B[28][25] +
                  mat_A[15][29] * mat_B[29][25] +
                  mat_A[15][30] * mat_B[30][25] +
                  mat_A[15][31] * mat_B[31][25];
    mat_C[15][26] <= 
                  mat_A[15][0] * mat_B[0][26] +
                  mat_A[15][1] * mat_B[1][26] +
                  mat_A[15][2] * mat_B[2][26] +
                  mat_A[15][3] * mat_B[3][26] +
                  mat_A[15][4] * mat_B[4][26] +
                  mat_A[15][5] * mat_B[5][26] +
                  mat_A[15][6] * mat_B[6][26] +
                  mat_A[15][7] * mat_B[7][26] +
                  mat_A[15][8] * mat_B[8][26] +
                  mat_A[15][9] * mat_B[9][26] +
                  mat_A[15][10] * mat_B[10][26] +
                  mat_A[15][11] * mat_B[11][26] +
                  mat_A[15][12] * mat_B[12][26] +
                  mat_A[15][13] * mat_B[13][26] +
                  mat_A[15][14] * mat_B[14][26] +
                  mat_A[15][15] * mat_B[15][26] +
                  mat_A[15][16] * mat_B[16][26] +
                  mat_A[15][17] * mat_B[17][26] +
                  mat_A[15][18] * mat_B[18][26] +
                  mat_A[15][19] * mat_B[19][26] +
                  mat_A[15][20] * mat_B[20][26] +
                  mat_A[15][21] * mat_B[21][26] +
                  mat_A[15][22] * mat_B[22][26] +
                  mat_A[15][23] * mat_B[23][26] +
                  mat_A[15][24] * mat_B[24][26] +
                  mat_A[15][25] * mat_B[25][26] +
                  mat_A[15][26] * mat_B[26][26] +
                  mat_A[15][27] * mat_B[27][26] +
                  mat_A[15][28] * mat_B[28][26] +
                  mat_A[15][29] * mat_B[29][26] +
                  mat_A[15][30] * mat_B[30][26] +
                  mat_A[15][31] * mat_B[31][26];
    mat_C[15][27] <= 
                  mat_A[15][0] * mat_B[0][27] +
                  mat_A[15][1] * mat_B[1][27] +
                  mat_A[15][2] * mat_B[2][27] +
                  mat_A[15][3] * mat_B[3][27] +
                  mat_A[15][4] * mat_B[4][27] +
                  mat_A[15][5] * mat_B[5][27] +
                  mat_A[15][6] * mat_B[6][27] +
                  mat_A[15][7] * mat_B[7][27] +
                  mat_A[15][8] * mat_B[8][27] +
                  mat_A[15][9] * mat_B[9][27] +
                  mat_A[15][10] * mat_B[10][27] +
                  mat_A[15][11] * mat_B[11][27] +
                  mat_A[15][12] * mat_B[12][27] +
                  mat_A[15][13] * mat_B[13][27] +
                  mat_A[15][14] * mat_B[14][27] +
                  mat_A[15][15] * mat_B[15][27] +
                  mat_A[15][16] * mat_B[16][27] +
                  mat_A[15][17] * mat_B[17][27] +
                  mat_A[15][18] * mat_B[18][27] +
                  mat_A[15][19] * mat_B[19][27] +
                  mat_A[15][20] * mat_B[20][27] +
                  mat_A[15][21] * mat_B[21][27] +
                  mat_A[15][22] * mat_B[22][27] +
                  mat_A[15][23] * mat_B[23][27] +
                  mat_A[15][24] * mat_B[24][27] +
                  mat_A[15][25] * mat_B[25][27] +
                  mat_A[15][26] * mat_B[26][27] +
                  mat_A[15][27] * mat_B[27][27] +
                  mat_A[15][28] * mat_B[28][27] +
                  mat_A[15][29] * mat_B[29][27] +
                  mat_A[15][30] * mat_B[30][27] +
                  mat_A[15][31] * mat_B[31][27];
    mat_C[15][28] <= 
                  mat_A[15][0] * mat_B[0][28] +
                  mat_A[15][1] * mat_B[1][28] +
                  mat_A[15][2] * mat_B[2][28] +
                  mat_A[15][3] * mat_B[3][28] +
                  mat_A[15][4] * mat_B[4][28] +
                  mat_A[15][5] * mat_B[5][28] +
                  mat_A[15][6] * mat_B[6][28] +
                  mat_A[15][7] * mat_B[7][28] +
                  mat_A[15][8] * mat_B[8][28] +
                  mat_A[15][9] * mat_B[9][28] +
                  mat_A[15][10] * mat_B[10][28] +
                  mat_A[15][11] * mat_B[11][28] +
                  mat_A[15][12] * mat_B[12][28] +
                  mat_A[15][13] * mat_B[13][28] +
                  mat_A[15][14] * mat_B[14][28] +
                  mat_A[15][15] * mat_B[15][28] +
                  mat_A[15][16] * mat_B[16][28] +
                  mat_A[15][17] * mat_B[17][28] +
                  mat_A[15][18] * mat_B[18][28] +
                  mat_A[15][19] * mat_B[19][28] +
                  mat_A[15][20] * mat_B[20][28] +
                  mat_A[15][21] * mat_B[21][28] +
                  mat_A[15][22] * mat_B[22][28] +
                  mat_A[15][23] * mat_B[23][28] +
                  mat_A[15][24] * mat_B[24][28] +
                  mat_A[15][25] * mat_B[25][28] +
                  mat_A[15][26] * mat_B[26][28] +
                  mat_A[15][27] * mat_B[27][28] +
                  mat_A[15][28] * mat_B[28][28] +
                  mat_A[15][29] * mat_B[29][28] +
                  mat_A[15][30] * mat_B[30][28] +
                  mat_A[15][31] * mat_B[31][28];
    mat_C[15][29] <= 
                  mat_A[15][0] * mat_B[0][29] +
                  mat_A[15][1] * mat_B[1][29] +
                  mat_A[15][2] * mat_B[2][29] +
                  mat_A[15][3] * mat_B[3][29] +
                  mat_A[15][4] * mat_B[4][29] +
                  mat_A[15][5] * mat_B[5][29] +
                  mat_A[15][6] * mat_B[6][29] +
                  mat_A[15][7] * mat_B[7][29] +
                  mat_A[15][8] * mat_B[8][29] +
                  mat_A[15][9] * mat_B[9][29] +
                  mat_A[15][10] * mat_B[10][29] +
                  mat_A[15][11] * mat_B[11][29] +
                  mat_A[15][12] * mat_B[12][29] +
                  mat_A[15][13] * mat_B[13][29] +
                  mat_A[15][14] * mat_B[14][29] +
                  mat_A[15][15] * mat_B[15][29] +
                  mat_A[15][16] * mat_B[16][29] +
                  mat_A[15][17] * mat_B[17][29] +
                  mat_A[15][18] * mat_B[18][29] +
                  mat_A[15][19] * mat_B[19][29] +
                  mat_A[15][20] * mat_B[20][29] +
                  mat_A[15][21] * mat_B[21][29] +
                  mat_A[15][22] * mat_B[22][29] +
                  mat_A[15][23] * mat_B[23][29] +
                  mat_A[15][24] * mat_B[24][29] +
                  mat_A[15][25] * mat_B[25][29] +
                  mat_A[15][26] * mat_B[26][29] +
                  mat_A[15][27] * mat_B[27][29] +
                  mat_A[15][28] * mat_B[28][29] +
                  mat_A[15][29] * mat_B[29][29] +
                  mat_A[15][30] * mat_B[30][29] +
                  mat_A[15][31] * mat_B[31][29];
    mat_C[15][30] <= 
                  mat_A[15][0] * mat_B[0][30] +
                  mat_A[15][1] * mat_B[1][30] +
                  mat_A[15][2] * mat_B[2][30] +
                  mat_A[15][3] * mat_B[3][30] +
                  mat_A[15][4] * mat_B[4][30] +
                  mat_A[15][5] * mat_B[5][30] +
                  mat_A[15][6] * mat_B[6][30] +
                  mat_A[15][7] * mat_B[7][30] +
                  mat_A[15][8] * mat_B[8][30] +
                  mat_A[15][9] * mat_B[9][30] +
                  mat_A[15][10] * mat_B[10][30] +
                  mat_A[15][11] * mat_B[11][30] +
                  mat_A[15][12] * mat_B[12][30] +
                  mat_A[15][13] * mat_B[13][30] +
                  mat_A[15][14] * mat_B[14][30] +
                  mat_A[15][15] * mat_B[15][30] +
                  mat_A[15][16] * mat_B[16][30] +
                  mat_A[15][17] * mat_B[17][30] +
                  mat_A[15][18] * mat_B[18][30] +
                  mat_A[15][19] * mat_B[19][30] +
                  mat_A[15][20] * mat_B[20][30] +
                  mat_A[15][21] * mat_B[21][30] +
                  mat_A[15][22] * mat_B[22][30] +
                  mat_A[15][23] * mat_B[23][30] +
                  mat_A[15][24] * mat_B[24][30] +
                  mat_A[15][25] * mat_B[25][30] +
                  mat_A[15][26] * mat_B[26][30] +
                  mat_A[15][27] * mat_B[27][30] +
                  mat_A[15][28] * mat_B[28][30] +
                  mat_A[15][29] * mat_B[29][30] +
                  mat_A[15][30] * mat_B[30][30] +
                  mat_A[15][31] * mat_B[31][30];
    mat_C[15][31] <= 
                  mat_A[15][0] * mat_B[0][31] +
                  mat_A[15][1] * mat_B[1][31] +
                  mat_A[15][2] * mat_B[2][31] +
                  mat_A[15][3] * mat_B[3][31] +
                  mat_A[15][4] * mat_B[4][31] +
                  mat_A[15][5] * mat_B[5][31] +
                  mat_A[15][6] * mat_B[6][31] +
                  mat_A[15][7] * mat_B[7][31] +
                  mat_A[15][8] * mat_B[8][31] +
                  mat_A[15][9] * mat_B[9][31] +
                  mat_A[15][10] * mat_B[10][31] +
                  mat_A[15][11] * mat_B[11][31] +
                  mat_A[15][12] * mat_B[12][31] +
                  mat_A[15][13] * mat_B[13][31] +
                  mat_A[15][14] * mat_B[14][31] +
                  mat_A[15][15] * mat_B[15][31] +
                  mat_A[15][16] * mat_B[16][31] +
                  mat_A[15][17] * mat_B[17][31] +
                  mat_A[15][18] * mat_B[18][31] +
                  mat_A[15][19] * mat_B[19][31] +
                  mat_A[15][20] * mat_B[20][31] +
                  mat_A[15][21] * mat_B[21][31] +
                  mat_A[15][22] * mat_B[22][31] +
                  mat_A[15][23] * mat_B[23][31] +
                  mat_A[15][24] * mat_B[24][31] +
                  mat_A[15][25] * mat_B[25][31] +
                  mat_A[15][26] * mat_B[26][31] +
                  mat_A[15][27] * mat_B[27][31] +
                  mat_A[15][28] * mat_B[28][31] +
                  mat_A[15][29] * mat_B[29][31] +
                  mat_A[15][30] * mat_B[30][31] +
                  mat_A[15][31] * mat_B[31][31];
    mat_C[16][0] <= 
                  mat_A[16][0] * mat_B[0][0] +
                  mat_A[16][1] * mat_B[1][0] +
                  mat_A[16][2] * mat_B[2][0] +
                  mat_A[16][3] * mat_B[3][0] +
                  mat_A[16][4] * mat_B[4][0] +
                  mat_A[16][5] * mat_B[5][0] +
                  mat_A[16][6] * mat_B[6][0] +
                  mat_A[16][7] * mat_B[7][0] +
                  mat_A[16][8] * mat_B[8][0] +
                  mat_A[16][9] * mat_B[9][0] +
                  mat_A[16][10] * mat_B[10][0] +
                  mat_A[16][11] * mat_B[11][0] +
                  mat_A[16][12] * mat_B[12][0] +
                  mat_A[16][13] * mat_B[13][0] +
                  mat_A[16][14] * mat_B[14][0] +
                  mat_A[16][15] * mat_B[15][0] +
                  mat_A[16][16] * mat_B[16][0] +
                  mat_A[16][17] * mat_B[17][0] +
                  mat_A[16][18] * mat_B[18][0] +
                  mat_A[16][19] * mat_B[19][0] +
                  mat_A[16][20] * mat_B[20][0] +
                  mat_A[16][21] * mat_B[21][0] +
                  mat_A[16][22] * mat_B[22][0] +
                  mat_A[16][23] * mat_B[23][0] +
                  mat_A[16][24] * mat_B[24][0] +
                  mat_A[16][25] * mat_B[25][0] +
                  mat_A[16][26] * mat_B[26][0] +
                  mat_A[16][27] * mat_B[27][0] +
                  mat_A[16][28] * mat_B[28][0] +
                  mat_A[16][29] * mat_B[29][0] +
                  mat_A[16][30] * mat_B[30][0] +
                  mat_A[16][31] * mat_B[31][0];
    mat_C[16][1] <= 
                  mat_A[16][0] * mat_B[0][1] +
                  mat_A[16][1] * mat_B[1][1] +
                  mat_A[16][2] * mat_B[2][1] +
                  mat_A[16][3] * mat_B[3][1] +
                  mat_A[16][4] * mat_B[4][1] +
                  mat_A[16][5] * mat_B[5][1] +
                  mat_A[16][6] * mat_B[6][1] +
                  mat_A[16][7] * mat_B[7][1] +
                  mat_A[16][8] * mat_B[8][1] +
                  mat_A[16][9] * mat_B[9][1] +
                  mat_A[16][10] * mat_B[10][1] +
                  mat_A[16][11] * mat_B[11][1] +
                  mat_A[16][12] * mat_B[12][1] +
                  mat_A[16][13] * mat_B[13][1] +
                  mat_A[16][14] * mat_B[14][1] +
                  mat_A[16][15] * mat_B[15][1] +
                  mat_A[16][16] * mat_B[16][1] +
                  mat_A[16][17] * mat_B[17][1] +
                  mat_A[16][18] * mat_B[18][1] +
                  mat_A[16][19] * mat_B[19][1] +
                  mat_A[16][20] * mat_B[20][1] +
                  mat_A[16][21] * mat_B[21][1] +
                  mat_A[16][22] * mat_B[22][1] +
                  mat_A[16][23] * mat_B[23][1] +
                  mat_A[16][24] * mat_B[24][1] +
                  mat_A[16][25] * mat_B[25][1] +
                  mat_A[16][26] * mat_B[26][1] +
                  mat_A[16][27] * mat_B[27][1] +
                  mat_A[16][28] * mat_B[28][1] +
                  mat_A[16][29] * mat_B[29][1] +
                  mat_A[16][30] * mat_B[30][1] +
                  mat_A[16][31] * mat_B[31][1];
    mat_C[16][2] <= 
                  mat_A[16][0] * mat_B[0][2] +
                  mat_A[16][1] * mat_B[1][2] +
                  mat_A[16][2] * mat_B[2][2] +
                  mat_A[16][3] * mat_B[3][2] +
                  mat_A[16][4] * mat_B[4][2] +
                  mat_A[16][5] * mat_B[5][2] +
                  mat_A[16][6] * mat_B[6][2] +
                  mat_A[16][7] * mat_B[7][2] +
                  mat_A[16][8] * mat_B[8][2] +
                  mat_A[16][9] * mat_B[9][2] +
                  mat_A[16][10] * mat_B[10][2] +
                  mat_A[16][11] * mat_B[11][2] +
                  mat_A[16][12] * mat_B[12][2] +
                  mat_A[16][13] * mat_B[13][2] +
                  mat_A[16][14] * mat_B[14][2] +
                  mat_A[16][15] * mat_B[15][2] +
                  mat_A[16][16] * mat_B[16][2] +
                  mat_A[16][17] * mat_B[17][2] +
                  mat_A[16][18] * mat_B[18][2] +
                  mat_A[16][19] * mat_B[19][2] +
                  mat_A[16][20] * mat_B[20][2] +
                  mat_A[16][21] * mat_B[21][2] +
                  mat_A[16][22] * mat_B[22][2] +
                  mat_A[16][23] * mat_B[23][2] +
                  mat_A[16][24] * mat_B[24][2] +
                  mat_A[16][25] * mat_B[25][2] +
                  mat_A[16][26] * mat_B[26][2] +
                  mat_A[16][27] * mat_B[27][2] +
                  mat_A[16][28] * mat_B[28][2] +
                  mat_A[16][29] * mat_B[29][2] +
                  mat_A[16][30] * mat_B[30][2] +
                  mat_A[16][31] * mat_B[31][2];
    mat_C[16][3] <= 
                  mat_A[16][0] * mat_B[0][3] +
                  mat_A[16][1] * mat_B[1][3] +
                  mat_A[16][2] * mat_B[2][3] +
                  mat_A[16][3] * mat_B[3][3] +
                  mat_A[16][4] * mat_B[4][3] +
                  mat_A[16][5] * mat_B[5][3] +
                  mat_A[16][6] * mat_B[6][3] +
                  mat_A[16][7] * mat_B[7][3] +
                  mat_A[16][8] * mat_B[8][3] +
                  mat_A[16][9] * mat_B[9][3] +
                  mat_A[16][10] * mat_B[10][3] +
                  mat_A[16][11] * mat_B[11][3] +
                  mat_A[16][12] * mat_B[12][3] +
                  mat_A[16][13] * mat_B[13][3] +
                  mat_A[16][14] * mat_B[14][3] +
                  mat_A[16][15] * mat_B[15][3] +
                  mat_A[16][16] * mat_B[16][3] +
                  mat_A[16][17] * mat_B[17][3] +
                  mat_A[16][18] * mat_B[18][3] +
                  mat_A[16][19] * mat_B[19][3] +
                  mat_A[16][20] * mat_B[20][3] +
                  mat_A[16][21] * mat_B[21][3] +
                  mat_A[16][22] * mat_B[22][3] +
                  mat_A[16][23] * mat_B[23][3] +
                  mat_A[16][24] * mat_B[24][3] +
                  mat_A[16][25] * mat_B[25][3] +
                  mat_A[16][26] * mat_B[26][3] +
                  mat_A[16][27] * mat_B[27][3] +
                  mat_A[16][28] * mat_B[28][3] +
                  mat_A[16][29] * mat_B[29][3] +
                  mat_A[16][30] * mat_B[30][3] +
                  mat_A[16][31] * mat_B[31][3];
    mat_C[16][4] <= 
                  mat_A[16][0] * mat_B[0][4] +
                  mat_A[16][1] * mat_B[1][4] +
                  mat_A[16][2] * mat_B[2][4] +
                  mat_A[16][3] * mat_B[3][4] +
                  mat_A[16][4] * mat_B[4][4] +
                  mat_A[16][5] * mat_B[5][4] +
                  mat_A[16][6] * mat_B[6][4] +
                  mat_A[16][7] * mat_B[7][4] +
                  mat_A[16][8] * mat_B[8][4] +
                  mat_A[16][9] * mat_B[9][4] +
                  mat_A[16][10] * mat_B[10][4] +
                  mat_A[16][11] * mat_B[11][4] +
                  mat_A[16][12] * mat_B[12][4] +
                  mat_A[16][13] * mat_B[13][4] +
                  mat_A[16][14] * mat_B[14][4] +
                  mat_A[16][15] * mat_B[15][4] +
                  mat_A[16][16] * mat_B[16][4] +
                  mat_A[16][17] * mat_B[17][4] +
                  mat_A[16][18] * mat_B[18][4] +
                  mat_A[16][19] * mat_B[19][4] +
                  mat_A[16][20] * mat_B[20][4] +
                  mat_A[16][21] * mat_B[21][4] +
                  mat_A[16][22] * mat_B[22][4] +
                  mat_A[16][23] * mat_B[23][4] +
                  mat_A[16][24] * mat_B[24][4] +
                  mat_A[16][25] * mat_B[25][4] +
                  mat_A[16][26] * mat_B[26][4] +
                  mat_A[16][27] * mat_B[27][4] +
                  mat_A[16][28] * mat_B[28][4] +
                  mat_A[16][29] * mat_B[29][4] +
                  mat_A[16][30] * mat_B[30][4] +
                  mat_A[16][31] * mat_B[31][4];
    mat_C[16][5] <= 
                  mat_A[16][0] * mat_B[0][5] +
                  mat_A[16][1] * mat_B[1][5] +
                  mat_A[16][2] * mat_B[2][5] +
                  mat_A[16][3] * mat_B[3][5] +
                  mat_A[16][4] * mat_B[4][5] +
                  mat_A[16][5] * mat_B[5][5] +
                  mat_A[16][6] * mat_B[6][5] +
                  mat_A[16][7] * mat_B[7][5] +
                  mat_A[16][8] * mat_B[8][5] +
                  mat_A[16][9] * mat_B[9][5] +
                  mat_A[16][10] * mat_B[10][5] +
                  mat_A[16][11] * mat_B[11][5] +
                  mat_A[16][12] * mat_B[12][5] +
                  mat_A[16][13] * mat_B[13][5] +
                  mat_A[16][14] * mat_B[14][5] +
                  mat_A[16][15] * mat_B[15][5] +
                  mat_A[16][16] * mat_B[16][5] +
                  mat_A[16][17] * mat_B[17][5] +
                  mat_A[16][18] * mat_B[18][5] +
                  mat_A[16][19] * mat_B[19][5] +
                  mat_A[16][20] * mat_B[20][5] +
                  mat_A[16][21] * mat_B[21][5] +
                  mat_A[16][22] * mat_B[22][5] +
                  mat_A[16][23] * mat_B[23][5] +
                  mat_A[16][24] * mat_B[24][5] +
                  mat_A[16][25] * mat_B[25][5] +
                  mat_A[16][26] * mat_B[26][5] +
                  mat_A[16][27] * mat_B[27][5] +
                  mat_A[16][28] * mat_B[28][5] +
                  mat_A[16][29] * mat_B[29][5] +
                  mat_A[16][30] * mat_B[30][5] +
                  mat_A[16][31] * mat_B[31][5];
    mat_C[16][6] <= 
                  mat_A[16][0] * mat_B[0][6] +
                  mat_A[16][1] * mat_B[1][6] +
                  mat_A[16][2] * mat_B[2][6] +
                  mat_A[16][3] * mat_B[3][6] +
                  mat_A[16][4] * mat_B[4][6] +
                  mat_A[16][5] * mat_B[5][6] +
                  mat_A[16][6] * mat_B[6][6] +
                  mat_A[16][7] * mat_B[7][6] +
                  mat_A[16][8] * mat_B[8][6] +
                  mat_A[16][9] * mat_B[9][6] +
                  mat_A[16][10] * mat_B[10][6] +
                  mat_A[16][11] * mat_B[11][6] +
                  mat_A[16][12] * mat_B[12][6] +
                  mat_A[16][13] * mat_B[13][6] +
                  mat_A[16][14] * mat_B[14][6] +
                  mat_A[16][15] * mat_B[15][6] +
                  mat_A[16][16] * mat_B[16][6] +
                  mat_A[16][17] * mat_B[17][6] +
                  mat_A[16][18] * mat_B[18][6] +
                  mat_A[16][19] * mat_B[19][6] +
                  mat_A[16][20] * mat_B[20][6] +
                  mat_A[16][21] * mat_B[21][6] +
                  mat_A[16][22] * mat_B[22][6] +
                  mat_A[16][23] * mat_B[23][6] +
                  mat_A[16][24] * mat_B[24][6] +
                  mat_A[16][25] * mat_B[25][6] +
                  mat_A[16][26] * mat_B[26][6] +
                  mat_A[16][27] * mat_B[27][6] +
                  mat_A[16][28] * mat_B[28][6] +
                  mat_A[16][29] * mat_B[29][6] +
                  mat_A[16][30] * mat_B[30][6] +
                  mat_A[16][31] * mat_B[31][6];
    mat_C[16][7] <= 
                  mat_A[16][0] * mat_B[0][7] +
                  mat_A[16][1] * mat_B[1][7] +
                  mat_A[16][2] * mat_B[2][7] +
                  mat_A[16][3] * mat_B[3][7] +
                  mat_A[16][4] * mat_B[4][7] +
                  mat_A[16][5] * mat_B[5][7] +
                  mat_A[16][6] * mat_B[6][7] +
                  mat_A[16][7] * mat_B[7][7] +
                  mat_A[16][8] * mat_B[8][7] +
                  mat_A[16][9] * mat_B[9][7] +
                  mat_A[16][10] * mat_B[10][7] +
                  mat_A[16][11] * mat_B[11][7] +
                  mat_A[16][12] * mat_B[12][7] +
                  mat_A[16][13] * mat_B[13][7] +
                  mat_A[16][14] * mat_B[14][7] +
                  mat_A[16][15] * mat_B[15][7] +
                  mat_A[16][16] * mat_B[16][7] +
                  mat_A[16][17] * mat_B[17][7] +
                  mat_A[16][18] * mat_B[18][7] +
                  mat_A[16][19] * mat_B[19][7] +
                  mat_A[16][20] * mat_B[20][7] +
                  mat_A[16][21] * mat_B[21][7] +
                  mat_A[16][22] * mat_B[22][7] +
                  mat_A[16][23] * mat_B[23][7] +
                  mat_A[16][24] * mat_B[24][7] +
                  mat_A[16][25] * mat_B[25][7] +
                  mat_A[16][26] * mat_B[26][7] +
                  mat_A[16][27] * mat_B[27][7] +
                  mat_A[16][28] * mat_B[28][7] +
                  mat_A[16][29] * mat_B[29][7] +
                  mat_A[16][30] * mat_B[30][7] +
                  mat_A[16][31] * mat_B[31][7];
    mat_C[16][8] <= 
                  mat_A[16][0] * mat_B[0][8] +
                  mat_A[16][1] * mat_B[1][8] +
                  mat_A[16][2] * mat_B[2][8] +
                  mat_A[16][3] * mat_B[3][8] +
                  mat_A[16][4] * mat_B[4][8] +
                  mat_A[16][5] * mat_B[5][8] +
                  mat_A[16][6] * mat_B[6][8] +
                  mat_A[16][7] * mat_B[7][8] +
                  mat_A[16][8] * mat_B[8][8] +
                  mat_A[16][9] * mat_B[9][8] +
                  mat_A[16][10] * mat_B[10][8] +
                  mat_A[16][11] * mat_B[11][8] +
                  mat_A[16][12] * mat_B[12][8] +
                  mat_A[16][13] * mat_B[13][8] +
                  mat_A[16][14] * mat_B[14][8] +
                  mat_A[16][15] * mat_B[15][8] +
                  mat_A[16][16] * mat_B[16][8] +
                  mat_A[16][17] * mat_B[17][8] +
                  mat_A[16][18] * mat_B[18][8] +
                  mat_A[16][19] * mat_B[19][8] +
                  mat_A[16][20] * mat_B[20][8] +
                  mat_A[16][21] * mat_B[21][8] +
                  mat_A[16][22] * mat_B[22][8] +
                  mat_A[16][23] * mat_B[23][8] +
                  mat_A[16][24] * mat_B[24][8] +
                  mat_A[16][25] * mat_B[25][8] +
                  mat_A[16][26] * mat_B[26][8] +
                  mat_A[16][27] * mat_B[27][8] +
                  mat_A[16][28] * mat_B[28][8] +
                  mat_A[16][29] * mat_B[29][8] +
                  mat_A[16][30] * mat_B[30][8] +
                  mat_A[16][31] * mat_B[31][8];
    mat_C[16][9] <= 
                  mat_A[16][0] * mat_B[0][9] +
                  mat_A[16][1] * mat_B[1][9] +
                  mat_A[16][2] * mat_B[2][9] +
                  mat_A[16][3] * mat_B[3][9] +
                  mat_A[16][4] * mat_B[4][9] +
                  mat_A[16][5] * mat_B[5][9] +
                  mat_A[16][6] * mat_B[6][9] +
                  mat_A[16][7] * mat_B[7][9] +
                  mat_A[16][8] * mat_B[8][9] +
                  mat_A[16][9] * mat_B[9][9] +
                  mat_A[16][10] * mat_B[10][9] +
                  mat_A[16][11] * mat_B[11][9] +
                  mat_A[16][12] * mat_B[12][9] +
                  mat_A[16][13] * mat_B[13][9] +
                  mat_A[16][14] * mat_B[14][9] +
                  mat_A[16][15] * mat_B[15][9] +
                  mat_A[16][16] * mat_B[16][9] +
                  mat_A[16][17] * mat_B[17][9] +
                  mat_A[16][18] * mat_B[18][9] +
                  mat_A[16][19] * mat_B[19][9] +
                  mat_A[16][20] * mat_B[20][9] +
                  mat_A[16][21] * mat_B[21][9] +
                  mat_A[16][22] * mat_B[22][9] +
                  mat_A[16][23] * mat_B[23][9] +
                  mat_A[16][24] * mat_B[24][9] +
                  mat_A[16][25] * mat_B[25][9] +
                  mat_A[16][26] * mat_B[26][9] +
                  mat_A[16][27] * mat_B[27][9] +
                  mat_A[16][28] * mat_B[28][9] +
                  mat_A[16][29] * mat_B[29][9] +
                  mat_A[16][30] * mat_B[30][9] +
                  mat_A[16][31] * mat_B[31][9];
    mat_C[16][10] <= 
                  mat_A[16][0] * mat_B[0][10] +
                  mat_A[16][1] * mat_B[1][10] +
                  mat_A[16][2] * mat_B[2][10] +
                  mat_A[16][3] * mat_B[3][10] +
                  mat_A[16][4] * mat_B[4][10] +
                  mat_A[16][5] * mat_B[5][10] +
                  mat_A[16][6] * mat_B[6][10] +
                  mat_A[16][7] * mat_B[7][10] +
                  mat_A[16][8] * mat_B[8][10] +
                  mat_A[16][9] * mat_B[9][10] +
                  mat_A[16][10] * mat_B[10][10] +
                  mat_A[16][11] * mat_B[11][10] +
                  mat_A[16][12] * mat_B[12][10] +
                  mat_A[16][13] * mat_B[13][10] +
                  mat_A[16][14] * mat_B[14][10] +
                  mat_A[16][15] * mat_B[15][10] +
                  mat_A[16][16] * mat_B[16][10] +
                  mat_A[16][17] * mat_B[17][10] +
                  mat_A[16][18] * mat_B[18][10] +
                  mat_A[16][19] * mat_B[19][10] +
                  mat_A[16][20] * mat_B[20][10] +
                  mat_A[16][21] * mat_B[21][10] +
                  mat_A[16][22] * mat_B[22][10] +
                  mat_A[16][23] * mat_B[23][10] +
                  mat_A[16][24] * mat_B[24][10] +
                  mat_A[16][25] * mat_B[25][10] +
                  mat_A[16][26] * mat_B[26][10] +
                  mat_A[16][27] * mat_B[27][10] +
                  mat_A[16][28] * mat_B[28][10] +
                  mat_A[16][29] * mat_B[29][10] +
                  mat_A[16][30] * mat_B[30][10] +
                  mat_A[16][31] * mat_B[31][10];
    mat_C[16][11] <= 
                  mat_A[16][0] * mat_B[0][11] +
                  mat_A[16][1] * mat_B[1][11] +
                  mat_A[16][2] * mat_B[2][11] +
                  mat_A[16][3] * mat_B[3][11] +
                  mat_A[16][4] * mat_B[4][11] +
                  mat_A[16][5] * mat_B[5][11] +
                  mat_A[16][6] * mat_B[6][11] +
                  mat_A[16][7] * mat_B[7][11] +
                  mat_A[16][8] * mat_B[8][11] +
                  mat_A[16][9] * mat_B[9][11] +
                  mat_A[16][10] * mat_B[10][11] +
                  mat_A[16][11] * mat_B[11][11] +
                  mat_A[16][12] * mat_B[12][11] +
                  mat_A[16][13] * mat_B[13][11] +
                  mat_A[16][14] * mat_B[14][11] +
                  mat_A[16][15] * mat_B[15][11] +
                  mat_A[16][16] * mat_B[16][11] +
                  mat_A[16][17] * mat_B[17][11] +
                  mat_A[16][18] * mat_B[18][11] +
                  mat_A[16][19] * mat_B[19][11] +
                  mat_A[16][20] * mat_B[20][11] +
                  mat_A[16][21] * mat_B[21][11] +
                  mat_A[16][22] * mat_B[22][11] +
                  mat_A[16][23] * mat_B[23][11] +
                  mat_A[16][24] * mat_B[24][11] +
                  mat_A[16][25] * mat_B[25][11] +
                  mat_A[16][26] * mat_B[26][11] +
                  mat_A[16][27] * mat_B[27][11] +
                  mat_A[16][28] * mat_B[28][11] +
                  mat_A[16][29] * mat_B[29][11] +
                  mat_A[16][30] * mat_B[30][11] +
                  mat_A[16][31] * mat_B[31][11];
    mat_C[16][12] <= 
                  mat_A[16][0] * mat_B[0][12] +
                  mat_A[16][1] * mat_B[1][12] +
                  mat_A[16][2] * mat_B[2][12] +
                  mat_A[16][3] * mat_B[3][12] +
                  mat_A[16][4] * mat_B[4][12] +
                  mat_A[16][5] * mat_B[5][12] +
                  mat_A[16][6] * mat_B[6][12] +
                  mat_A[16][7] * mat_B[7][12] +
                  mat_A[16][8] * mat_B[8][12] +
                  mat_A[16][9] * mat_B[9][12] +
                  mat_A[16][10] * mat_B[10][12] +
                  mat_A[16][11] * mat_B[11][12] +
                  mat_A[16][12] * mat_B[12][12] +
                  mat_A[16][13] * mat_B[13][12] +
                  mat_A[16][14] * mat_B[14][12] +
                  mat_A[16][15] * mat_B[15][12] +
                  mat_A[16][16] * mat_B[16][12] +
                  mat_A[16][17] * mat_B[17][12] +
                  mat_A[16][18] * mat_B[18][12] +
                  mat_A[16][19] * mat_B[19][12] +
                  mat_A[16][20] * mat_B[20][12] +
                  mat_A[16][21] * mat_B[21][12] +
                  mat_A[16][22] * mat_B[22][12] +
                  mat_A[16][23] * mat_B[23][12] +
                  mat_A[16][24] * mat_B[24][12] +
                  mat_A[16][25] * mat_B[25][12] +
                  mat_A[16][26] * mat_B[26][12] +
                  mat_A[16][27] * mat_B[27][12] +
                  mat_A[16][28] * mat_B[28][12] +
                  mat_A[16][29] * mat_B[29][12] +
                  mat_A[16][30] * mat_B[30][12] +
                  mat_A[16][31] * mat_B[31][12];
    mat_C[16][13] <= 
                  mat_A[16][0] * mat_B[0][13] +
                  mat_A[16][1] * mat_B[1][13] +
                  mat_A[16][2] * mat_B[2][13] +
                  mat_A[16][3] * mat_B[3][13] +
                  mat_A[16][4] * mat_B[4][13] +
                  mat_A[16][5] * mat_B[5][13] +
                  mat_A[16][6] * mat_B[6][13] +
                  mat_A[16][7] * mat_B[7][13] +
                  mat_A[16][8] * mat_B[8][13] +
                  mat_A[16][9] * mat_B[9][13] +
                  mat_A[16][10] * mat_B[10][13] +
                  mat_A[16][11] * mat_B[11][13] +
                  mat_A[16][12] * mat_B[12][13] +
                  mat_A[16][13] * mat_B[13][13] +
                  mat_A[16][14] * mat_B[14][13] +
                  mat_A[16][15] * mat_B[15][13] +
                  mat_A[16][16] * mat_B[16][13] +
                  mat_A[16][17] * mat_B[17][13] +
                  mat_A[16][18] * mat_B[18][13] +
                  mat_A[16][19] * mat_B[19][13] +
                  mat_A[16][20] * mat_B[20][13] +
                  mat_A[16][21] * mat_B[21][13] +
                  mat_A[16][22] * mat_B[22][13] +
                  mat_A[16][23] * mat_B[23][13] +
                  mat_A[16][24] * mat_B[24][13] +
                  mat_A[16][25] * mat_B[25][13] +
                  mat_A[16][26] * mat_B[26][13] +
                  mat_A[16][27] * mat_B[27][13] +
                  mat_A[16][28] * mat_B[28][13] +
                  mat_A[16][29] * mat_B[29][13] +
                  mat_A[16][30] * mat_B[30][13] +
                  mat_A[16][31] * mat_B[31][13];
    mat_C[16][14] <= 
                  mat_A[16][0] * mat_B[0][14] +
                  mat_A[16][1] * mat_B[1][14] +
                  mat_A[16][2] * mat_B[2][14] +
                  mat_A[16][3] * mat_B[3][14] +
                  mat_A[16][4] * mat_B[4][14] +
                  mat_A[16][5] * mat_B[5][14] +
                  mat_A[16][6] * mat_B[6][14] +
                  mat_A[16][7] * mat_B[7][14] +
                  mat_A[16][8] * mat_B[8][14] +
                  mat_A[16][9] * mat_B[9][14] +
                  mat_A[16][10] * mat_B[10][14] +
                  mat_A[16][11] * mat_B[11][14] +
                  mat_A[16][12] * mat_B[12][14] +
                  mat_A[16][13] * mat_B[13][14] +
                  mat_A[16][14] * mat_B[14][14] +
                  mat_A[16][15] * mat_B[15][14] +
                  mat_A[16][16] * mat_B[16][14] +
                  mat_A[16][17] * mat_B[17][14] +
                  mat_A[16][18] * mat_B[18][14] +
                  mat_A[16][19] * mat_B[19][14] +
                  mat_A[16][20] * mat_B[20][14] +
                  mat_A[16][21] * mat_B[21][14] +
                  mat_A[16][22] * mat_B[22][14] +
                  mat_A[16][23] * mat_B[23][14] +
                  mat_A[16][24] * mat_B[24][14] +
                  mat_A[16][25] * mat_B[25][14] +
                  mat_A[16][26] * mat_B[26][14] +
                  mat_A[16][27] * mat_B[27][14] +
                  mat_A[16][28] * mat_B[28][14] +
                  mat_A[16][29] * mat_B[29][14] +
                  mat_A[16][30] * mat_B[30][14] +
                  mat_A[16][31] * mat_B[31][14];
    mat_C[16][15] <= 
                  mat_A[16][0] * mat_B[0][15] +
                  mat_A[16][1] * mat_B[1][15] +
                  mat_A[16][2] * mat_B[2][15] +
                  mat_A[16][3] * mat_B[3][15] +
                  mat_A[16][4] * mat_B[4][15] +
                  mat_A[16][5] * mat_B[5][15] +
                  mat_A[16][6] * mat_B[6][15] +
                  mat_A[16][7] * mat_B[7][15] +
                  mat_A[16][8] * mat_B[8][15] +
                  mat_A[16][9] * mat_B[9][15] +
                  mat_A[16][10] * mat_B[10][15] +
                  mat_A[16][11] * mat_B[11][15] +
                  mat_A[16][12] * mat_B[12][15] +
                  mat_A[16][13] * mat_B[13][15] +
                  mat_A[16][14] * mat_B[14][15] +
                  mat_A[16][15] * mat_B[15][15] +
                  mat_A[16][16] * mat_B[16][15] +
                  mat_A[16][17] * mat_B[17][15] +
                  mat_A[16][18] * mat_B[18][15] +
                  mat_A[16][19] * mat_B[19][15] +
                  mat_A[16][20] * mat_B[20][15] +
                  mat_A[16][21] * mat_B[21][15] +
                  mat_A[16][22] * mat_B[22][15] +
                  mat_A[16][23] * mat_B[23][15] +
                  mat_A[16][24] * mat_B[24][15] +
                  mat_A[16][25] * mat_B[25][15] +
                  mat_A[16][26] * mat_B[26][15] +
                  mat_A[16][27] * mat_B[27][15] +
                  mat_A[16][28] * mat_B[28][15] +
                  mat_A[16][29] * mat_B[29][15] +
                  mat_A[16][30] * mat_B[30][15] +
                  mat_A[16][31] * mat_B[31][15];
    mat_C[16][16] <= 
                  mat_A[16][0] * mat_B[0][16] +
                  mat_A[16][1] * mat_B[1][16] +
                  mat_A[16][2] * mat_B[2][16] +
                  mat_A[16][3] * mat_B[3][16] +
                  mat_A[16][4] * mat_B[4][16] +
                  mat_A[16][5] * mat_B[5][16] +
                  mat_A[16][6] * mat_B[6][16] +
                  mat_A[16][7] * mat_B[7][16] +
                  mat_A[16][8] * mat_B[8][16] +
                  mat_A[16][9] * mat_B[9][16] +
                  mat_A[16][10] * mat_B[10][16] +
                  mat_A[16][11] * mat_B[11][16] +
                  mat_A[16][12] * mat_B[12][16] +
                  mat_A[16][13] * mat_B[13][16] +
                  mat_A[16][14] * mat_B[14][16] +
                  mat_A[16][15] * mat_B[15][16] +
                  mat_A[16][16] * mat_B[16][16] +
                  mat_A[16][17] * mat_B[17][16] +
                  mat_A[16][18] * mat_B[18][16] +
                  mat_A[16][19] * mat_B[19][16] +
                  mat_A[16][20] * mat_B[20][16] +
                  mat_A[16][21] * mat_B[21][16] +
                  mat_A[16][22] * mat_B[22][16] +
                  mat_A[16][23] * mat_B[23][16] +
                  mat_A[16][24] * mat_B[24][16] +
                  mat_A[16][25] * mat_B[25][16] +
                  mat_A[16][26] * mat_B[26][16] +
                  mat_A[16][27] * mat_B[27][16] +
                  mat_A[16][28] * mat_B[28][16] +
                  mat_A[16][29] * mat_B[29][16] +
                  mat_A[16][30] * mat_B[30][16] +
                  mat_A[16][31] * mat_B[31][16];
    mat_C[16][17] <= 
                  mat_A[16][0] * mat_B[0][17] +
                  mat_A[16][1] * mat_B[1][17] +
                  mat_A[16][2] * mat_B[2][17] +
                  mat_A[16][3] * mat_B[3][17] +
                  mat_A[16][4] * mat_B[4][17] +
                  mat_A[16][5] * mat_B[5][17] +
                  mat_A[16][6] * mat_B[6][17] +
                  mat_A[16][7] * mat_B[7][17] +
                  mat_A[16][8] * mat_B[8][17] +
                  mat_A[16][9] * mat_B[9][17] +
                  mat_A[16][10] * mat_B[10][17] +
                  mat_A[16][11] * mat_B[11][17] +
                  mat_A[16][12] * mat_B[12][17] +
                  mat_A[16][13] * mat_B[13][17] +
                  mat_A[16][14] * mat_B[14][17] +
                  mat_A[16][15] * mat_B[15][17] +
                  mat_A[16][16] * mat_B[16][17] +
                  mat_A[16][17] * mat_B[17][17] +
                  mat_A[16][18] * mat_B[18][17] +
                  mat_A[16][19] * mat_B[19][17] +
                  mat_A[16][20] * mat_B[20][17] +
                  mat_A[16][21] * mat_B[21][17] +
                  mat_A[16][22] * mat_B[22][17] +
                  mat_A[16][23] * mat_B[23][17] +
                  mat_A[16][24] * mat_B[24][17] +
                  mat_A[16][25] * mat_B[25][17] +
                  mat_A[16][26] * mat_B[26][17] +
                  mat_A[16][27] * mat_B[27][17] +
                  mat_A[16][28] * mat_B[28][17] +
                  mat_A[16][29] * mat_B[29][17] +
                  mat_A[16][30] * mat_B[30][17] +
                  mat_A[16][31] * mat_B[31][17];
    mat_C[16][18] <= 
                  mat_A[16][0] * mat_B[0][18] +
                  mat_A[16][1] * mat_B[1][18] +
                  mat_A[16][2] * mat_B[2][18] +
                  mat_A[16][3] * mat_B[3][18] +
                  mat_A[16][4] * mat_B[4][18] +
                  mat_A[16][5] * mat_B[5][18] +
                  mat_A[16][6] * mat_B[6][18] +
                  mat_A[16][7] * mat_B[7][18] +
                  mat_A[16][8] * mat_B[8][18] +
                  mat_A[16][9] * mat_B[9][18] +
                  mat_A[16][10] * mat_B[10][18] +
                  mat_A[16][11] * mat_B[11][18] +
                  mat_A[16][12] * mat_B[12][18] +
                  mat_A[16][13] * mat_B[13][18] +
                  mat_A[16][14] * mat_B[14][18] +
                  mat_A[16][15] * mat_B[15][18] +
                  mat_A[16][16] * mat_B[16][18] +
                  mat_A[16][17] * mat_B[17][18] +
                  mat_A[16][18] * mat_B[18][18] +
                  mat_A[16][19] * mat_B[19][18] +
                  mat_A[16][20] * mat_B[20][18] +
                  mat_A[16][21] * mat_B[21][18] +
                  mat_A[16][22] * mat_B[22][18] +
                  mat_A[16][23] * mat_B[23][18] +
                  mat_A[16][24] * mat_B[24][18] +
                  mat_A[16][25] * mat_B[25][18] +
                  mat_A[16][26] * mat_B[26][18] +
                  mat_A[16][27] * mat_B[27][18] +
                  mat_A[16][28] * mat_B[28][18] +
                  mat_A[16][29] * mat_B[29][18] +
                  mat_A[16][30] * mat_B[30][18] +
                  mat_A[16][31] * mat_B[31][18];
    mat_C[16][19] <= 
                  mat_A[16][0] * mat_B[0][19] +
                  mat_A[16][1] * mat_B[1][19] +
                  mat_A[16][2] * mat_B[2][19] +
                  mat_A[16][3] * mat_B[3][19] +
                  mat_A[16][4] * mat_B[4][19] +
                  mat_A[16][5] * mat_B[5][19] +
                  mat_A[16][6] * mat_B[6][19] +
                  mat_A[16][7] * mat_B[7][19] +
                  mat_A[16][8] * mat_B[8][19] +
                  mat_A[16][9] * mat_B[9][19] +
                  mat_A[16][10] * mat_B[10][19] +
                  mat_A[16][11] * mat_B[11][19] +
                  mat_A[16][12] * mat_B[12][19] +
                  mat_A[16][13] * mat_B[13][19] +
                  mat_A[16][14] * mat_B[14][19] +
                  mat_A[16][15] * mat_B[15][19] +
                  mat_A[16][16] * mat_B[16][19] +
                  mat_A[16][17] * mat_B[17][19] +
                  mat_A[16][18] * mat_B[18][19] +
                  mat_A[16][19] * mat_B[19][19] +
                  mat_A[16][20] * mat_B[20][19] +
                  mat_A[16][21] * mat_B[21][19] +
                  mat_A[16][22] * mat_B[22][19] +
                  mat_A[16][23] * mat_B[23][19] +
                  mat_A[16][24] * mat_B[24][19] +
                  mat_A[16][25] * mat_B[25][19] +
                  mat_A[16][26] * mat_B[26][19] +
                  mat_A[16][27] * mat_B[27][19] +
                  mat_A[16][28] * mat_B[28][19] +
                  mat_A[16][29] * mat_B[29][19] +
                  mat_A[16][30] * mat_B[30][19] +
                  mat_A[16][31] * mat_B[31][19];
    mat_C[16][20] <= 
                  mat_A[16][0] * mat_B[0][20] +
                  mat_A[16][1] * mat_B[1][20] +
                  mat_A[16][2] * mat_B[2][20] +
                  mat_A[16][3] * mat_B[3][20] +
                  mat_A[16][4] * mat_B[4][20] +
                  mat_A[16][5] * mat_B[5][20] +
                  mat_A[16][6] * mat_B[6][20] +
                  mat_A[16][7] * mat_B[7][20] +
                  mat_A[16][8] * mat_B[8][20] +
                  mat_A[16][9] * mat_B[9][20] +
                  mat_A[16][10] * mat_B[10][20] +
                  mat_A[16][11] * mat_B[11][20] +
                  mat_A[16][12] * mat_B[12][20] +
                  mat_A[16][13] * mat_B[13][20] +
                  mat_A[16][14] * mat_B[14][20] +
                  mat_A[16][15] * mat_B[15][20] +
                  mat_A[16][16] * mat_B[16][20] +
                  mat_A[16][17] * mat_B[17][20] +
                  mat_A[16][18] * mat_B[18][20] +
                  mat_A[16][19] * mat_B[19][20] +
                  mat_A[16][20] * mat_B[20][20] +
                  mat_A[16][21] * mat_B[21][20] +
                  mat_A[16][22] * mat_B[22][20] +
                  mat_A[16][23] * mat_B[23][20] +
                  mat_A[16][24] * mat_B[24][20] +
                  mat_A[16][25] * mat_B[25][20] +
                  mat_A[16][26] * mat_B[26][20] +
                  mat_A[16][27] * mat_B[27][20] +
                  mat_A[16][28] * mat_B[28][20] +
                  mat_A[16][29] * mat_B[29][20] +
                  mat_A[16][30] * mat_B[30][20] +
                  mat_A[16][31] * mat_B[31][20];
    mat_C[16][21] <= 
                  mat_A[16][0] * mat_B[0][21] +
                  mat_A[16][1] * mat_B[1][21] +
                  mat_A[16][2] * mat_B[2][21] +
                  mat_A[16][3] * mat_B[3][21] +
                  mat_A[16][4] * mat_B[4][21] +
                  mat_A[16][5] * mat_B[5][21] +
                  mat_A[16][6] * mat_B[6][21] +
                  mat_A[16][7] * mat_B[7][21] +
                  mat_A[16][8] * mat_B[8][21] +
                  mat_A[16][9] * mat_B[9][21] +
                  mat_A[16][10] * mat_B[10][21] +
                  mat_A[16][11] * mat_B[11][21] +
                  mat_A[16][12] * mat_B[12][21] +
                  mat_A[16][13] * mat_B[13][21] +
                  mat_A[16][14] * mat_B[14][21] +
                  mat_A[16][15] * mat_B[15][21] +
                  mat_A[16][16] * mat_B[16][21] +
                  mat_A[16][17] * mat_B[17][21] +
                  mat_A[16][18] * mat_B[18][21] +
                  mat_A[16][19] * mat_B[19][21] +
                  mat_A[16][20] * mat_B[20][21] +
                  mat_A[16][21] * mat_B[21][21] +
                  mat_A[16][22] * mat_B[22][21] +
                  mat_A[16][23] * mat_B[23][21] +
                  mat_A[16][24] * mat_B[24][21] +
                  mat_A[16][25] * mat_B[25][21] +
                  mat_A[16][26] * mat_B[26][21] +
                  mat_A[16][27] * mat_B[27][21] +
                  mat_A[16][28] * mat_B[28][21] +
                  mat_A[16][29] * mat_B[29][21] +
                  mat_A[16][30] * mat_B[30][21] +
                  mat_A[16][31] * mat_B[31][21];
    mat_C[16][22] <= 
                  mat_A[16][0] * mat_B[0][22] +
                  mat_A[16][1] * mat_B[1][22] +
                  mat_A[16][2] * mat_B[2][22] +
                  mat_A[16][3] * mat_B[3][22] +
                  mat_A[16][4] * mat_B[4][22] +
                  mat_A[16][5] * mat_B[5][22] +
                  mat_A[16][6] * mat_B[6][22] +
                  mat_A[16][7] * mat_B[7][22] +
                  mat_A[16][8] * mat_B[8][22] +
                  mat_A[16][9] * mat_B[9][22] +
                  mat_A[16][10] * mat_B[10][22] +
                  mat_A[16][11] * mat_B[11][22] +
                  mat_A[16][12] * mat_B[12][22] +
                  mat_A[16][13] * mat_B[13][22] +
                  mat_A[16][14] * mat_B[14][22] +
                  mat_A[16][15] * mat_B[15][22] +
                  mat_A[16][16] * mat_B[16][22] +
                  mat_A[16][17] * mat_B[17][22] +
                  mat_A[16][18] * mat_B[18][22] +
                  mat_A[16][19] * mat_B[19][22] +
                  mat_A[16][20] * mat_B[20][22] +
                  mat_A[16][21] * mat_B[21][22] +
                  mat_A[16][22] * mat_B[22][22] +
                  mat_A[16][23] * mat_B[23][22] +
                  mat_A[16][24] * mat_B[24][22] +
                  mat_A[16][25] * mat_B[25][22] +
                  mat_A[16][26] * mat_B[26][22] +
                  mat_A[16][27] * mat_B[27][22] +
                  mat_A[16][28] * mat_B[28][22] +
                  mat_A[16][29] * mat_B[29][22] +
                  mat_A[16][30] * mat_B[30][22] +
                  mat_A[16][31] * mat_B[31][22];
    mat_C[16][23] <= 
                  mat_A[16][0] * mat_B[0][23] +
                  mat_A[16][1] * mat_B[1][23] +
                  mat_A[16][2] * mat_B[2][23] +
                  mat_A[16][3] * mat_B[3][23] +
                  mat_A[16][4] * mat_B[4][23] +
                  mat_A[16][5] * mat_B[5][23] +
                  mat_A[16][6] * mat_B[6][23] +
                  mat_A[16][7] * mat_B[7][23] +
                  mat_A[16][8] * mat_B[8][23] +
                  mat_A[16][9] * mat_B[9][23] +
                  mat_A[16][10] * mat_B[10][23] +
                  mat_A[16][11] * mat_B[11][23] +
                  mat_A[16][12] * mat_B[12][23] +
                  mat_A[16][13] * mat_B[13][23] +
                  mat_A[16][14] * mat_B[14][23] +
                  mat_A[16][15] * mat_B[15][23] +
                  mat_A[16][16] * mat_B[16][23] +
                  mat_A[16][17] * mat_B[17][23] +
                  mat_A[16][18] * mat_B[18][23] +
                  mat_A[16][19] * mat_B[19][23] +
                  mat_A[16][20] * mat_B[20][23] +
                  mat_A[16][21] * mat_B[21][23] +
                  mat_A[16][22] * mat_B[22][23] +
                  mat_A[16][23] * mat_B[23][23] +
                  mat_A[16][24] * mat_B[24][23] +
                  mat_A[16][25] * mat_B[25][23] +
                  mat_A[16][26] * mat_B[26][23] +
                  mat_A[16][27] * mat_B[27][23] +
                  mat_A[16][28] * mat_B[28][23] +
                  mat_A[16][29] * mat_B[29][23] +
                  mat_A[16][30] * mat_B[30][23] +
                  mat_A[16][31] * mat_B[31][23];
    mat_C[16][24] <= 
                  mat_A[16][0] * mat_B[0][24] +
                  mat_A[16][1] * mat_B[1][24] +
                  mat_A[16][2] * mat_B[2][24] +
                  mat_A[16][3] * mat_B[3][24] +
                  mat_A[16][4] * mat_B[4][24] +
                  mat_A[16][5] * mat_B[5][24] +
                  mat_A[16][6] * mat_B[6][24] +
                  mat_A[16][7] * mat_B[7][24] +
                  mat_A[16][8] * mat_B[8][24] +
                  mat_A[16][9] * mat_B[9][24] +
                  mat_A[16][10] * mat_B[10][24] +
                  mat_A[16][11] * mat_B[11][24] +
                  mat_A[16][12] * mat_B[12][24] +
                  mat_A[16][13] * mat_B[13][24] +
                  mat_A[16][14] * mat_B[14][24] +
                  mat_A[16][15] * mat_B[15][24] +
                  mat_A[16][16] * mat_B[16][24] +
                  mat_A[16][17] * mat_B[17][24] +
                  mat_A[16][18] * mat_B[18][24] +
                  mat_A[16][19] * mat_B[19][24] +
                  mat_A[16][20] * mat_B[20][24] +
                  mat_A[16][21] * mat_B[21][24] +
                  mat_A[16][22] * mat_B[22][24] +
                  mat_A[16][23] * mat_B[23][24] +
                  mat_A[16][24] * mat_B[24][24] +
                  mat_A[16][25] * mat_B[25][24] +
                  mat_A[16][26] * mat_B[26][24] +
                  mat_A[16][27] * mat_B[27][24] +
                  mat_A[16][28] * mat_B[28][24] +
                  mat_A[16][29] * mat_B[29][24] +
                  mat_A[16][30] * mat_B[30][24] +
                  mat_A[16][31] * mat_B[31][24];
    mat_C[16][25] <= 
                  mat_A[16][0] * mat_B[0][25] +
                  mat_A[16][1] * mat_B[1][25] +
                  mat_A[16][2] * mat_B[2][25] +
                  mat_A[16][3] * mat_B[3][25] +
                  mat_A[16][4] * mat_B[4][25] +
                  mat_A[16][5] * mat_B[5][25] +
                  mat_A[16][6] * mat_B[6][25] +
                  mat_A[16][7] * mat_B[7][25] +
                  mat_A[16][8] * mat_B[8][25] +
                  mat_A[16][9] * mat_B[9][25] +
                  mat_A[16][10] * mat_B[10][25] +
                  mat_A[16][11] * mat_B[11][25] +
                  mat_A[16][12] * mat_B[12][25] +
                  mat_A[16][13] * mat_B[13][25] +
                  mat_A[16][14] * mat_B[14][25] +
                  mat_A[16][15] * mat_B[15][25] +
                  mat_A[16][16] * mat_B[16][25] +
                  mat_A[16][17] * mat_B[17][25] +
                  mat_A[16][18] * mat_B[18][25] +
                  mat_A[16][19] * mat_B[19][25] +
                  mat_A[16][20] * mat_B[20][25] +
                  mat_A[16][21] * mat_B[21][25] +
                  mat_A[16][22] * mat_B[22][25] +
                  mat_A[16][23] * mat_B[23][25] +
                  mat_A[16][24] * mat_B[24][25] +
                  mat_A[16][25] * mat_B[25][25] +
                  mat_A[16][26] * mat_B[26][25] +
                  mat_A[16][27] * mat_B[27][25] +
                  mat_A[16][28] * mat_B[28][25] +
                  mat_A[16][29] * mat_B[29][25] +
                  mat_A[16][30] * mat_B[30][25] +
                  mat_A[16][31] * mat_B[31][25];
    mat_C[16][26] <= 
                  mat_A[16][0] * mat_B[0][26] +
                  mat_A[16][1] * mat_B[1][26] +
                  mat_A[16][2] * mat_B[2][26] +
                  mat_A[16][3] * mat_B[3][26] +
                  mat_A[16][4] * mat_B[4][26] +
                  mat_A[16][5] * mat_B[5][26] +
                  mat_A[16][6] * mat_B[6][26] +
                  mat_A[16][7] * mat_B[7][26] +
                  mat_A[16][8] * mat_B[8][26] +
                  mat_A[16][9] * mat_B[9][26] +
                  mat_A[16][10] * mat_B[10][26] +
                  mat_A[16][11] * mat_B[11][26] +
                  mat_A[16][12] * mat_B[12][26] +
                  mat_A[16][13] * mat_B[13][26] +
                  mat_A[16][14] * mat_B[14][26] +
                  mat_A[16][15] * mat_B[15][26] +
                  mat_A[16][16] * mat_B[16][26] +
                  mat_A[16][17] * mat_B[17][26] +
                  mat_A[16][18] * mat_B[18][26] +
                  mat_A[16][19] * mat_B[19][26] +
                  mat_A[16][20] * mat_B[20][26] +
                  mat_A[16][21] * mat_B[21][26] +
                  mat_A[16][22] * mat_B[22][26] +
                  mat_A[16][23] * mat_B[23][26] +
                  mat_A[16][24] * mat_B[24][26] +
                  mat_A[16][25] * mat_B[25][26] +
                  mat_A[16][26] * mat_B[26][26] +
                  mat_A[16][27] * mat_B[27][26] +
                  mat_A[16][28] * mat_B[28][26] +
                  mat_A[16][29] * mat_B[29][26] +
                  mat_A[16][30] * mat_B[30][26] +
                  mat_A[16][31] * mat_B[31][26];
    mat_C[16][27] <= 
                  mat_A[16][0] * mat_B[0][27] +
                  mat_A[16][1] * mat_B[1][27] +
                  mat_A[16][2] * mat_B[2][27] +
                  mat_A[16][3] * mat_B[3][27] +
                  mat_A[16][4] * mat_B[4][27] +
                  mat_A[16][5] * mat_B[5][27] +
                  mat_A[16][6] * mat_B[6][27] +
                  mat_A[16][7] * mat_B[7][27] +
                  mat_A[16][8] * mat_B[8][27] +
                  mat_A[16][9] * mat_B[9][27] +
                  mat_A[16][10] * mat_B[10][27] +
                  mat_A[16][11] * mat_B[11][27] +
                  mat_A[16][12] * mat_B[12][27] +
                  mat_A[16][13] * mat_B[13][27] +
                  mat_A[16][14] * mat_B[14][27] +
                  mat_A[16][15] * mat_B[15][27] +
                  mat_A[16][16] * mat_B[16][27] +
                  mat_A[16][17] * mat_B[17][27] +
                  mat_A[16][18] * mat_B[18][27] +
                  mat_A[16][19] * mat_B[19][27] +
                  mat_A[16][20] * mat_B[20][27] +
                  mat_A[16][21] * mat_B[21][27] +
                  mat_A[16][22] * mat_B[22][27] +
                  mat_A[16][23] * mat_B[23][27] +
                  mat_A[16][24] * mat_B[24][27] +
                  mat_A[16][25] * mat_B[25][27] +
                  mat_A[16][26] * mat_B[26][27] +
                  mat_A[16][27] * mat_B[27][27] +
                  mat_A[16][28] * mat_B[28][27] +
                  mat_A[16][29] * mat_B[29][27] +
                  mat_A[16][30] * mat_B[30][27] +
                  mat_A[16][31] * mat_B[31][27];
    mat_C[16][28] <= 
                  mat_A[16][0] * mat_B[0][28] +
                  mat_A[16][1] * mat_B[1][28] +
                  mat_A[16][2] * mat_B[2][28] +
                  mat_A[16][3] * mat_B[3][28] +
                  mat_A[16][4] * mat_B[4][28] +
                  mat_A[16][5] * mat_B[5][28] +
                  mat_A[16][6] * mat_B[6][28] +
                  mat_A[16][7] * mat_B[7][28] +
                  mat_A[16][8] * mat_B[8][28] +
                  mat_A[16][9] * mat_B[9][28] +
                  mat_A[16][10] * mat_B[10][28] +
                  mat_A[16][11] * mat_B[11][28] +
                  mat_A[16][12] * mat_B[12][28] +
                  mat_A[16][13] * mat_B[13][28] +
                  mat_A[16][14] * mat_B[14][28] +
                  mat_A[16][15] * mat_B[15][28] +
                  mat_A[16][16] * mat_B[16][28] +
                  mat_A[16][17] * mat_B[17][28] +
                  mat_A[16][18] * mat_B[18][28] +
                  mat_A[16][19] * mat_B[19][28] +
                  mat_A[16][20] * mat_B[20][28] +
                  mat_A[16][21] * mat_B[21][28] +
                  mat_A[16][22] * mat_B[22][28] +
                  mat_A[16][23] * mat_B[23][28] +
                  mat_A[16][24] * mat_B[24][28] +
                  mat_A[16][25] * mat_B[25][28] +
                  mat_A[16][26] * mat_B[26][28] +
                  mat_A[16][27] * mat_B[27][28] +
                  mat_A[16][28] * mat_B[28][28] +
                  mat_A[16][29] * mat_B[29][28] +
                  mat_A[16][30] * mat_B[30][28] +
                  mat_A[16][31] * mat_B[31][28];
    mat_C[16][29] <= 
                  mat_A[16][0] * mat_B[0][29] +
                  mat_A[16][1] * mat_B[1][29] +
                  mat_A[16][2] * mat_B[2][29] +
                  mat_A[16][3] * mat_B[3][29] +
                  mat_A[16][4] * mat_B[4][29] +
                  mat_A[16][5] * mat_B[5][29] +
                  mat_A[16][6] * mat_B[6][29] +
                  mat_A[16][7] * mat_B[7][29] +
                  mat_A[16][8] * mat_B[8][29] +
                  mat_A[16][9] * mat_B[9][29] +
                  mat_A[16][10] * mat_B[10][29] +
                  mat_A[16][11] * mat_B[11][29] +
                  mat_A[16][12] * mat_B[12][29] +
                  mat_A[16][13] * mat_B[13][29] +
                  mat_A[16][14] * mat_B[14][29] +
                  mat_A[16][15] * mat_B[15][29] +
                  mat_A[16][16] * mat_B[16][29] +
                  mat_A[16][17] * mat_B[17][29] +
                  mat_A[16][18] * mat_B[18][29] +
                  mat_A[16][19] * mat_B[19][29] +
                  mat_A[16][20] * mat_B[20][29] +
                  mat_A[16][21] * mat_B[21][29] +
                  mat_A[16][22] * mat_B[22][29] +
                  mat_A[16][23] * mat_B[23][29] +
                  mat_A[16][24] * mat_B[24][29] +
                  mat_A[16][25] * mat_B[25][29] +
                  mat_A[16][26] * mat_B[26][29] +
                  mat_A[16][27] * mat_B[27][29] +
                  mat_A[16][28] * mat_B[28][29] +
                  mat_A[16][29] * mat_B[29][29] +
                  mat_A[16][30] * mat_B[30][29] +
                  mat_A[16][31] * mat_B[31][29];
    mat_C[16][30] <= 
                  mat_A[16][0] * mat_B[0][30] +
                  mat_A[16][1] * mat_B[1][30] +
                  mat_A[16][2] * mat_B[2][30] +
                  mat_A[16][3] * mat_B[3][30] +
                  mat_A[16][4] * mat_B[4][30] +
                  mat_A[16][5] * mat_B[5][30] +
                  mat_A[16][6] * mat_B[6][30] +
                  mat_A[16][7] * mat_B[7][30] +
                  mat_A[16][8] * mat_B[8][30] +
                  mat_A[16][9] * mat_B[9][30] +
                  mat_A[16][10] * mat_B[10][30] +
                  mat_A[16][11] * mat_B[11][30] +
                  mat_A[16][12] * mat_B[12][30] +
                  mat_A[16][13] * mat_B[13][30] +
                  mat_A[16][14] * mat_B[14][30] +
                  mat_A[16][15] * mat_B[15][30] +
                  mat_A[16][16] * mat_B[16][30] +
                  mat_A[16][17] * mat_B[17][30] +
                  mat_A[16][18] * mat_B[18][30] +
                  mat_A[16][19] * mat_B[19][30] +
                  mat_A[16][20] * mat_B[20][30] +
                  mat_A[16][21] * mat_B[21][30] +
                  mat_A[16][22] * mat_B[22][30] +
                  mat_A[16][23] * mat_B[23][30] +
                  mat_A[16][24] * mat_B[24][30] +
                  mat_A[16][25] * mat_B[25][30] +
                  mat_A[16][26] * mat_B[26][30] +
                  mat_A[16][27] * mat_B[27][30] +
                  mat_A[16][28] * mat_B[28][30] +
                  mat_A[16][29] * mat_B[29][30] +
                  mat_A[16][30] * mat_B[30][30] +
                  mat_A[16][31] * mat_B[31][30];
    mat_C[16][31] <= 
                  mat_A[16][0] * mat_B[0][31] +
                  mat_A[16][1] * mat_B[1][31] +
                  mat_A[16][2] * mat_B[2][31] +
                  mat_A[16][3] * mat_B[3][31] +
                  mat_A[16][4] * mat_B[4][31] +
                  mat_A[16][5] * mat_B[5][31] +
                  mat_A[16][6] * mat_B[6][31] +
                  mat_A[16][7] * mat_B[7][31] +
                  mat_A[16][8] * mat_B[8][31] +
                  mat_A[16][9] * mat_B[9][31] +
                  mat_A[16][10] * mat_B[10][31] +
                  mat_A[16][11] * mat_B[11][31] +
                  mat_A[16][12] * mat_B[12][31] +
                  mat_A[16][13] * mat_B[13][31] +
                  mat_A[16][14] * mat_B[14][31] +
                  mat_A[16][15] * mat_B[15][31] +
                  mat_A[16][16] * mat_B[16][31] +
                  mat_A[16][17] * mat_B[17][31] +
                  mat_A[16][18] * mat_B[18][31] +
                  mat_A[16][19] * mat_B[19][31] +
                  mat_A[16][20] * mat_B[20][31] +
                  mat_A[16][21] * mat_B[21][31] +
                  mat_A[16][22] * mat_B[22][31] +
                  mat_A[16][23] * mat_B[23][31] +
                  mat_A[16][24] * mat_B[24][31] +
                  mat_A[16][25] * mat_B[25][31] +
                  mat_A[16][26] * mat_B[26][31] +
                  mat_A[16][27] * mat_B[27][31] +
                  mat_A[16][28] * mat_B[28][31] +
                  mat_A[16][29] * mat_B[29][31] +
                  mat_A[16][30] * mat_B[30][31] +
                  mat_A[16][31] * mat_B[31][31];
    mat_C[17][0] <= 
                  mat_A[17][0] * mat_B[0][0] +
                  mat_A[17][1] * mat_B[1][0] +
                  mat_A[17][2] * mat_B[2][0] +
                  mat_A[17][3] * mat_B[3][0] +
                  mat_A[17][4] * mat_B[4][0] +
                  mat_A[17][5] * mat_B[5][0] +
                  mat_A[17][6] * mat_B[6][0] +
                  mat_A[17][7] * mat_B[7][0] +
                  mat_A[17][8] * mat_B[8][0] +
                  mat_A[17][9] * mat_B[9][0] +
                  mat_A[17][10] * mat_B[10][0] +
                  mat_A[17][11] * mat_B[11][0] +
                  mat_A[17][12] * mat_B[12][0] +
                  mat_A[17][13] * mat_B[13][0] +
                  mat_A[17][14] * mat_B[14][0] +
                  mat_A[17][15] * mat_B[15][0] +
                  mat_A[17][16] * mat_B[16][0] +
                  mat_A[17][17] * mat_B[17][0] +
                  mat_A[17][18] * mat_B[18][0] +
                  mat_A[17][19] * mat_B[19][0] +
                  mat_A[17][20] * mat_B[20][0] +
                  mat_A[17][21] * mat_B[21][0] +
                  mat_A[17][22] * mat_B[22][0] +
                  mat_A[17][23] * mat_B[23][0] +
                  mat_A[17][24] * mat_B[24][0] +
                  mat_A[17][25] * mat_B[25][0] +
                  mat_A[17][26] * mat_B[26][0] +
                  mat_A[17][27] * mat_B[27][0] +
                  mat_A[17][28] * mat_B[28][0] +
                  mat_A[17][29] * mat_B[29][0] +
                  mat_A[17][30] * mat_B[30][0] +
                  mat_A[17][31] * mat_B[31][0];
    mat_C[17][1] <= 
                  mat_A[17][0] * mat_B[0][1] +
                  mat_A[17][1] * mat_B[1][1] +
                  mat_A[17][2] * mat_B[2][1] +
                  mat_A[17][3] * mat_B[3][1] +
                  mat_A[17][4] * mat_B[4][1] +
                  mat_A[17][5] * mat_B[5][1] +
                  mat_A[17][6] * mat_B[6][1] +
                  mat_A[17][7] * mat_B[7][1] +
                  mat_A[17][8] * mat_B[8][1] +
                  mat_A[17][9] * mat_B[9][1] +
                  mat_A[17][10] * mat_B[10][1] +
                  mat_A[17][11] * mat_B[11][1] +
                  mat_A[17][12] * mat_B[12][1] +
                  mat_A[17][13] * mat_B[13][1] +
                  mat_A[17][14] * mat_B[14][1] +
                  mat_A[17][15] * mat_B[15][1] +
                  mat_A[17][16] * mat_B[16][1] +
                  mat_A[17][17] * mat_B[17][1] +
                  mat_A[17][18] * mat_B[18][1] +
                  mat_A[17][19] * mat_B[19][1] +
                  mat_A[17][20] * mat_B[20][1] +
                  mat_A[17][21] * mat_B[21][1] +
                  mat_A[17][22] * mat_B[22][1] +
                  mat_A[17][23] * mat_B[23][1] +
                  mat_A[17][24] * mat_B[24][1] +
                  mat_A[17][25] * mat_B[25][1] +
                  mat_A[17][26] * mat_B[26][1] +
                  mat_A[17][27] * mat_B[27][1] +
                  mat_A[17][28] * mat_B[28][1] +
                  mat_A[17][29] * mat_B[29][1] +
                  mat_A[17][30] * mat_B[30][1] +
                  mat_A[17][31] * mat_B[31][1];
    mat_C[17][2] <= 
                  mat_A[17][0] * mat_B[0][2] +
                  mat_A[17][1] * mat_B[1][2] +
                  mat_A[17][2] * mat_B[2][2] +
                  mat_A[17][3] * mat_B[3][2] +
                  mat_A[17][4] * mat_B[4][2] +
                  mat_A[17][5] * mat_B[5][2] +
                  mat_A[17][6] * mat_B[6][2] +
                  mat_A[17][7] * mat_B[7][2] +
                  mat_A[17][8] * mat_B[8][2] +
                  mat_A[17][9] * mat_B[9][2] +
                  mat_A[17][10] * mat_B[10][2] +
                  mat_A[17][11] * mat_B[11][2] +
                  mat_A[17][12] * mat_B[12][2] +
                  mat_A[17][13] * mat_B[13][2] +
                  mat_A[17][14] * mat_B[14][2] +
                  mat_A[17][15] * mat_B[15][2] +
                  mat_A[17][16] * mat_B[16][2] +
                  mat_A[17][17] * mat_B[17][2] +
                  mat_A[17][18] * mat_B[18][2] +
                  mat_A[17][19] * mat_B[19][2] +
                  mat_A[17][20] * mat_B[20][2] +
                  mat_A[17][21] * mat_B[21][2] +
                  mat_A[17][22] * mat_B[22][2] +
                  mat_A[17][23] * mat_B[23][2] +
                  mat_A[17][24] * mat_B[24][2] +
                  mat_A[17][25] * mat_B[25][2] +
                  mat_A[17][26] * mat_B[26][2] +
                  mat_A[17][27] * mat_B[27][2] +
                  mat_A[17][28] * mat_B[28][2] +
                  mat_A[17][29] * mat_B[29][2] +
                  mat_A[17][30] * mat_B[30][2] +
                  mat_A[17][31] * mat_B[31][2];
    mat_C[17][3] <= 
                  mat_A[17][0] * mat_B[0][3] +
                  mat_A[17][1] * mat_B[1][3] +
                  mat_A[17][2] * mat_B[2][3] +
                  mat_A[17][3] * mat_B[3][3] +
                  mat_A[17][4] * mat_B[4][3] +
                  mat_A[17][5] * mat_B[5][3] +
                  mat_A[17][6] * mat_B[6][3] +
                  mat_A[17][7] * mat_B[7][3] +
                  mat_A[17][8] * mat_B[8][3] +
                  mat_A[17][9] * mat_B[9][3] +
                  mat_A[17][10] * mat_B[10][3] +
                  mat_A[17][11] * mat_B[11][3] +
                  mat_A[17][12] * mat_B[12][3] +
                  mat_A[17][13] * mat_B[13][3] +
                  mat_A[17][14] * mat_B[14][3] +
                  mat_A[17][15] * mat_B[15][3] +
                  mat_A[17][16] * mat_B[16][3] +
                  mat_A[17][17] * mat_B[17][3] +
                  mat_A[17][18] * mat_B[18][3] +
                  mat_A[17][19] * mat_B[19][3] +
                  mat_A[17][20] * mat_B[20][3] +
                  mat_A[17][21] * mat_B[21][3] +
                  mat_A[17][22] * mat_B[22][3] +
                  mat_A[17][23] * mat_B[23][3] +
                  mat_A[17][24] * mat_B[24][3] +
                  mat_A[17][25] * mat_B[25][3] +
                  mat_A[17][26] * mat_B[26][3] +
                  mat_A[17][27] * mat_B[27][3] +
                  mat_A[17][28] * mat_B[28][3] +
                  mat_A[17][29] * mat_B[29][3] +
                  mat_A[17][30] * mat_B[30][3] +
                  mat_A[17][31] * mat_B[31][3];
    mat_C[17][4] <= 
                  mat_A[17][0] * mat_B[0][4] +
                  mat_A[17][1] * mat_B[1][4] +
                  mat_A[17][2] * mat_B[2][4] +
                  mat_A[17][3] * mat_B[3][4] +
                  mat_A[17][4] * mat_B[4][4] +
                  mat_A[17][5] * mat_B[5][4] +
                  mat_A[17][6] * mat_B[6][4] +
                  mat_A[17][7] * mat_B[7][4] +
                  mat_A[17][8] * mat_B[8][4] +
                  mat_A[17][9] * mat_B[9][4] +
                  mat_A[17][10] * mat_B[10][4] +
                  mat_A[17][11] * mat_B[11][4] +
                  mat_A[17][12] * mat_B[12][4] +
                  mat_A[17][13] * mat_B[13][4] +
                  mat_A[17][14] * mat_B[14][4] +
                  mat_A[17][15] * mat_B[15][4] +
                  mat_A[17][16] * mat_B[16][4] +
                  mat_A[17][17] * mat_B[17][4] +
                  mat_A[17][18] * mat_B[18][4] +
                  mat_A[17][19] * mat_B[19][4] +
                  mat_A[17][20] * mat_B[20][4] +
                  mat_A[17][21] * mat_B[21][4] +
                  mat_A[17][22] * mat_B[22][4] +
                  mat_A[17][23] * mat_B[23][4] +
                  mat_A[17][24] * mat_B[24][4] +
                  mat_A[17][25] * mat_B[25][4] +
                  mat_A[17][26] * mat_B[26][4] +
                  mat_A[17][27] * mat_B[27][4] +
                  mat_A[17][28] * mat_B[28][4] +
                  mat_A[17][29] * mat_B[29][4] +
                  mat_A[17][30] * mat_B[30][4] +
                  mat_A[17][31] * mat_B[31][4];
    mat_C[17][5] <= 
                  mat_A[17][0] * mat_B[0][5] +
                  mat_A[17][1] * mat_B[1][5] +
                  mat_A[17][2] * mat_B[2][5] +
                  mat_A[17][3] * mat_B[3][5] +
                  mat_A[17][4] * mat_B[4][5] +
                  mat_A[17][5] * mat_B[5][5] +
                  mat_A[17][6] * mat_B[6][5] +
                  mat_A[17][7] * mat_B[7][5] +
                  mat_A[17][8] * mat_B[8][5] +
                  mat_A[17][9] * mat_B[9][5] +
                  mat_A[17][10] * mat_B[10][5] +
                  mat_A[17][11] * mat_B[11][5] +
                  mat_A[17][12] * mat_B[12][5] +
                  mat_A[17][13] * mat_B[13][5] +
                  mat_A[17][14] * mat_B[14][5] +
                  mat_A[17][15] * mat_B[15][5] +
                  mat_A[17][16] * mat_B[16][5] +
                  mat_A[17][17] * mat_B[17][5] +
                  mat_A[17][18] * mat_B[18][5] +
                  mat_A[17][19] * mat_B[19][5] +
                  mat_A[17][20] * mat_B[20][5] +
                  mat_A[17][21] * mat_B[21][5] +
                  mat_A[17][22] * mat_B[22][5] +
                  mat_A[17][23] * mat_B[23][5] +
                  mat_A[17][24] * mat_B[24][5] +
                  mat_A[17][25] * mat_B[25][5] +
                  mat_A[17][26] * mat_B[26][5] +
                  mat_A[17][27] * mat_B[27][5] +
                  mat_A[17][28] * mat_B[28][5] +
                  mat_A[17][29] * mat_B[29][5] +
                  mat_A[17][30] * mat_B[30][5] +
                  mat_A[17][31] * mat_B[31][5];
    mat_C[17][6] <= 
                  mat_A[17][0] * mat_B[0][6] +
                  mat_A[17][1] * mat_B[1][6] +
                  mat_A[17][2] * mat_B[2][6] +
                  mat_A[17][3] * mat_B[3][6] +
                  mat_A[17][4] * mat_B[4][6] +
                  mat_A[17][5] * mat_B[5][6] +
                  mat_A[17][6] * mat_B[6][6] +
                  mat_A[17][7] * mat_B[7][6] +
                  mat_A[17][8] * mat_B[8][6] +
                  mat_A[17][9] * mat_B[9][6] +
                  mat_A[17][10] * mat_B[10][6] +
                  mat_A[17][11] * mat_B[11][6] +
                  mat_A[17][12] * mat_B[12][6] +
                  mat_A[17][13] * mat_B[13][6] +
                  mat_A[17][14] * mat_B[14][6] +
                  mat_A[17][15] * mat_B[15][6] +
                  mat_A[17][16] * mat_B[16][6] +
                  mat_A[17][17] * mat_B[17][6] +
                  mat_A[17][18] * mat_B[18][6] +
                  mat_A[17][19] * mat_B[19][6] +
                  mat_A[17][20] * mat_B[20][6] +
                  mat_A[17][21] * mat_B[21][6] +
                  mat_A[17][22] * mat_B[22][6] +
                  mat_A[17][23] * mat_B[23][6] +
                  mat_A[17][24] * mat_B[24][6] +
                  mat_A[17][25] * mat_B[25][6] +
                  mat_A[17][26] * mat_B[26][6] +
                  mat_A[17][27] * mat_B[27][6] +
                  mat_A[17][28] * mat_B[28][6] +
                  mat_A[17][29] * mat_B[29][6] +
                  mat_A[17][30] * mat_B[30][6] +
                  mat_A[17][31] * mat_B[31][6];
    mat_C[17][7] <= 
                  mat_A[17][0] * mat_B[0][7] +
                  mat_A[17][1] * mat_B[1][7] +
                  mat_A[17][2] * mat_B[2][7] +
                  mat_A[17][3] * mat_B[3][7] +
                  mat_A[17][4] * mat_B[4][7] +
                  mat_A[17][5] * mat_B[5][7] +
                  mat_A[17][6] * mat_B[6][7] +
                  mat_A[17][7] * mat_B[7][7] +
                  mat_A[17][8] * mat_B[8][7] +
                  mat_A[17][9] * mat_B[9][7] +
                  mat_A[17][10] * mat_B[10][7] +
                  mat_A[17][11] * mat_B[11][7] +
                  mat_A[17][12] * mat_B[12][7] +
                  mat_A[17][13] * mat_B[13][7] +
                  mat_A[17][14] * mat_B[14][7] +
                  mat_A[17][15] * mat_B[15][7] +
                  mat_A[17][16] * mat_B[16][7] +
                  mat_A[17][17] * mat_B[17][7] +
                  mat_A[17][18] * mat_B[18][7] +
                  mat_A[17][19] * mat_B[19][7] +
                  mat_A[17][20] * mat_B[20][7] +
                  mat_A[17][21] * mat_B[21][7] +
                  mat_A[17][22] * mat_B[22][7] +
                  mat_A[17][23] * mat_B[23][7] +
                  mat_A[17][24] * mat_B[24][7] +
                  mat_A[17][25] * mat_B[25][7] +
                  mat_A[17][26] * mat_B[26][7] +
                  mat_A[17][27] * mat_B[27][7] +
                  mat_A[17][28] * mat_B[28][7] +
                  mat_A[17][29] * mat_B[29][7] +
                  mat_A[17][30] * mat_B[30][7] +
                  mat_A[17][31] * mat_B[31][7];
    mat_C[17][8] <= 
                  mat_A[17][0] * mat_B[0][8] +
                  mat_A[17][1] * mat_B[1][8] +
                  mat_A[17][2] * mat_B[2][8] +
                  mat_A[17][3] * mat_B[3][8] +
                  mat_A[17][4] * mat_B[4][8] +
                  mat_A[17][5] * mat_B[5][8] +
                  mat_A[17][6] * mat_B[6][8] +
                  mat_A[17][7] * mat_B[7][8] +
                  mat_A[17][8] * mat_B[8][8] +
                  mat_A[17][9] * mat_B[9][8] +
                  mat_A[17][10] * mat_B[10][8] +
                  mat_A[17][11] * mat_B[11][8] +
                  mat_A[17][12] * mat_B[12][8] +
                  mat_A[17][13] * mat_B[13][8] +
                  mat_A[17][14] * mat_B[14][8] +
                  mat_A[17][15] * mat_B[15][8] +
                  mat_A[17][16] * mat_B[16][8] +
                  mat_A[17][17] * mat_B[17][8] +
                  mat_A[17][18] * mat_B[18][8] +
                  mat_A[17][19] * mat_B[19][8] +
                  mat_A[17][20] * mat_B[20][8] +
                  mat_A[17][21] * mat_B[21][8] +
                  mat_A[17][22] * mat_B[22][8] +
                  mat_A[17][23] * mat_B[23][8] +
                  mat_A[17][24] * mat_B[24][8] +
                  mat_A[17][25] * mat_B[25][8] +
                  mat_A[17][26] * mat_B[26][8] +
                  mat_A[17][27] * mat_B[27][8] +
                  mat_A[17][28] * mat_B[28][8] +
                  mat_A[17][29] * mat_B[29][8] +
                  mat_A[17][30] * mat_B[30][8] +
                  mat_A[17][31] * mat_B[31][8];
    mat_C[17][9] <= 
                  mat_A[17][0] * mat_B[0][9] +
                  mat_A[17][1] * mat_B[1][9] +
                  mat_A[17][2] * mat_B[2][9] +
                  mat_A[17][3] * mat_B[3][9] +
                  mat_A[17][4] * mat_B[4][9] +
                  mat_A[17][5] * mat_B[5][9] +
                  mat_A[17][6] * mat_B[6][9] +
                  mat_A[17][7] * mat_B[7][9] +
                  mat_A[17][8] * mat_B[8][9] +
                  mat_A[17][9] * mat_B[9][9] +
                  mat_A[17][10] * mat_B[10][9] +
                  mat_A[17][11] * mat_B[11][9] +
                  mat_A[17][12] * mat_B[12][9] +
                  mat_A[17][13] * mat_B[13][9] +
                  mat_A[17][14] * mat_B[14][9] +
                  mat_A[17][15] * mat_B[15][9] +
                  mat_A[17][16] * mat_B[16][9] +
                  mat_A[17][17] * mat_B[17][9] +
                  mat_A[17][18] * mat_B[18][9] +
                  mat_A[17][19] * mat_B[19][9] +
                  mat_A[17][20] * mat_B[20][9] +
                  mat_A[17][21] * mat_B[21][9] +
                  mat_A[17][22] * mat_B[22][9] +
                  mat_A[17][23] * mat_B[23][9] +
                  mat_A[17][24] * mat_B[24][9] +
                  mat_A[17][25] * mat_B[25][9] +
                  mat_A[17][26] * mat_B[26][9] +
                  mat_A[17][27] * mat_B[27][9] +
                  mat_A[17][28] * mat_B[28][9] +
                  mat_A[17][29] * mat_B[29][9] +
                  mat_A[17][30] * mat_B[30][9] +
                  mat_A[17][31] * mat_B[31][9];
    mat_C[17][10] <= 
                  mat_A[17][0] * mat_B[0][10] +
                  mat_A[17][1] * mat_B[1][10] +
                  mat_A[17][2] * mat_B[2][10] +
                  mat_A[17][3] * mat_B[3][10] +
                  mat_A[17][4] * mat_B[4][10] +
                  mat_A[17][5] * mat_B[5][10] +
                  mat_A[17][6] * mat_B[6][10] +
                  mat_A[17][7] * mat_B[7][10] +
                  mat_A[17][8] * mat_B[8][10] +
                  mat_A[17][9] * mat_B[9][10] +
                  mat_A[17][10] * mat_B[10][10] +
                  mat_A[17][11] * mat_B[11][10] +
                  mat_A[17][12] * mat_B[12][10] +
                  mat_A[17][13] * mat_B[13][10] +
                  mat_A[17][14] * mat_B[14][10] +
                  mat_A[17][15] * mat_B[15][10] +
                  mat_A[17][16] * mat_B[16][10] +
                  mat_A[17][17] * mat_B[17][10] +
                  mat_A[17][18] * mat_B[18][10] +
                  mat_A[17][19] * mat_B[19][10] +
                  mat_A[17][20] * mat_B[20][10] +
                  mat_A[17][21] * mat_B[21][10] +
                  mat_A[17][22] * mat_B[22][10] +
                  mat_A[17][23] * mat_B[23][10] +
                  mat_A[17][24] * mat_B[24][10] +
                  mat_A[17][25] * mat_B[25][10] +
                  mat_A[17][26] * mat_B[26][10] +
                  mat_A[17][27] * mat_B[27][10] +
                  mat_A[17][28] * mat_B[28][10] +
                  mat_A[17][29] * mat_B[29][10] +
                  mat_A[17][30] * mat_B[30][10] +
                  mat_A[17][31] * mat_B[31][10];
    mat_C[17][11] <= 
                  mat_A[17][0] * mat_B[0][11] +
                  mat_A[17][1] * mat_B[1][11] +
                  mat_A[17][2] * mat_B[2][11] +
                  mat_A[17][3] * mat_B[3][11] +
                  mat_A[17][4] * mat_B[4][11] +
                  mat_A[17][5] * mat_B[5][11] +
                  mat_A[17][6] * mat_B[6][11] +
                  mat_A[17][7] * mat_B[7][11] +
                  mat_A[17][8] * mat_B[8][11] +
                  mat_A[17][9] * mat_B[9][11] +
                  mat_A[17][10] * mat_B[10][11] +
                  mat_A[17][11] * mat_B[11][11] +
                  mat_A[17][12] * mat_B[12][11] +
                  mat_A[17][13] * mat_B[13][11] +
                  mat_A[17][14] * mat_B[14][11] +
                  mat_A[17][15] * mat_B[15][11] +
                  mat_A[17][16] * mat_B[16][11] +
                  mat_A[17][17] * mat_B[17][11] +
                  mat_A[17][18] * mat_B[18][11] +
                  mat_A[17][19] * mat_B[19][11] +
                  mat_A[17][20] * mat_B[20][11] +
                  mat_A[17][21] * mat_B[21][11] +
                  mat_A[17][22] * mat_B[22][11] +
                  mat_A[17][23] * mat_B[23][11] +
                  mat_A[17][24] * mat_B[24][11] +
                  mat_A[17][25] * mat_B[25][11] +
                  mat_A[17][26] * mat_B[26][11] +
                  mat_A[17][27] * mat_B[27][11] +
                  mat_A[17][28] * mat_B[28][11] +
                  mat_A[17][29] * mat_B[29][11] +
                  mat_A[17][30] * mat_B[30][11] +
                  mat_A[17][31] * mat_B[31][11];
    mat_C[17][12] <= 
                  mat_A[17][0] * mat_B[0][12] +
                  mat_A[17][1] * mat_B[1][12] +
                  mat_A[17][2] * mat_B[2][12] +
                  mat_A[17][3] * mat_B[3][12] +
                  mat_A[17][4] * mat_B[4][12] +
                  mat_A[17][5] * mat_B[5][12] +
                  mat_A[17][6] * mat_B[6][12] +
                  mat_A[17][7] * mat_B[7][12] +
                  mat_A[17][8] * mat_B[8][12] +
                  mat_A[17][9] * mat_B[9][12] +
                  mat_A[17][10] * mat_B[10][12] +
                  mat_A[17][11] * mat_B[11][12] +
                  mat_A[17][12] * mat_B[12][12] +
                  mat_A[17][13] * mat_B[13][12] +
                  mat_A[17][14] * mat_B[14][12] +
                  mat_A[17][15] * mat_B[15][12] +
                  mat_A[17][16] * mat_B[16][12] +
                  mat_A[17][17] * mat_B[17][12] +
                  mat_A[17][18] * mat_B[18][12] +
                  mat_A[17][19] * mat_B[19][12] +
                  mat_A[17][20] * mat_B[20][12] +
                  mat_A[17][21] * mat_B[21][12] +
                  mat_A[17][22] * mat_B[22][12] +
                  mat_A[17][23] * mat_B[23][12] +
                  mat_A[17][24] * mat_B[24][12] +
                  mat_A[17][25] * mat_B[25][12] +
                  mat_A[17][26] * mat_B[26][12] +
                  mat_A[17][27] * mat_B[27][12] +
                  mat_A[17][28] * mat_B[28][12] +
                  mat_A[17][29] * mat_B[29][12] +
                  mat_A[17][30] * mat_B[30][12] +
                  mat_A[17][31] * mat_B[31][12];
    mat_C[17][13] <= 
                  mat_A[17][0] * mat_B[0][13] +
                  mat_A[17][1] * mat_B[1][13] +
                  mat_A[17][2] * mat_B[2][13] +
                  mat_A[17][3] * mat_B[3][13] +
                  mat_A[17][4] * mat_B[4][13] +
                  mat_A[17][5] * mat_B[5][13] +
                  mat_A[17][6] * mat_B[6][13] +
                  mat_A[17][7] * mat_B[7][13] +
                  mat_A[17][8] * mat_B[8][13] +
                  mat_A[17][9] * mat_B[9][13] +
                  mat_A[17][10] * mat_B[10][13] +
                  mat_A[17][11] * mat_B[11][13] +
                  mat_A[17][12] * mat_B[12][13] +
                  mat_A[17][13] * mat_B[13][13] +
                  mat_A[17][14] * mat_B[14][13] +
                  mat_A[17][15] * mat_B[15][13] +
                  mat_A[17][16] * mat_B[16][13] +
                  mat_A[17][17] * mat_B[17][13] +
                  mat_A[17][18] * mat_B[18][13] +
                  mat_A[17][19] * mat_B[19][13] +
                  mat_A[17][20] * mat_B[20][13] +
                  mat_A[17][21] * mat_B[21][13] +
                  mat_A[17][22] * mat_B[22][13] +
                  mat_A[17][23] * mat_B[23][13] +
                  mat_A[17][24] * mat_B[24][13] +
                  mat_A[17][25] * mat_B[25][13] +
                  mat_A[17][26] * mat_B[26][13] +
                  mat_A[17][27] * mat_B[27][13] +
                  mat_A[17][28] * mat_B[28][13] +
                  mat_A[17][29] * mat_B[29][13] +
                  mat_A[17][30] * mat_B[30][13] +
                  mat_A[17][31] * mat_B[31][13];
    mat_C[17][14] <= 
                  mat_A[17][0] * mat_B[0][14] +
                  mat_A[17][1] * mat_B[1][14] +
                  mat_A[17][2] * mat_B[2][14] +
                  mat_A[17][3] * mat_B[3][14] +
                  mat_A[17][4] * mat_B[4][14] +
                  mat_A[17][5] * mat_B[5][14] +
                  mat_A[17][6] * mat_B[6][14] +
                  mat_A[17][7] * mat_B[7][14] +
                  mat_A[17][8] * mat_B[8][14] +
                  mat_A[17][9] * mat_B[9][14] +
                  mat_A[17][10] * mat_B[10][14] +
                  mat_A[17][11] * mat_B[11][14] +
                  mat_A[17][12] * mat_B[12][14] +
                  mat_A[17][13] * mat_B[13][14] +
                  mat_A[17][14] * mat_B[14][14] +
                  mat_A[17][15] * mat_B[15][14] +
                  mat_A[17][16] * mat_B[16][14] +
                  mat_A[17][17] * mat_B[17][14] +
                  mat_A[17][18] * mat_B[18][14] +
                  mat_A[17][19] * mat_B[19][14] +
                  mat_A[17][20] * mat_B[20][14] +
                  mat_A[17][21] * mat_B[21][14] +
                  mat_A[17][22] * mat_B[22][14] +
                  mat_A[17][23] * mat_B[23][14] +
                  mat_A[17][24] * mat_B[24][14] +
                  mat_A[17][25] * mat_B[25][14] +
                  mat_A[17][26] * mat_B[26][14] +
                  mat_A[17][27] * mat_B[27][14] +
                  mat_A[17][28] * mat_B[28][14] +
                  mat_A[17][29] * mat_B[29][14] +
                  mat_A[17][30] * mat_B[30][14] +
                  mat_A[17][31] * mat_B[31][14];
    mat_C[17][15] <= 
                  mat_A[17][0] * mat_B[0][15] +
                  mat_A[17][1] * mat_B[1][15] +
                  mat_A[17][2] * mat_B[2][15] +
                  mat_A[17][3] * mat_B[3][15] +
                  mat_A[17][4] * mat_B[4][15] +
                  mat_A[17][5] * mat_B[5][15] +
                  mat_A[17][6] * mat_B[6][15] +
                  mat_A[17][7] * mat_B[7][15] +
                  mat_A[17][8] * mat_B[8][15] +
                  mat_A[17][9] * mat_B[9][15] +
                  mat_A[17][10] * mat_B[10][15] +
                  mat_A[17][11] * mat_B[11][15] +
                  mat_A[17][12] * mat_B[12][15] +
                  mat_A[17][13] * mat_B[13][15] +
                  mat_A[17][14] * mat_B[14][15] +
                  mat_A[17][15] * mat_B[15][15] +
                  mat_A[17][16] * mat_B[16][15] +
                  mat_A[17][17] * mat_B[17][15] +
                  mat_A[17][18] * mat_B[18][15] +
                  mat_A[17][19] * mat_B[19][15] +
                  mat_A[17][20] * mat_B[20][15] +
                  mat_A[17][21] * mat_B[21][15] +
                  mat_A[17][22] * mat_B[22][15] +
                  mat_A[17][23] * mat_B[23][15] +
                  mat_A[17][24] * mat_B[24][15] +
                  mat_A[17][25] * mat_B[25][15] +
                  mat_A[17][26] * mat_B[26][15] +
                  mat_A[17][27] * mat_B[27][15] +
                  mat_A[17][28] * mat_B[28][15] +
                  mat_A[17][29] * mat_B[29][15] +
                  mat_A[17][30] * mat_B[30][15] +
                  mat_A[17][31] * mat_B[31][15];
    mat_C[17][16] <= 
                  mat_A[17][0] * mat_B[0][16] +
                  mat_A[17][1] * mat_B[1][16] +
                  mat_A[17][2] * mat_B[2][16] +
                  mat_A[17][3] * mat_B[3][16] +
                  mat_A[17][4] * mat_B[4][16] +
                  mat_A[17][5] * mat_B[5][16] +
                  mat_A[17][6] * mat_B[6][16] +
                  mat_A[17][7] * mat_B[7][16] +
                  mat_A[17][8] * mat_B[8][16] +
                  mat_A[17][9] * mat_B[9][16] +
                  mat_A[17][10] * mat_B[10][16] +
                  mat_A[17][11] * mat_B[11][16] +
                  mat_A[17][12] * mat_B[12][16] +
                  mat_A[17][13] * mat_B[13][16] +
                  mat_A[17][14] * mat_B[14][16] +
                  mat_A[17][15] * mat_B[15][16] +
                  mat_A[17][16] * mat_B[16][16] +
                  mat_A[17][17] * mat_B[17][16] +
                  mat_A[17][18] * mat_B[18][16] +
                  mat_A[17][19] * mat_B[19][16] +
                  mat_A[17][20] * mat_B[20][16] +
                  mat_A[17][21] * mat_B[21][16] +
                  mat_A[17][22] * mat_B[22][16] +
                  mat_A[17][23] * mat_B[23][16] +
                  mat_A[17][24] * mat_B[24][16] +
                  mat_A[17][25] * mat_B[25][16] +
                  mat_A[17][26] * mat_B[26][16] +
                  mat_A[17][27] * mat_B[27][16] +
                  mat_A[17][28] * mat_B[28][16] +
                  mat_A[17][29] * mat_B[29][16] +
                  mat_A[17][30] * mat_B[30][16] +
                  mat_A[17][31] * mat_B[31][16];
    mat_C[17][17] <= 
                  mat_A[17][0] * mat_B[0][17] +
                  mat_A[17][1] * mat_B[1][17] +
                  mat_A[17][2] * mat_B[2][17] +
                  mat_A[17][3] * mat_B[3][17] +
                  mat_A[17][4] * mat_B[4][17] +
                  mat_A[17][5] * mat_B[5][17] +
                  mat_A[17][6] * mat_B[6][17] +
                  mat_A[17][7] * mat_B[7][17] +
                  mat_A[17][8] * mat_B[8][17] +
                  mat_A[17][9] * mat_B[9][17] +
                  mat_A[17][10] * mat_B[10][17] +
                  mat_A[17][11] * mat_B[11][17] +
                  mat_A[17][12] * mat_B[12][17] +
                  mat_A[17][13] * mat_B[13][17] +
                  mat_A[17][14] * mat_B[14][17] +
                  mat_A[17][15] * mat_B[15][17] +
                  mat_A[17][16] * mat_B[16][17] +
                  mat_A[17][17] * mat_B[17][17] +
                  mat_A[17][18] * mat_B[18][17] +
                  mat_A[17][19] * mat_B[19][17] +
                  mat_A[17][20] * mat_B[20][17] +
                  mat_A[17][21] * mat_B[21][17] +
                  mat_A[17][22] * mat_B[22][17] +
                  mat_A[17][23] * mat_B[23][17] +
                  mat_A[17][24] * mat_B[24][17] +
                  mat_A[17][25] * mat_B[25][17] +
                  mat_A[17][26] * mat_B[26][17] +
                  mat_A[17][27] * mat_B[27][17] +
                  mat_A[17][28] * mat_B[28][17] +
                  mat_A[17][29] * mat_B[29][17] +
                  mat_A[17][30] * mat_B[30][17] +
                  mat_A[17][31] * mat_B[31][17];
    mat_C[17][18] <= 
                  mat_A[17][0] * mat_B[0][18] +
                  mat_A[17][1] * mat_B[1][18] +
                  mat_A[17][2] * mat_B[2][18] +
                  mat_A[17][3] * mat_B[3][18] +
                  mat_A[17][4] * mat_B[4][18] +
                  mat_A[17][5] * mat_B[5][18] +
                  mat_A[17][6] * mat_B[6][18] +
                  mat_A[17][7] * mat_B[7][18] +
                  mat_A[17][8] * mat_B[8][18] +
                  mat_A[17][9] * mat_B[9][18] +
                  mat_A[17][10] * mat_B[10][18] +
                  mat_A[17][11] * mat_B[11][18] +
                  mat_A[17][12] * mat_B[12][18] +
                  mat_A[17][13] * mat_B[13][18] +
                  mat_A[17][14] * mat_B[14][18] +
                  mat_A[17][15] * mat_B[15][18] +
                  mat_A[17][16] * mat_B[16][18] +
                  mat_A[17][17] * mat_B[17][18] +
                  mat_A[17][18] * mat_B[18][18] +
                  mat_A[17][19] * mat_B[19][18] +
                  mat_A[17][20] * mat_B[20][18] +
                  mat_A[17][21] * mat_B[21][18] +
                  mat_A[17][22] * mat_B[22][18] +
                  mat_A[17][23] * mat_B[23][18] +
                  mat_A[17][24] * mat_B[24][18] +
                  mat_A[17][25] * mat_B[25][18] +
                  mat_A[17][26] * mat_B[26][18] +
                  mat_A[17][27] * mat_B[27][18] +
                  mat_A[17][28] * mat_B[28][18] +
                  mat_A[17][29] * mat_B[29][18] +
                  mat_A[17][30] * mat_B[30][18] +
                  mat_A[17][31] * mat_B[31][18];
    mat_C[17][19] <= 
                  mat_A[17][0] * mat_B[0][19] +
                  mat_A[17][1] * mat_B[1][19] +
                  mat_A[17][2] * mat_B[2][19] +
                  mat_A[17][3] * mat_B[3][19] +
                  mat_A[17][4] * mat_B[4][19] +
                  mat_A[17][5] * mat_B[5][19] +
                  mat_A[17][6] * mat_B[6][19] +
                  mat_A[17][7] * mat_B[7][19] +
                  mat_A[17][8] * mat_B[8][19] +
                  mat_A[17][9] * mat_B[9][19] +
                  mat_A[17][10] * mat_B[10][19] +
                  mat_A[17][11] * mat_B[11][19] +
                  mat_A[17][12] * mat_B[12][19] +
                  mat_A[17][13] * mat_B[13][19] +
                  mat_A[17][14] * mat_B[14][19] +
                  mat_A[17][15] * mat_B[15][19] +
                  mat_A[17][16] * mat_B[16][19] +
                  mat_A[17][17] * mat_B[17][19] +
                  mat_A[17][18] * mat_B[18][19] +
                  mat_A[17][19] * mat_B[19][19] +
                  mat_A[17][20] * mat_B[20][19] +
                  mat_A[17][21] * mat_B[21][19] +
                  mat_A[17][22] * mat_B[22][19] +
                  mat_A[17][23] * mat_B[23][19] +
                  mat_A[17][24] * mat_B[24][19] +
                  mat_A[17][25] * mat_B[25][19] +
                  mat_A[17][26] * mat_B[26][19] +
                  mat_A[17][27] * mat_B[27][19] +
                  mat_A[17][28] * mat_B[28][19] +
                  mat_A[17][29] * mat_B[29][19] +
                  mat_A[17][30] * mat_B[30][19] +
                  mat_A[17][31] * mat_B[31][19];
    mat_C[17][20] <= 
                  mat_A[17][0] * mat_B[0][20] +
                  mat_A[17][1] * mat_B[1][20] +
                  mat_A[17][2] * mat_B[2][20] +
                  mat_A[17][3] * mat_B[3][20] +
                  mat_A[17][4] * mat_B[4][20] +
                  mat_A[17][5] * mat_B[5][20] +
                  mat_A[17][6] * mat_B[6][20] +
                  mat_A[17][7] * mat_B[7][20] +
                  mat_A[17][8] * mat_B[8][20] +
                  mat_A[17][9] * mat_B[9][20] +
                  mat_A[17][10] * mat_B[10][20] +
                  mat_A[17][11] * mat_B[11][20] +
                  mat_A[17][12] * mat_B[12][20] +
                  mat_A[17][13] * mat_B[13][20] +
                  mat_A[17][14] * mat_B[14][20] +
                  mat_A[17][15] * mat_B[15][20] +
                  mat_A[17][16] * mat_B[16][20] +
                  mat_A[17][17] * mat_B[17][20] +
                  mat_A[17][18] * mat_B[18][20] +
                  mat_A[17][19] * mat_B[19][20] +
                  mat_A[17][20] * mat_B[20][20] +
                  mat_A[17][21] * mat_B[21][20] +
                  mat_A[17][22] * mat_B[22][20] +
                  mat_A[17][23] * mat_B[23][20] +
                  mat_A[17][24] * mat_B[24][20] +
                  mat_A[17][25] * mat_B[25][20] +
                  mat_A[17][26] * mat_B[26][20] +
                  mat_A[17][27] * mat_B[27][20] +
                  mat_A[17][28] * mat_B[28][20] +
                  mat_A[17][29] * mat_B[29][20] +
                  mat_A[17][30] * mat_B[30][20] +
                  mat_A[17][31] * mat_B[31][20];
    mat_C[17][21] <= 
                  mat_A[17][0] * mat_B[0][21] +
                  mat_A[17][1] * mat_B[1][21] +
                  mat_A[17][2] * mat_B[2][21] +
                  mat_A[17][3] * mat_B[3][21] +
                  mat_A[17][4] * mat_B[4][21] +
                  mat_A[17][5] * mat_B[5][21] +
                  mat_A[17][6] * mat_B[6][21] +
                  mat_A[17][7] * mat_B[7][21] +
                  mat_A[17][8] * mat_B[8][21] +
                  mat_A[17][9] * mat_B[9][21] +
                  mat_A[17][10] * mat_B[10][21] +
                  mat_A[17][11] * mat_B[11][21] +
                  mat_A[17][12] * mat_B[12][21] +
                  mat_A[17][13] * mat_B[13][21] +
                  mat_A[17][14] * mat_B[14][21] +
                  mat_A[17][15] * mat_B[15][21] +
                  mat_A[17][16] * mat_B[16][21] +
                  mat_A[17][17] * mat_B[17][21] +
                  mat_A[17][18] * mat_B[18][21] +
                  mat_A[17][19] * mat_B[19][21] +
                  mat_A[17][20] * mat_B[20][21] +
                  mat_A[17][21] * mat_B[21][21] +
                  mat_A[17][22] * mat_B[22][21] +
                  mat_A[17][23] * mat_B[23][21] +
                  mat_A[17][24] * mat_B[24][21] +
                  mat_A[17][25] * mat_B[25][21] +
                  mat_A[17][26] * mat_B[26][21] +
                  mat_A[17][27] * mat_B[27][21] +
                  mat_A[17][28] * mat_B[28][21] +
                  mat_A[17][29] * mat_B[29][21] +
                  mat_A[17][30] * mat_B[30][21] +
                  mat_A[17][31] * mat_B[31][21];
    mat_C[17][22] <= 
                  mat_A[17][0] * mat_B[0][22] +
                  mat_A[17][1] * mat_B[1][22] +
                  mat_A[17][2] * mat_B[2][22] +
                  mat_A[17][3] * mat_B[3][22] +
                  mat_A[17][4] * mat_B[4][22] +
                  mat_A[17][5] * mat_B[5][22] +
                  mat_A[17][6] * mat_B[6][22] +
                  mat_A[17][7] * mat_B[7][22] +
                  mat_A[17][8] * mat_B[8][22] +
                  mat_A[17][9] * mat_B[9][22] +
                  mat_A[17][10] * mat_B[10][22] +
                  mat_A[17][11] * mat_B[11][22] +
                  mat_A[17][12] * mat_B[12][22] +
                  mat_A[17][13] * mat_B[13][22] +
                  mat_A[17][14] * mat_B[14][22] +
                  mat_A[17][15] * mat_B[15][22] +
                  mat_A[17][16] * mat_B[16][22] +
                  mat_A[17][17] * mat_B[17][22] +
                  mat_A[17][18] * mat_B[18][22] +
                  mat_A[17][19] * mat_B[19][22] +
                  mat_A[17][20] * mat_B[20][22] +
                  mat_A[17][21] * mat_B[21][22] +
                  mat_A[17][22] * mat_B[22][22] +
                  mat_A[17][23] * mat_B[23][22] +
                  mat_A[17][24] * mat_B[24][22] +
                  mat_A[17][25] * mat_B[25][22] +
                  mat_A[17][26] * mat_B[26][22] +
                  mat_A[17][27] * mat_B[27][22] +
                  mat_A[17][28] * mat_B[28][22] +
                  mat_A[17][29] * mat_B[29][22] +
                  mat_A[17][30] * mat_B[30][22] +
                  mat_A[17][31] * mat_B[31][22];
    mat_C[17][23] <= 
                  mat_A[17][0] * mat_B[0][23] +
                  mat_A[17][1] * mat_B[1][23] +
                  mat_A[17][2] * mat_B[2][23] +
                  mat_A[17][3] * mat_B[3][23] +
                  mat_A[17][4] * mat_B[4][23] +
                  mat_A[17][5] * mat_B[5][23] +
                  mat_A[17][6] * mat_B[6][23] +
                  mat_A[17][7] * mat_B[7][23] +
                  mat_A[17][8] * mat_B[8][23] +
                  mat_A[17][9] * mat_B[9][23] +
                  mat_A[17][10] * mat_B[10][23] +
                  mat_A[17][11] * mat_B[11][23] +
                  mat_A[17][12] * mat_B[12][23] +
                  mat_A[17][13] * mat_B[13][23] +
                  mat_A[17][14] * mat_B[14][23] +
                  mat_A[17][15] * mat_B[15][23] +
                  mat_A[17][16] * mat_B[16][23] +
                  mat_A[17][17] * mat_B[17][23] +
                  mat_A[17][18] * mat_B[18][23] +
                  mat_A[17][19] * mat_B[19][23] +
                  mat_A[17][20] * mat_B[20][23] +
                  mat_A[17][21] * mat_B[21][23] +
                  mat_A[17][22] * mat_B[22][23] +
                  mat_A[17][23] * mat_B[23][23] +
                  mat_A[17][24] * mat_B[24][23] +
                  mat_A[17][25] * mat_B[25][23] +
                  mat_A[17][26] * mat_B[26][23] +
                  mat_A[17][27] * mat_B[27][23] +
                  mat_A[17][28] * mat_B[28][23] +
                  mat_A[17][29] * mat_B[29][23] +
                  mat_A[17][30] * mat_B[30][23] +
                  mat_A[17][31] * mat_B[31][23];
    mat_C[17][24] <= 
                  mat_A[17][0] * mat_B[0][24] +
                  mat_A[17][1] * mat_B[1][24] +
                  mat_A[17][2] * mat_B[2][24] +
                  mat_A[17][3] * mat_B[3][24] +
                  mat_A[17][4] * mat_B[4][24] +
                  mat_A[17][5] * mat_B[5][24] +
                  mat_A[17][6] * mat_B[6][24] +
                  mat_A[17][7] * mat_B[7][24] +
                  mat_A[17][8] * mat_B[8][24] +
                  mat_A[17][9] * mat_B[9][24] +
                  mat_A[17][10] * mat_B[10][24] +
                  mat_A[17][11] * mat_B[11][24] +
                  mat_A[17][12] * mat_B[12][24] +
                  mat_A[17][13] * mat_B[13][24] +
                  mat_A[17][14] * mat_B[14][24] +
                  mat_A[17][15] * mat_B[15][24] +
                  mat_A[17][16] * mat_B[16][24] +
                  mat_A[17][17] * mat_B[17][24] +
                  mat_A[17][18] * mat_B[18][24] +
                  mat_A[17][19] * mat_B[19][24] +
                  mat_A[17][20] * mat_B[20][24] +
                  mat_A[17][21] * mat_B[21][24] +
                  mat_A[17][22] * mat_B[22][24] +
                  mat_A[17][23] * mat_B[23][24] +
                  mat_A[17][24] * mat_B[24][24] +
                  mat_A[17][25] * mat_B[25][24] +
                  mat_A[17][26] * mat_B[26][24] +
                  mat_A[17][27] * mat_B[27][24] +
                  mat_A[17][28] * mat_B[28][24] +
                  mat_A[17][29] * mat_B[29][24] +
                  mat_A[17][30] * mat_B[30][24] +
                  mat_A[17][31] * mat_B[31][24];
    mat_C[17][25] <= 
                  mat_A[17][0] * mat_B[0][25] +
                  mat_A[17][1] * mat_B[1][25] +
                  mat_A[17][2] * mat_B[2][25] +
                  mat_A[17][3] * mat_B[3][25] +
                  mat_A[17][4] * mat_B[4][25] +
                  mat_A[17][5] * mat_B[5][25] +
                  mat_A[17][6] * mat_B[6][25] +
                  mat_A[17][7] * mat_B[7][25] +
                  mat_A[17][8] * mat_B[8][25] +
                  mat_A[17][9] * mat_B[9][25] +
                  mat_A[17][10] * mat_B[10][25] +
                  mat_A[17][11] * mat_B[11][25] +
                  mat_A[17][12] * mat_B[12][25] +
                  mat_A[17][13] * mat_B[13][25] +
                  mat_A[17][14] * mat_B[14][25] +
                  mat_A[17][15] * mat_B[15][25] +
                  mat_A[17][16] * mat_B[16][25] +
                  mat_A[17][17] * mat_B[17][25] +
                  mat_A[17][18] * mat_B[18][25] +
                  mat_A[17][19] * mat_B[19][25] +
                  mat_A[17][20] * mat_B[20][25] +
                  mat_A[17][21] * mat_B[21][25] +
                  mat_A[17][22] * mat_B[22][25] +
                  mat_A[17][23] * mat_B[23][25] +
                  mat_A[17][24] * mat_B[24][25] +
                  mat_A[17][25] * mat_B[25][25] +
                  mat_A[17][26] * mat_B[26][25] +
                  mat_A[17][27] * mat_B[27][25] +
                  mat_A[17][28] * mat_B[28][25] +
                  mat_A[17][29] * mat_B[29][25] +
                  mat_A[17][30] * mat_B[30][25] +
                  mat_A[17][31] * mat_B[31][25];
    mat_C[17][26] <= 
                  mat_A[17][0] * mat_B[0][26] +
                  mat_A[17][1] * mat_B[1][26] +
                  mat_A[17][2] * mat_B[2][26] +
                  mat_A[17][3] * mat_B[3][26] +
                  mat_A[17][4] * mat_B[4][26] +
                  mat_A[17][5] * mat_B[5][26] +
                  mat_A[17][6] * mat_B[6][26] +
                  mat_A[17][7] * mat_B[7][26] +
                  mat_A[17][8] * mat_B[8][26] +
                  mat_A[17][9] * mat_B[9][26] +
                  mat_A[17][10] * mat_B[10][26] +
                  mat_A[17][11] * mat_B[11][26] +
                  mat_A[17][12] * mat_B[12][26] +
                  mat_A[17][13] * mat_B[13][26] +
                  mat_A[17][14] * mat_B[14][26] +
                  mat_A[17][15] * mat_B[15][26] +
                  mat_A[17][16] * mat_B[16][26] +
                  mat_A[17][17] * mat_B[17][26] +
                  mat_A[17][18] * mat_B[18][26] +
                  mat_A[17][19] * mat_B[19][26] +
                  mat_A[17][20] * mat_B[20][26] +
                  mat_A[17][21] * mat_B[21][26] +
                  mat_A[17][22] * mat_B[22][26] +
                  mat_A[17][23] * mat_B[23][26] +
                  mat_A[17][24] * mat_B[24][26] +
                  mat_A[17][25] * mat_B[25][26] +
                  mat_A[17][26] * mat_B[26][26] +
                  mat_A[17][27] * mat_B[27][26] +
                  mat_A[17][28] * mat_B[28][26] +
                  mat_A[17][29] * mat_B[29][26] +
                  mat_A[17][30] * mat_B[30][26] +
                  mat_A[17][31] * mat_B[31][26];
    mat_C[17][27] <= 
                  mat_A[17][0] * mat_B[0][27] +
                  mat_A[17][1] * mat_B[1][27] +
                  mat_A[17][2] * mat_B[2][27] +
                  mat_A[17][3] * mat_B[3][27] +
                  mat_A[17][4] * mat_B[4][27] +
                  mat_A[17][5] * mat_B[5][27] +
                  mat_A[17][6] * mat_B[6][27] +
                  mat_A[17][7] * mat_B[7][27] +
                  mat_A[17][8] * mat_B[8][27] +
                  mat_A[17][9] * mat_B[9][27] +
                  mat_A[17][10] * mat_B[10][27] +
                  mat_A[17][11] * mat_B[11][27] +
                  mat_A[17][12] * mat_B[12][27] +
                  mat_A[17][13] * mat_B[13][27] +
                  mat_A[17][14] * mat_B[14][27] +
                  mat_A[17][15] * mat_B[15][27] +
                  mat_A[17][16] * mat_B[16][27] +
                  mat_A[17][17] * mat_B[17][27] +
                  mat_A[17][18] * mat_B[18][27] +
                  mat_A[17][19] * mat_B[19][27] +
                  mat_A[17][20] * mat_B[20][27] +
                  mat_A[17][21] * mat_B[21][27] +
                  mat_A[17][22] * mat_B[22][27] +
                  mat_A[17][23] * mat_B[23][27] +
                  mat_A[17][24] * mat_B[24][27] +
                  mat_A[17][25] * mat_B[25][27] +
                  mat_A[17][26] * mat_B[26][27] +
                  mat_A[17][27] * mat_B[27][27] +
                  mat_A[17][28] * mat_B[28][27] +
                  mat_A[17][29] * mat_B[29][27] +
                  mat_A[17][30] * mat_B[30][27] +
                  mat_A[17][31] * mat_B[31][27];
    mat_C[17][28] <= 
                  mat_A[17][0] * mat_B[0][28] +
                  mat_A[17][1] * mat_B[1][28] +
                  mat_A[17][2] * mat_B[2][28] +
                  mat_A[17][3] * mat_B[3][28] +
                  mat_A[17][4] * mat_B[4][28] +
                  mat_A[17][5] * mat_B[5][28] +
                  mat_A[17][6] * mat_B[6][28] +
                  mat_A[17][7] * mat_B[7][28] +
                  mat_A[17][8] * mat_B[8][28] +
                  mat_A[17][9] * mat_B[9][28] +
                  mat_A[17][10] * mat_B[10][28] +
                  mat_A[17][11] * mat_B[11][28] +
                  mat_A[17][12] * mat_B[12][28] +
                  mat_A[17][13] * mat_B[13][28] +
                  mat_A[17][14] * mat_B[14][28] +
                  mat_A[17][15] * mat_B[15][28] +
                  mat_A[17][16] * mat_B[16][28] +
                  mat_A[17][17] * mat_B[17][28] +
                  mat_A[17][18] * mat_B[18][28] +
                  mat_A[17][19] * mat_B[19][28] +
                  mat_A[17][20] * mat_B[20][28] +
                  mat_A[17][21] * mat_B[21][28] +
                  mat_A[17][22] * mat_B[22][28] +
                  mat_A[17][23] * mat_B[23][28] +
                  mat_A[17][24] * mat_B[24][28] +
                  mat_A[17][25] * mat_B[25][28] +
                  mat_A[17][26] * mat_B[26][28] +
                  mat_A[17][27] * mat_B[27][28] +
                  mat_A[17][28] * mat_B[28][28] +
                  mat_A[17][29] * mat_B[29][28] +
                  mat_A[17][30] * mat_B[30][28] +
                  mat_A[17][31] * mat_B[31][28];
    mat_C[17][29] <= 
                  mat_A[17][0] * mat_B[0][29] +
                  mat_A[17][1] * mat_B[1][29] +
                  mat_A[17][2] * mat_B[2][29] +
                  mat_A[17][3] * mat_B[3][29] +
                  mat_A[17][4] * mat_B[4][29] +
                  mat_A[17][5] * mat_B[5][29] +
                  mat_A[17][6] * mat_B[6][29] +
                  mat_A[17][7] * mat_B[7][29] +
                  mat_A[17][8] * mat_B[8][29] +
                  mat_A[17][9] * mat_B[9][29] +
                  mat_A[17][10] * mat_B[10][29] +
                  mat_A[17][11] * mat_B[11][29] +
                  mat_A[17][12] * mat_B[12][29] +
                  mat_A[17][13] * mat_B[13][29] +
                  mat_A[17][14] * mat_B[14][29] +
                  mat_A[17][15] * mat_B[15][29] +
                  mat_A[17][16] * mat_B[16][29] +
                  mat_A[17][17] * mat_B[17][29] +
                  mat_A[17][18] * mat_B[18][29] +
                  mat_A[17][19] * mat_B[19][29] +
                  mat_A[17][20] * mat_B[20][29] +
                  mat_A[17][21] * mat_B[21][29] +
                  mat_A[17][22] * mat_B[22][29] +
                  mat_A[17][23] * mat_B[23][29] +
                  mat_A[17][24] * mat_B[24][29] +
                  mat_A[17][25] * mat_B[25][29] +
                  mat_A[17][26] * mat_B[26][29] +
                  mat_A[17][27] * mat_B[27][29] +
                  mat_A[17][28] * mat_B[28][29] +
                  mat_A[17][29] * mat_B[29][29] +
                  mat_A[17][30] * mat_B[30][29] +
                  mat_A[17][31] * mat_B[31][29];
    mat_C[17][30] <= 
                  mat_A[17][0] * mat_B[0][30] +
                  mat_A[17][1] * mat_B[1][30] +
                  mat_A[17][2] * mat_B[2][30] +
                  mat_A[17][3] * mat_B[3][30] +
                  mat_A[17][4] * mat_B[4][30] +
                  mat_A[17][5] * mat_B[5][30] +
                  mat_A[17][6] * mat_B[6][30] +
                  mat_A[17][7] * mat_B[7][30] +
                  mat_A[17][8] * mat_B[8][30] +
                  mat_A[17][9] * mat_B[9][30] +
                  mat_A[17][10] * mat_B[10][30] +
                  mat_A[17][11] * mat_B[11][30] +
                  mat_A[17][12] * mat_B[12][30] +
                  mat_A[17][13] * mat_B[13][30] +
                  mat_A[17][14] * mat_B[14][30] +
                  mat_A[17][15] * mat_B[15][30] +
                  mat_A[17][16] * mat_B[16][30] +
                  mat_A[17][17] * mat_B[17][30] +
                  mat_A[17][18] * mat_B[18][30] +
                  mat_A[17][19] * mat_B[19][30] +
                  mat_A[17][20] * mat_B[20][30] +
                  mat_A[17][21] * mat_B[21][30] +
                  mat_A[17][22] * mat_B[22][30] +
                  mat_A[17][23] * mat_B[23][30] +
                  mat_A[17][24] * mat_B[24][30] +
                  mat_A[17][25] * mat_B[25][30] +
                  mat_A[17][26] * mat_B[26][30] +
                  mat_A[17][27] * mat_B[27][30] +
                  mat_A[17][28] * mat_B[28][30] +
                  mat_A[17][29] * mat_B[29][30] +
                  mat_A[17][30] * mat_B[30][30] +
                  mat_A[17][31] * mat_B[31][30];
    mat_C[17][31] <= 
                  mat_A[17][0] * mat_B[0][31] +
                  mat_A[17][1] * mat_B[1][31] +
                  mat_A[17][2] * mat_B[2][31] +
                  mat_A[17][3] * mat_B[3][31] +
                  mat_A[17][4] * mat_B[4][31] +
                  mat_A[17][5] * mat_B[5][31] +
                  mat_A[17][6] * mat_B[6][31] +
                  mat_A[17][7] * mat_B[7][31] +
                  mat_A[17][8] * mat_B[8][31] +
                  mat_A[17][9] * mat_B[9][31] +
                  mat_A[17][10] * mat_B[10][31] +
                  mat_A[17][11] * mat_B[11][31] +
                  mat_A[17][12] * mat_B[12][31] +
                  mat_A[17][13] * mat_B[13][31] +
                  mat_A[17][14] * mat_B[14][31] +
                  mat_A[17][15] * mat_B[15][31] +
                  mat_A[17][16] * mat_B[16][31] +
                  mat_A[17][17] * mat_B[17][31] +
                  mat_A[17][18] * mat_B[18][31] +
                  mat_A[17][19] * mat_B[19][31] +
                  mat_A[17][20] * mat_B[20][31] +
                  mat_A[17][21] * mat_B[21][31] +
                  mat_A[17][22] * mat_B[22][31] +
                  mat_A[17][23] * mat_B[23][31] +
                  mat_A[17][24] * mat_B[24][31] +
                  mat_A[17][25] * mat_B[25][31] +
                  mat_A[17][26] * mat_B[26][31] +
                  mat_A[17][27] * mat_B[27][31] +
                  mat_A[17][28] * mat_B[28][31] +
                  mat_A[17][29] * mat_B[29][31] +
                  mat_A[17][30] * mat_B[30][31] +
                  mat_A[17][31] * mat_B[31][31];
    mat_C[18][0] <= 
                  mat_A[18][0] * mat_B[0][0] +
                  mat_A[18][1] * mat_B[1][0] +
                  mat_A[18][2] * mat_B[2][0] +
                  mat_A[18][3] * mat_B[3][0] +
                  mat_A[18][4] * mat_B[4][0] +
                  mat_A[18][5] * mat_B[5][0] +
                  mat_A[18][6] * mat_B[6][0] +
                  mat_A[18][7] * mat_B[7][0] +
                  mat_A[18][8] * mat_B[8][0] +
                  mat_A[18][9] * mat_B[9][0] +
                  mat_A[18][10] * mat_B[10][0] +
                  mat_A[18][11] * mat_B[11][0] +
                  mat_A[18][12] * mat_B[12][0] +
                  mat_A[18][13] * mat_B[13][0] +
                  mat_A[18][14] * mat_B[14][0] +
                  mat_A[18][15] * mat_B[15][0] +
                  mat_A[18][16] * mat_B[16][0] +
                  mat_A[18][17] * mat_B[17][0] +
                  mat_A[18][18] * mat_B[18][0] +
                  mat_A[18][19] * mat_B[19][0] +
                  mat_A[18][20] * mat_B[20][0] +
                  mat_A[18][21] * mat_B[21][0] +
                  mat_A[18][22] * mat_B[22][0] +
                  mat_A[18][23] * mat_B[23][0] +
                  mat_A[18][24] * mat_B[24][0] +
                  mat_A[18][25] * mat_B[25][0] +
                  mat_A[18][26] * mat_B[26][0] +
                  mat_A[18][27] * mat_B[27][0] +
                  mat_A[18][28] * mat_B[28][0] +
                  mat_A[18][29] * mat_B[29][0] +
                  mat_A[18][30] * mat_B[30][0] +
                  mat_A[18][31] * mat_B[31][0];
    mat_C[18][1] <= 
                  mat_A[18][0] * mat_B[0][1] +
                  mat_A[18][1] * mat_B[1][1] +
                  mat_A[18][2] * mat_B[2][1] +
                  mat_A[18][3] * mat_B[3][1] +
                  mat_A[18][4] * mat_B[4][1] +
                  mat_A[18][5] * mat_B[5][1] +
                  mat_A[18][6] * mat_B[6][1] +
                  mat_A[18][7] * mat_B[7][1] +
                  mat_A[18][8] * mat_B[8][1] +
                  mat_A[18][9] * mat_B[9][1] +
                  mat_A[18][10] * mat_B[10][1] +
                  mat_A[18][11] * mat_B[11][1] +
                  mat_A[18][12] * mat_B[12][1] +
                  mat_A[18][13] * mat_B[13][1] +
                  mat_A[18][14] * mat_B[14][1] +
                  mat_A[18][15] * mat_B[15][1] +
                  mat_A[18][16] * mat_B[16][1] +
                  mat_A[18][17] * mat_B[17][1] +
                  mat_A[18][18] * mat_B[18][1] +
                  mat_A[18][19] * mat_B[19][1] +
                  mat_A[18][20] * mat_B[20][1] +
                  mat_A[18][21] * mat_B[21][1] +
                  mat_A[18][22] * mat_B[22][1] +
                  mat_A[18][23] * mat_B[23][1] +
                  mat_A[18][24] * mat_B[24][1] +
                  mat_A[18][25] * mat_B[25][1] +
                  mat_A[18][26] * mat_B[26][1] +
                  mat_A[18][27] * mat_B[27][1] +
                  mat_A[18][28] * mat_B[28][1] +
                  mat_A[18][29] * mat_B[29][1] +
                  mat_A[18][30] * mat_B[30][1] +
                  mat_A[18][31] * mat_B[31][1];
    mat_C[18][2] <= 
                  mat_A[18][0] * mat_B[0][2] +
                  mat_A[18][1] * mat_B[1][2] +
                  mat_A[18][2] * mat_B[2][2] +
                  mat_A[18][3] * mat_B[3][2] +
                  mat_A[18][4] * mat_B[4][2] +
                  mat_A[18][5] * mat_B[5][2] +
                  mat_A[18][6] * mat_B[6][2] +
                  mat_A[18][7] * mat_B[7][2] +
                  mat_A[18][8] * mat_B[8][2] +
                  mat_A[18][9] * mat_B[9][2] +
                  mat_A[18][10] * mat_B[10][2] +
                  mat_A[18][11] * mat_B[11][2] +
                  mat_A[18][12] * mat_B[12][2] +
                  mat_A[18][13] * mat_B[13][2] +
                  mat_A[18][14] * mat_B[14][2] +
                  mat_A[18][15] * mat_B[15][2] +
                  mat_A[18][16] * mat_B[16][2] +
                  mat_A[18][17] * mat_B[17][2] +
                  mat_A[18][18] * mat_B[18][2] +
                  mat_A[18][19] * mat_B[19][2] +
                  mat_A[18][20] * mat_B[20][2] +
                  mat_A[18][21] * mat_B[21][2] +
                  mat_A[18][22] * mat_B[22][2] +
                  mat_A[18][23] * mat_B[23][2] +
                  mat_A[18][24] * mat_B[24][2] +
                  mat_A[18][25] * mat_B[25][2] +
                  mat_A[18][26] * mat_B[26][2] +
                  mat_A[18][27] * mat_B[27][2] +
                  mat_A[18][28] * mat_B[28][2] +
                  mat_A[18][29] * mat_B[29][2] +
                  mat_A[18][30] * mat_B[30][2] +
                  mat_A[18][31] * mat_B[31][2];
    mat_C[18][3] <= 
                  mat_A[18][0] * mat_B[0][3] +
                  mat_A[18][1] * mat_B[1][3] +
                  mat_A[18][2] * mat_B[2][3] +
                  mat_A[18][3] * mat_B[3][3] +
                  mat_A[18][4] * mat_B[4][3] +
                  mat_A[18][5] * mat_B[5][3] +
                  mat_A[18][6] * mat_B[6][3] +
                  mat_A[18][7] * mat_B[7][3] +
                  mat_A[18][8] * mat_B[8][3] +
                  mat_A[18][9] * mat_B[9][3] +
                  mat_A[18][10] * mat_B[10][3] +
                  mat_A[18][11] * mat_B[11][3] +
                  mat_A[18][12] * mat_B[12][3] +
                  mat_A[18][13] * mat_B[13][3] +
                  mat_A[18][14] * mat_B[14][3] +
                  mat_A[18][15] * mat_B[15][3] +
                  mat_A[18][16] * mat_B[16][3] +
                  mat_A[18][17] * mat_B[17][3] +
                  mat_A[18][18] * mat_B[18][3] +
                  mat_A[18][19] * mat_B[19][3] +
                  mat_A[18][20] * mat_B[20][3] +
                  mat_A[18][21] * mat_B[21][3] +
                  mat_A[18][22] * mat_B[22][3] +
                  mat_A[18][23] * mat_B[23][3] +
                  mat_A[18][24] * mat_B[24][3] +
                  mat_A[18][25] * mat_B[25][3] +
                  mat_A[18][26] * mat_B[26][3] +
                  mat_A[18][27] * mat_B[27][3] +
                  mat_A[18][28] * mat_B[28][3] +
                  mat_A[18][29] * mat_B[29][3] +
                  mat_A[18][30] * mat_B[30][3] +
                  mat_A[18][31] * mat_B[31][3];
    mat_C[18][4] <= 
                  mat_A[18][0] * mat_B[0][4] +
                  mat_A[18][1] * mat_B[1][4] +
                  mat_A[18][2] * mat_B[2][4] +
                  mat_A[18][3] * mat_B[3][4] +
                  mat_A[18][4] * mat_B[4][4] +
                  mat_A[18][5] * mat_B[5][4] +
                  mat_A[18][6] * mat_B[6][4] +
                  mat_A[18][7] * mat_B[7][4] +
                  mat_A[18][8] * mat_B[8][4] +
                  mat_A[18][9] * mat_B[9][4] +
                  mat_A[18][10] * mat_B[10][4] +
                  mat_A[18][11] * mat_B[11][4] +
                  mat_A[18][12] * mat_B[12][4] +
                  mat_A[18][13] * mat_B[13][4] +
                  mat_A[18][14] * mat_B[14][4] +
                  mat_A[18][15] * mat_B[15][4] +
                  mat_A[18][16] * mat_B[16][4] +
                  mat_A[18][17] * mat_B[17][4] +
                  mat_A[18][18] * mat_B[18][4] +
                  mat_A[18][19] * mat_B[19][4] +
                  mat_A[18][20] * mat_B[20][4] +
                  mat_A[18][21] * mat_B[21][4] +
                  mat_A[18][22] * mat_B[22][4] +
                  mat_A[18][23] * mat_B[23][4] +
                  mat_A[18][24] * mat_B[24][4] +
                  mat_A[18][25] * mat_B[25][4] +
                  mat_A[18][26] * mat_B[26][4] +
                  mat_A[18][27] * mat_B[27][4] +
                  mat_A[18][28] * mat_B[28][4] +
                  mat_A[18][29] * mat_B[29][4] +
                  mat_A[18][30] * mat_B[30][4] +
                  mat_A[18][31] * mat_B[31][4];
    mat_C[18][5] <= 
                  mat_A[18][0] * mat_B[0][5] +
                  mat_A[18][1] * mat_B[1][5] +
                  mat_A[18][2] * mat_B[2][5] +
                  mat_A[18][3] * mat_B[3][5] +
                  mat_A[18][4] * mat_B[4][5] +
                  mat_A[18][5] * mat_B[5][5] +
                  mat_A[18][6] * mat_B[6][5] +
                  mat_A[18][7] * mat_B[7][5] +
                  mat_A[18][8] * mat_B[8][5] +
                  mat_A[18][9] * mat_B[9][5] +
                  mat_A[18][10] * mat_B[10][5] +
                  mat_A[18][11] * mat_B[11][5] +
                  mat_A[18][12] * mat_B[12][5] +
                  mat_A[18][13] * mat_B[13][5] +
                  mat_A[18][14] * mat_B[14][5] +
                  mat_A[18][15] * mat_B[15][5] +
                  mat_A[18][16] * mat_B[16][5] +
                  mat_A[18][17] * mat_B[17][5] +
                  mat_A[18][18] * mat_B[18][5] +
                  mat_A[18][19] * mat_B[19][5] +
                  mat_A[18][20] * mat_B[20][5] +
                  mat_A[18][21] * mat_B[21][5] +
                  mat_A[18][22] * mat_B[22][5] +
                  mat_A[18][23] * mat_B[23][5] +
                  mat_A[18][24] * mat_B[24][5] +
                  mat_A[18][25] * mat_B[25][5] +
                  mat_A[18][26] * mat_B[26][5] +
                  mat_A[18][27] * mat_B[27][5] +
                  mat_A[18][28] * mat_B[28][5] +
                  mat_A[18][29] * mat_B[29][5] +
                  mat_A[18][30] * mat_B[30][5] +
                  mat_A[18][31] * mat_B[31][5];
    mat_C[18][6] <= 
                  mat_A[18][0] * mat_B[0][6] +
                  mat_A[18][1] * mat_B[1][6] +
                  mat_A[18][2] * mat_B[2][6] +
                  mat_A[18][3] * mat_B[3][6] +
                  mat_A[18][4] * mat_B[4][6] +
                  mat_A[18][5] * mat_B[5][6] +
                  mat_A[18][6] * mat_B[6][6] +
                  mat_A[18][7] * mat_B[7][6] +
                  mat_A[18][8] * mat_B[8][6] +
                  mat_A[18][9] * mat_B[9][6] +
                  mat_A[18][10] * mat_B[10][6] +
                  mat_A[18][11] * mat_B[11][6] +
                  mat_A[18][12] * mat_B[12][6] +
                  mat_A[18][13] * mat_B[13][6] +
                  mat_A[18][14] * mat_B[14][6] +
                  mat_A[18][15] * mat_B[15][6] +
                  mat_A[18][16] * mat_B[16][6] +
                  mat_A[18][17] * mat_B[17][6] +
                  mat_A[18][18] * mat_B[18][6] +
                  mat_A[18][19] * mat_B[19][6] +
                  mat_A[18][20] * mat_B[20][6] +
                  mat_A[18][21] * mat_B[21][6] +
                  mat_A[18][22] * mat_B[22][6] +
                  mat_A[18][23] * mat_B[23][6] +
                  mat_A[18][24] * mat_B[24][6] +
                  mat_A[18][25] * mat_B[25][6] +
                  mat_A[18][26] * mat_B[26][6] +
                  mat_A[18][27] * mat_B[27][6] +
                  mat_A[18][28] * mat_B[28][6] +
                  mat_A[18][29] * mat_B[29][6] +
                  mat_A[18][30] * mat_B[30][6] +
                  mat_A[18][31] * mat_B[31][6];
    mat_C[18][7] <= 
                  mat_A[18][0] * mat_B[0][7] +
                  mat_A[18][1] * mat_B[1][7] +
                  mat_A[18][2] * mat_B[2][7] +
                  mat_A[18][3] * mat_B[3][7] +
                  mat_A[18][4] * mat_B[4][7] +
                  mat_A[18][5] * mat_B[5][7] +
                  mat_A[18][6] * mat_B[6][7] +
                  mat_A[18][7] * mat_B[7][7] +
                  mat_A[18][8] * mat_B[8][7] +
                  mat_A[18][9] * mat_B[9][7] +
                  mat_A[18][10] * mat_B[10][7] +
                  mat_A[18][11] * mat_B[11][7] +
                  mat_A[18][12] * mat_B[12][7] +
                  mat_A[18][13] * mat_B[13][7] +
                  mat_A[18][14] * mat_B[14][7] +
                  mat_A[18][15] * mat_B[15][7] +
                  mat_A[18][16] * mat_B[16][7] +
                  mat_A[18][17] * mat_B[17][7] +
                  mat_A[18][18] * mat_B[18][7] +
                  mat_A[18][19] * mat_B[19][7] +
                  mat_A[18][20] * mat_B[20][7] +
                  mat_A[18][21] * mat_B[21][7] +
                  mat_A[18][22] * mat_B[22][7] +
                  mat_A[18][23] * mat_B[23][7] +
                  mat_A[18][24] * mat_B[24][7] +
                  mat_A[18][25] * mat_B[25][7] +
                  mat_A[18][26] * mat_B[26][7] +
                  mat_A[18][27] * mat_B[27][7] +
                  mat_A[18][28] * mat_B[28][7] +
                  mat_A[18][29] * mat_B[29][7] +
                  mat_A[18][30] * mat_B[30][7] +
                  mat_A[18][31] * mat_B[31][7];
    mat_C[18][8] <= 
                  mat_A[18][0] * mat_B[0][8] +
                  mat_A[18][1] * mat_B[1][8] +
                  mat_A[18][2] * mat_B[2][8] +
                  mat_A[18][3] * mat_B[3][8] +
                  mat_A[18][4] * mat_B[4][8] +
                  mat_A[18][5] * mat_B[5][8] +
                  mat_A[18][6] * mat_B[6][8] +
                  mat_A[18][7] * mat_B[7][8] +
                  mat_A[18][8] * mat_B[8][8] +
                  mat_A[18][9] * mat_B[9][8] +
                  mat_A[18][10] * mat_B[10][8] +
                  mat_A[18][11] * mat_B[11][8] +
                  mat_A[18][12] * mat_B[12][8] +
                  mat_A[18][13] * mat_B[13][8] +
                  mat_A[18][14] * mat_B[14][8] +
                  mat_A[18][15] * mat_B[15][8] +
                  mat_A[18][16] * mat_B[16][8] +
                  mat_A[18][17] * mat_B[17][8] +
                  mat_A[18][18] * mat_B[18][8] +
                  mat_A[18][19] * mat_B[19][8] +
                  mat_A[18][20] * mat_B[20][8] +
                  mat_A[18][21] * mat_B[21][8] +
                  mat_A[18][22] * mat_B[22][8] +
                  mat_A[18][23] * mat_B[23][8] +
                  mat_A[18][24] * mat_B[24][8] +
                  mat_A[18][25] * mat_B[25][8] +
                  mat_A[18][26] * mat_B[26][8] +
                  mat_A[18][27] * mat_B[27][8] +
                  mat_A[18][28] * mat_B[28][8] +
                  mat_A[18][29] * mat_B[29][8] +
                  mat_A[18][30] * mat_B[30][8] +
                  mat_A[18][31] * mat_B[31][8];
    mat_C[18][9] <= 
                  mat_A[18][0] * mat_B[0][9] +
                  mat_A[18][1] * mat_B[1][9] +
                  mat_A[18][2] * mat_B[2][9] +
                  mat_A[18][3] * mat_B[3][9] +
                  mat_A[18][4] * mat_B[4][9] +
                  mat_A[18][5] * mat_B[5][9] +
                  mat_A[18][6] * mat_B[6][9] +
                  mat_A[18][7] * mat_B[7][9] +
                  mat_A[18][8] * mat_B[8][9] +
                  mat_A[18][9] * mat_B[9][9] +
                  mat_A[18][10] * mat_B[10][9] +
                  mat_A[18][11] * mat_B[11][9] +
                  mat_A[18][12] * mat_B[12][9] +
                  mat_A[18][13] * mat_B[13][9] +
                  mat_A[18][14] * mat_B[14][9] +
                  mat_A[18][15] * mat_B[15][9] +
                  mat_A[18][16] * mat_B[16][9] +
                  mat_A[18][17] * mat_B[17][9] +
                  mat_A[18][18] * mat_B[18][9] +
                  mat_A[18][19] * mat_B[19][9] +
                  mat_A[18][20] * mat_B[20][9] +
                  mat_A[18][21] * mat_B[21][9] +
                  mat_A[18][22] * mat_B[22][9] +
                  mat_A[18][23] * mat_B[23][9] +
                  mat_A[18][24] * mat_B[24][9] +
                  mat_A[18][25] * mat_B[25][9] +
                  mat_A[18][26] * mat_B[26][9] +
                  mat_A[18][27] * mat_B[27][9] +
                  mat_A[18][28] * mat_B[28][9] +
                  mat_A[18][29] * mat_B[29][9] +
                  mat_A[18][30] * mat_B[30][9] +
                  mat_A[18][31] * mat_B[31][9];
    mat_C[18][10] <= 
                  mat_A[18][0] * mat_B[0][10] +
                  mat_A[18][1] * mat_B[1][10] +
                  mat_A[18][2] * mat_B[2][10] +
                  mat_A[18][3] * mat_B[3][10] +
                  mat_A[18][4] * mat_B[4][10] +
                  mat_A[18][5] * mat_B[5][10] +
                  mat_A[18][6] * mat_B[6][10] +
                  mat_A[18][7] * mat_B[7][10] +
                  mat_A[18][8] * mat_B[8][10] +
                  mat_A[18][9] * mat_B[9][10] +
                  mat_A[18][10] * mat_B[10][10] +
                  mat_A[18][11] * mat_B[11][10] +
                  mat_A[18][12] * mat_B[12][10] +
                  mat_A[18][13] * mat_B[13][10] +
                  mat_A[18][14] * mat_B[14][10] +
                  mat_A[18][15] * mat_B[15][10] +
                  mat_A[18][16] * mat_B[16][10] +
                  mat_A[18][17] * mat_B[17][10] +
                  mat_A[18][18] * mat_B[18][10] +
                  mat_A[18][19] * mat_B[19][10] +
                  mat_A[18][20] * mat_B[20][10] +
                  mat_A[18][21] * mat_B[21][10] +
                  mat_A[18][22] * mat_B[22][10] +
                  mat_A[18][23] * mat_B[23][10] +
                  mat_A[18][24] * mat_B[24][10] +
                  mat_A[18][25] * mat_B[25][10] +
                  mat_A[18][26] * mat_B[26][10] +
                  mat_A[18][27] * mat_B[27][10] +
                  mat_A[18][28] * mat_B[28][10] +
                  mat_A[18][29] * mat_B[29][10] +
                  mat_A[18][30] * mat_B[30][10] +
                  mat_A[18][31] * mat_B[31][10];
    mat_C[18][11] <= 
                  mat_A[18][0] * mat_B[0][11] +
                  mat_A[18][1] * mat_B[1][11] +
                  mat_A[18][2] * mat_B[2][11] +
                  mat_A[18][3] * mat_B[3][11] +
                  mat_A[18][4] * mat_B[4][11] +
                  mat_A[18][5] * mat_B[5][11] +
                  mat_A[18][6] * mat_B[6][11] +
                  mat_A[18][7] * mat_B[7][11] +
                  mat_A[18][8] * mat_B[8][11] +
                  mat_A[18][9] * mat_B[9][11] +
                  mat_A[18][10] * mat_B[10][11] +
                  mat_A[18][11] * mat_B[11][11] +
                  mat_A[18][12] * mat_B[12][11] +
                  mat_A[18][13] * mat_B[13][11] +
                  mat_A[18][14] * mat_B[14][11] +
                  mat_A[18][15] * mat_B[15][11] +
                  mat_A[18][16] * mat_B[16][11] +
                  mat_A[18][17] * mat_B[17][11] +
                  mat_A[18][18] * mat_B[18][11] +
                  mat_A[18][19] * mat_B[19][11] +
                  mat_A[18][20] * mat_B[20][11] +
                  mat_A[18][21] * mat_B[21][11] +
                  mat_A[18][22] * mat_B[22][11] +
                  mat_A[18][23] * mat_B[23][11] +
                  mat_A[18][24] * mat_B[24][11] +
                  mat_A[18][25] * mat_B[25][11] +
                  mat_A[18][26] * mat_B[26][11] +
                  mat_A[18][27] * mat_B[27][11] +
                  mat_A[18][28] * mat_B[28][11] +
                  mat_A[18][29] * mat_B[29][11] +
                  mat_A[18][30] * mat_B[30][11] +
                  mat_A[18][31] * mat_B[31][11];
    mat_C[18][12] <= 
                  mat_A[18][0] * mat_B[0][12] +
                  mat_A[18][1] * mat_B[1][12] +
                  mat_A[18][2] * mat_B[2][12] +
                  mat_A[18][3] * mat_B[3][12] +
                  mat_A[18][4] * mat_B[4][12] +
                  mat_A[18][5] * mat_B[5][12] +
                  mat_A[18][6] * mat_B[6][12] +
                  mat_A[18][7] * mat_B[7][12] +
                  mat_A[18][8] * mat_B[8][12] +
                  mat_A[18][9] * mat_B[9][12] +
                  mat_A[18][10] * mat_B[10][12] +
                  mat_A[18][11] * mat_B[11][12] +
                  mat_A[18][12] * mat_B[12][12] +
                  mat_A[18][13] * mat_B[13][12] +
                  mat_A[18][14] * mat_B[14][12] +
                  mat_A[18][15] * mat_B[15][12] +
                  mat_A[18][16] * mat_B[16][12] +
                  mat_A[18][17] * mat_B[17][12] +
                  mat_A[18][18] * mat_B[18][12] +
                  mat_A[18][19] * mat_B[19][12] +
                  mat_A[18][20] * mat_B[20][12] +
                  mat_A[18][21] * mat_B[21][12] +
                  mat_A[18][22] * mat_B[22][12] +
                  mat_A[18][23] * mat_B[23][12] +
                  mat_A[18][24] * mat_B[24][12] +
                  mat_A[18][25] * mat_B[25][12] +
                  mat_A[18][26] * mat_B[26][12] +
                  mat_A[18][27] * mat_B[27][12] +
                  mat_A[18][28] * mat_B[28][12] +
                  mat_A[18][29] * mat_B[29][12] +
                  mat_A[18][30] * mat_B[30][12] +
                  mat_A[18][31] * mat_B[31][12];
    mat_C[18][13] <= 
                  mat_A[18][0] * mat_B[0][13] +
                  mat_A[18][1] * mat_B[1][13] +
                  mat_A[18][2] * mat_B[2][13] +
                  mat_A[18][3] * mat_B[3][13] +
                  mat_A[18][4] * mat_B[4][13] +
                  mat_A[18][5] * mat_B[5][13] +
                  mat_A[18][6] * mat_B[6][13] +
                  mat_A[18][7] * mat_B[7][13] +
                  mat_A[18][8] * mat_B[8][13] +
                  mat_A[18][9] * mat_B[9][13] +
                  mat_A[18][10] * mat_B[10][13] +
                  mat_A[18][11] * mat_B[11][13] +
                  mat_A[18][12] * mat_B[12][13] +
                  mat_A[18][13] * mat_B[13][13] +
                  mat_A[18][14] * mat_B[14][13] +
                  mat_A[18][15] * mat_B[15][13] +
                  mat_A[18][16] * mat_B[16][13] +
                  mat_A[18][17] * mat_B[17][13] +
                  mat_A[18][18] * mat_B[18][13] +
                  mat_A[18][19] * mat_B[19][13] +
                  mat_A[18][20] * mat_B[20][13] +
                  mat_A[18][21] * mat_B[21][13] +
                  mat_A[18][22] * mat_B[22][13] +
                  mat_A[18][23] * mat_B[23][13] +
                  mat_A[18][24] * mat_B[24][13] +
                  mat_A[18][25] * mat_B[25][13] +
                  mat_A[18][26] * mat_B[26][13] +
                  mat_A[18][27] * mat_B[27][13] +
                  mat_A[18][28] * mat_B[28][13] +
                  mat_A[18][29] * mat_B[29][13] +
                  mat_A[18][30] * mat_B[30][13] +
                  mat_A[18][31] * mat_B[31][13];
    mat_C[18][14] <= 
                  mat_A[18][0] * mat_B[0][14] +
                  mat_A[18][1] * mat_B[1][14] +
                  mat_A[18][2] * mat_B[2][14] +
                  mat_A[18][3] * mat_B[3][14] +
                  mat_A[18][4] * mat_B[4][14] +
                  mat_A[18][5] * mat_B[5][14] +
                  mat_A[18][6] * mat_B[6][14] +
                  mat_A[18][7] * mat_B[7][14] +
                  mat_A[18][8] * mat_B[8][14] +
                  mat_A[18][9] * mat_B[9][14] +
                  mat_A[18][10] * mat_B[10][14] +
                  mat_A[18][11] * mat_B[11][14] +
                  mat_A[18][12] * mat_B[12][14] +
                  mat_A[18][13] * mat_B[13][14] +
                  mat_A[18][14] * mat_B[14][14] +
                  mat_A[18][15] * mat_B[15][14] +
                  mat_A[18][16] * mat_B[16][14] +
                  mat_A[18][17] * mat_B[17][14] +
                  mat_A[18][18] * mat_B[18][14] +
                  mat_A[18][19] * mat_B[19][14] +
                  mat_A[18][20] * mat_B[20][14] +
                  mat_A[18][21] * mat_B[21][14] +
                  mat_A[18][22] * mat_B[22][14] +
                  mat_A[18][23] * mat_B[23][14] +
                  mat_A[18][24] * mat_B[24][14] +
                  mat_A[18][25] * mat_B[25][14] +
                  mat_A[18][26] * mat_B[26][14] +
                  mat_A[18][27] * mat_B[27][14] +
                  mat_A[18][28] * mat_B[28][14] +
                  mat_A[18][29] * mat_B[29][14] +
                  mat_A[18][30] * mat_B[30][14] +
                  mat_A[18][31] * mat_B[31][14];
    mat_C[18][15] <= 
                  mat_A[18][0] * mat_B[0][15] +
                  mat_A[18][1] * mat_B[1][15] +
                  mat_A[18][2] * mat_B[2][15] +
                  mat_A[18][3] * mat_B[3][15] +
                  mat_A[18][4] * mat_B[4][15] +
                  mat_A[18][5] * mat_B[5][15] +
                  mat_A[18][6] * mat_B[6][15] +
                  mat_A[18][7] * mat_B[7][15] +
                  mat_A[18][8] * mat_B[8][15] +
                  mat_A[18][9] * mat_B[9][15] +
                  mat_A[18][10] * mat_B[10][15] +
                  mat_A[18][11] * mat_B[11][15] +
                  mat_A[18][12] * mat_B[12][15] +
                  mat_A[18][13] * mat_B[13][15] +
                  mat_A[18][14] * mat_B[14][15] +
                  mat_A[18][15] * mat_B[15][15] +
                  mat_A[18][16] * mat_B[16][15] +
                  mat_A[18][17] * mat_B[17][15] +
                  mat_A[18][18] * mat_B[18][15] +
                  mat_A[18][19] * mat_B[19][15] +
                  mat_A[18][20] * mat_B[20][15] +
                  mat_A[18][21] * mat_B[21][15] +
                  mat_A[18][22] * mat_B[22][15] +
                  mat_A[18][23] * mat_B[23][15] +
                  mat_A[18][24] * mat_B[24][15] +
                  mat_A[18][25] * mat_B[25][15] +
                  mat_A[18][26] * mat_B[26][15] +
                  mat_A[18][27] * mat_B[27][15] +
                  mat_A[18][28] * mat_B[28][15] +
                  mat_A[18][29] * mat_B[29][15] +
                  mat_A[18][30] * mat_B[30][15] +
                  mat_A[18][31] * mat_B[31][15];
    mat_C[18][16] <= 
                  mat_A[18][0] * mat_B[0][16] +
                  mat_A[18][1] * mat_B[1][16] +
                  mat_A[18][2] * mat_B[2][16] +
                  mat_A[18][3] * mat_B[3][16] +
                  mat_A[18][4] * mat_B[4][16] +
                  mat_A[18][5] * mat_B[5][16] +
                  mat_A[18][6] * mat_B[6][16] +
                  mat_A[18][7] * mat_B[7][16] +
                  mat_A[18][8] * mat_B[8][16] +
                  mat_A[18][9] * mat_B[9][16] +
                  mat_A[18][10] * mat_B[10][16] +
                  mat_A[18][11] * mat_B[11][16] +
                  mat_A[18][12] * mat_B[12][16] +
                  mat_A[18][13] * mat_B[13][16] +
                  mat_A[18][14] * mat_B[14][16] +
                  mat_A[18][15] * mat_B[15][16] +
                  mat_A[18][16] * mat_B[16][16] +
                  mat_A[18][17] * mat_B[17][16] +
                  mat_A[18][18] * mat_B[18][16] +
                  mat_A[18][19] * mat_B[19][16] +
                  mat_A[18][20] * mat_B[20][16] +
                  mat_A[18][21] * mat_B[21][16] +
                  mat_A[18][22] * mat_B[22][16] +
                  mat_A[18][23] * mat_B[23][16] +
                  mat_A[18][24] * mat_B[24][16] +
                  mat_A[18][25] * mat_B[25][16] +
                  mat_A[18][26] * mat_B[26][16] +
                  mat_A[18][27] * mat_B[27][16] +
                  mat_A[18][28] * mat_B[28][16] +
                  mat_A[18][29] * mat_B[29][16] +
                  mat_A[18][30] * mat_B[30][16] +
                  mat_A[18][31] * mat_B[31][16];
    mat_C[18][17] <= 
                  mat_A[18][0] * mat_B[0][17] +
                  mat_A[18][1] * mat_B[1][17] +
                  mat_A[18][2] * mat_B[2][17] +
                  mat_A[18][3] * mat_B[3][17] +
                  mat_A[18][4] * mat_B[4][17] +
                  mat_A[18][5] * mat_B[5][17] +
                  mat_A[18][6] * mat_B[6][17] +
                  mat_A[18][7] * mat_B[7][17] +
                  mat_A[18][8] * mat_B[8][17] +
                  mat_A[18][9] * mat_B[9][17] +
                  mat_A[18][10] * mat_B[10][17] +
                  mat_A[18][11] * mat_B[11][17] +
                  mat_A[18][12] * mat_B[12][17] +
                  mat_A[18][13] * mat_B[13][17] +
                  mat_A[18][14] * mat_B[14][17] +
                  mat_A[18][15] * mat_B[15][17] +
                  mat_A[18][16] * mat_B[16][17] +
                  mat_A[18][17] * mat_B[17][17] +
                  mat_A[18][18] * mat_B[18][17] +
                  mat_A[18][19] * mat_B[19][17] +
                  mat_A[18][20] * mat_B[20][17] +
                  mat_A[18][21] * mat_B[21][17] +
                  mat_A[18][22] * mat_B[22][17] +
                  mat_A[18][23] * mat_B[23][17] +
                  mat_A[18][24] * mat_B[24][17] +
                  mat_A[18][25] * mat_B[25][17] +
                  mat_A[18][26] * mat_B[26][17] +
                  mat_A[18][27] * mat_B[27][17] +
                  mat_A[18][28] * mat_B[28][17] +
                  mat_A[18][29] * mat_B[29][17] +
                  mat_A[18][30] * mat_B[30][17] +
                  mat_A[18][31] * mat_B[31][17];
    mat_C[18][18] <= 
                  mat_A[18][0] * mat_B[0][18] +
                  mat_A[18][1] * mat_B[1][18] +
                  mat_A[18][2] * mat_B[2][18] +
                  mat_A[18][3] * mat_B[3][18] +
                  mat_A[18][4] * mat_B[4][18] +
                  mat_A[18][5] * mat_B[5][18] +
                  mat_A[18][6] * mat_B[6][18] +
                  mat_A[18][7] * mat_B[7][18] +
                  mat_A[18][8] * mat_B[8][18] +
                  mat_A[18][9] * mat_B[9][18] +
                  mat_A[18][10] * mat_B[10][18] +
                  mat_A[18][11] * mat_B[11][18] +
                  mat_A[18][12] * mat_B[12][18] +
                  mat_A[18][13] * mat_B[13][18] +
                  mat_A[18][14] * mat_B[14][18] +
                  mat_A[18][15] * mat_B[15][18] +
                  mat_A[18][16] * mat_B[16][18] +
                  mat_A[18][17] * mat_B[17][18] +
                  mat_A[18][18] * mat_B[18][18] +
                  mat_A[18][19] * mat_B[19][18] +
                  mat_A[18][20] * mat_B[20][18] +
                  mat_A[18][21] * mat_B[21][18] +
                  mat_A[18][22] * mat_B[22][18] +
                  mat_A[18][23] * mat_B[23][18] +
                  mat_A[18][24] * mat_B[24][18] +
                  mat_A[18][25] * mat_B[25][18] +
                  mat_A[18][26] * mat_B[26][18] +
                  mat_A[18][27] * mat_B[27][18] +
                  mat_A[18][28] * mat_B[28][18] +
                  mat_A[18][29] * mat_B[29][18] +
                  mat_A[18][30] * mat_B[30][18] +
                  mat_A[18][31] * mat_B[31][18];
    mat_C[18][19] <= 
                  mat_A[18][0] * mat_B[0][19] +
                  mat_A[18][1] * mat_B[1][19] +
                  mat_A[18][2] * mat_B[2][19] +
                  mat_A[18][3] * mat_B[3][19] +
                  mat_A[18][4] * mat_B[4][19] +
                  mat_A[18][5] * mat_B[5][19] +
                  mat_A[18][6] * mat_B[6][19] +
                  mat_A[18][7] * mat_B[7][19] +
                  mat_A[18][8] * mat_B[8][19] +
                  mat_A[18][9] * mat_B[9][19] +
                  mat_A[18][10] * mat_B[10][19] +
                  mat_A[18][11] * mat_B[11][19] +
                  mat_A[18][12] * mat_B[12][19] +
                  mat_A[18][13] * mat_B[13][19] +
                  mat_A[18][14] * mat_B[14][19] +
                  mat_A[18][15] * mat_B[15][19] +
                  mat_A[18][16] * mat_B[16][19] +
                  mat_A[18][17] * mat_B[17][19] +
                  mat_A[18][18] * mat_B[18][19] +
                  mat_A[18][19] * mat_B[19][19] +
                  mat_A[18][20] * mat_B[20][19] +
                  mat_A[18][21] * mat_B[21][19] +
                  mat_A[18][22] * mat_B[22][19] +
                  mat_A[18][23] * mat_B[23][19] +
                  mat_A[18][24] * mat_B[24][19] +
                  mat_A[18][25] * mat_B[25][19] +
                  mat_A[18][26] * mat_B[26][19] +
                  mat_A[18][27] * mat_B[27][19] +
                  mat_A[18][28] * mat_B[28][19] +
                  mat_A[18][29] * mat_B[29][19] +
                  mat_A[18][30] * mat_B[30][19] +
                  mat_A[18][31] * mat_B[31][19];
    mat_C[18][20] <= 
                  mat_A[18][0] * mat_B[0][20] +
                  mat_A[18][1] * mat_B[1][20] +
                  mat_A[18][2] * mat_B[2][20] +
                  mat_A[18][3] * mat_B[3][20] +
                  mat_A[18][4] * mat_B[4][20] +
                  mat_A[18][5] * mat_B[5][20] +
                  mat_A[18][6] * mat_B[6][20] +
                  mat_A[18][7] * mat_B[7][20] +
                  mat_A[18][8] * mat_B[8][20] +
                  mat_A[18][9] * mat_B[9][20] +
                  mat_A[18][10] * mat_B[10][20] +
                  mat_A[18][11] * mat_B[11][20] +
                  mat_A[18][12] * mat_B[12][20] +
                  mat_A[18][13] * mat_B[13][20] +
                  mat_A[18][14] * mat_B[14][20] +
                  mat_A[18][15] * mat_B[15][20] +
                  mat_A[18][16] * mat_B[16][20] +
                  mat_A[18][17] * mat_B[17][20] +
                  mat_A[18][18] * mat_B[18][20] +
                  mat_A[18][19] * mat_B[19][20] +
                  mat_A[18][20] * mat_B[20][20] +
                  mat_A[18][21] * mat_B[21][20] +
                  mat_A[18][22] * mat_B[22][20] +
                  mat_A[18][23] * mat_B[23][20] +
                  mat_A[18][24] * mat_B[24][20] +
                  mat_A[18][25] * mat_B[25][20] +
                  mat_A[18][26] * mat_B[26][20] +
                  mat_A[18][27] * mat_B[27][20] +
                  mat_A[18][28] * mat_B[28][20] +
                  mat_A[18][29] * mat_B[29][20] +
                  mat_A[18][30] * mat_B[30][20] +
                  mat_A[18][31] * mat_B[31][20];
    mat_C[18][21] <= 
                  mat_A[18][0] * mat_B[0][21] +
                  mat_A[18][1] * mat_B[1][21] +
                  mat_A[18][2] * mat_B[2][21] +
                  mat_A[18][3] * mat_B[3][21] +
                  mat_A[18][4] * mat_B[4][21] +
                  mat_A[18][5] * mat_B[5][21] +
                  mat_A[18][6] * mat_B[6][21] +
                  mat_A[18][7] * mat_B[7][21] +
                  mat_A[18][8] * mat_B[8][21] +
                  mat_A[18][9] * mat_B[9][21] +
                  mat_A[18][10] * mat_B[10][21] +
                  mat_A[18][11] * mat_B[11][21] +
                  mat_A[18][12] * mat_B[12][21] +
                  mat_A[18][13] * mat_B[13][21] +
                  mat_A[18][14] * mat_B[14][21] +
                  mat_A[18][15] * mat_B[15][21] +
                  mat_A[18][16] * mat_B[16][21] +
                  mat_A[18][17] * mat_B[17][21] +
                  mat_A[18][18] * mat_B[18][21] +
                  mat_A[18][19] * mat_B[19][21] +
                  mat_A[18][20] * mat_B[20][21] +
                  mat_A[18][21] * mat_B[21][21] +
                  mat_A[18][22] * mat_B[22][21] +
                  mat_A[18][23] * mat_B[23][21] +
                  mat_A[18][24] * mat_B[24][21] +
                  mat_A[18][25] * mat_B[25][21] +
                  mat_A[18][26] * mat_B[26][21] +
                  mat_A[18][27] * mat_B[27][21] +
                  mat_A[18][28] * mat_B[28][21] +
                  mat_A[18][29] * mat_B[29][21] +
                  mat_A[18][30] * mat_B[30][21] +
                  mat_A[18][31] * mat_B[31][21];
    mat_C[18][22] <= 
                  mat_A[18][0] * mat_B[0][22] +
                  mat_A[18][1] * mat_B[1][22] +
                  mat_A[18][2] * mat_B[2][22] +
                  mat_A[18][3] * mat_B[3][22] +
                  mat_A[18][4] * mat_B[4][22] +
                  mat_A[18][5] * mat_B[5][22] +
                  mat_A[18][6] * mat_B[6][22] +
                  mat_A[18][7] * mat_B[7][22] +
                  mat_A[18][8] * mat_B[8][22] +
                  mat_A[18][9] * mat_B[9][22] +
                  mat_A[18][10] * mat_B[10][22] +
                  mat_A[18][11] * mat_B[11][22] +
                  mat_A[18][12] * mat_B[12][22] +
                  mat_A[18][13] * mat_B[13][22] +
                  mat_A[18][14] * mat_B[14][22] +
                  mat_A[18][15] * mat_B[15][22] +
                  mat_A[18][16] * mat_B[16][22] +
                  mat_A[18][17] * mat_B[17][22] +
                  mat_A[18][18] * mat_B[18][22] +
                  mat_A[18][19] * mat_B[19][22] +
                  mat_A[18][20] * mat_B[20][22] +
                  mat_A[18][21] * mat_B[21][22] +
                  mat_A[18][22] * mat_B[22][22] +
                  mat_A[18][23] * mat_B[23][22] +
                  mat_A[18][24] * mat_B[24][22] +
                  mat_A[18][25] * mat_B[25][22] +
                  mat_A[18][26] * mat_B[26][22] +
                  mat_A[18][27] * mat_B[27][22] +
                  mat_A[18][28] * mat_B[28][22] +
                  mat_A[18][29] * mat_B[29][22] +
                  mat_A[18][30] * mat_B[30][22] +
                  mat_A[18][31] * mat_B[31][22];
    mat_C[18][23] <= 
                  mat_A[18][0] * mat_B[0][23] +
                  mat_A[18][1] * mat_B[1][23] +
                  mat_A[18][2] * mat_B[2][23] +
                  mat_A[18][3] * mat_B[3][23] +
                  mat_A[18][4] * mat_B[4][23] +
                  mat_A[18][5] * mat_B[5][23] +
                  mat_A[18][6] * mat_B[6][23] +
                  mat_A[18][7] * mat_B[7][23] +
                  mat_A[18][8] * mat_B[8][23] +
                  mat_A[18][9] * mat_B[9][23] +
                  mat_A[18][10] * mat_B[10][23] +
                  mat_A[18][11] * mat_B[11][23] +
                  mat_A[18][12] * mat_B[12][23] +
                  mat_A[18][13] * mat_B[13][23] +
                  mat_A[18][14] * mat_B[14][23] +
                  mat_A[18][15] * mat_B[15][23] +
                  mat_A[18][16] * mat_B[16][23] +
                  mat_A[18][17] * mat_B[17][23] +
                  mat_A[18][18] * mat_B[18][23] +
                  mat_A[18][19] * mat_B[19][23] +
                  mat_A[18][20] * mat_B[20][23] +
                  mat_A[18][21] * mat_B[21][23] +
                  mat_A[18][22] * mat_B[22][23] +
                  mat_A[18][23] * mat_B[23][23] +
                  mat_A[18][24] * mat_B[24][23] +
                  mat_A[18][25] * mat_B[25][23] +
                  mat_A[18][26] * mat_B[26][23] +
                  mat_A[18][27] * mat_B[27][23] +
                  mat_A[18][28] * mat_B[28][23] +
                  mat_A[18][29] * mat_B[29][23] +
                  mat_A[18][30] * mat_B[30][23] +
                  mat_A[18][31] * mat_B[31][23];
    mat_C[18][24] <= 
                  mat_A[18][0] * mat_B[0][24] +
                  mat_A[18][1] * mat_B[1][24] +
                  mat_A[18][2] * mat_B[2][24] +
                  mat_A[18][3] * mat_B[3][24] +
                  mat_A[18][4] * mat_B[4][24] +
                  mat_A[18][5] * mat_B[5][24] +
                  mat_A[18][6] * mat_B[6][24] +
                  mat_A[18][7] * mat_B[7][24] +
                  mat_A[18][8] * mat_B[8][24] +
                  mat_A[18][9] * mat_B[9][24] +
                  mat_A[18][10] * mat_B[10][24] +
                  mat_A[18][11] * mat_B[11][24] +
                  mat_A[18][12] * mat_B[12][24] +
                  mat_A[18][13] * mat_B[13][24] +
                  mat_A[18][14] * mat_B[14][24] +
                  mat_A[18][15] * mat_B[15][24] +
                  mat_A[18][16] * mat_B[16][24] +
                  mat_A[18][17] * mat_B[17][24] +
                  mat_A[18][18] * mat_B[18][24] +
                  mat_A[18][19] * mat_B[19][24] +
                  mat_A[18][20] * mat_B[20][24] +
                  mat_A[18][21] * mat_B[21][24] +
                  mat_A[18][22] * mat_B[22][24] +
                  mat_A[18][23] * mat_B[23][24] +
                  mat_A[18][24] * mat_B[24][24] +
                  mat_A[18][25] * mat_B[25][24] +
                  mat_A[18][26] * mat_B[26][24] +
                  mat_A[18][27] * mat_B[27][24] +
                  mat_A[18][28] * mat_B[28][24] +
                  mat_A[18][29] * mat_B[29][24] +
                  mat_A[18][30] * mat_B[30][24] +
                  mat_A[18][31] * mat_B[31][24];
    mat_C[18][25] <= 
                  mat_A[18][0] * mat_B[0][25] +
                  mat_A[18][1] * mat_B[1][25] +
                  mat_A[18][2] * mat_B[2][25] +
                  mat_A[18][3] * mat_B[3][25] +
                  mat_A[18][4] * mat_B[4][25] +
                  mat_A[18][5] * mat_B[5][25] +
                  mat_A[18][6] * mat_B[6][25] +
                  mat_A[18][7] * mat_B[7][25] +
                  mat_A[18][8] * mat_B[8][25] +
                  mat_A[18][9] * mat_B[9][25] +
                  mat_A[18][10] * mat_B[10][25] +
                  mat_A[18][11] * mat_B[11][25] +
                  mat_A[18][12] * mat_B[12][25] +
                  mat_A[18][13] * mat_B[13][25] +
                  mat_A[18][14] * mat_B[14][25] +
                  mat_A[18][15] * mat_B[15][25] +
                  mat_A[18][16] * mat_B[16][25] +
                  mat_A[18][17] * mat_B[17][25] +
                  mat_A[18][18] * mat_B[18][25] +
                  mat_A[18][19] * mat_B[19][25] +
                  mat_A[18][20] * mat_B[20][25] +
                  mat_A[18][21] * mat_B[21][25] +
                  mat_A[18][22] * mat_B[22][25] +
                  mat_A[18][23] * mat_B[23][25] +
                  mat_A[18][24] * mat_B[24][25] +
                  mat_A[18][25] * mat_B[25][25] +
                  mat_A[18][26] * mat_B[26][25] +
                  mat_A[18][27] * mat_B[27][25] +
                  mat_A[18][28] * mat_B[28][25] +
                  mat_A[18][29] * mat_B[29][25] +
                  mat_A[18][30] * mat_B[30][25] +
                  mat_A[18][31] * mat_B[31][25];
    mat_C[18][26] <= 
                  mat_A[18][0] * mat_B[0][26] +
                  mat_A[18][1] * mat_B[1][26] +
                  mat_A[18][2] * mat_B[2][26] +
                  mat_A[18][3] * mat_B[3][26] +
                  mat_A[18][4] * mat_B[4][26] +
                  mat_A[18][5] * mat_B[5][26] +
                  mat_A[18][6] * mat_B[6][26] +
                  mat_A[18][7] * mat_B[7][26] +
                  mat_A[18][8] * mat_B[8][26] +
                  mat_A[18][9] * mat_B[9][26] +
                  mat_A[18][10] * mat_B[10][26] +
                  mat_A[18][11] * mat_B[11][26] +
                  mat_A[18][12] * mat_B[12][26] +
                  mat_A[18][13] * mat_B[13][26] +
                  mat_A[18][14] * mat_B[14][26] +
                  mat_A[18][15] * mat_B[15][26] +
                  mat_A[18][16] * mat_B[16][26] +
                  mat_A[18][17] * mat_B[17][26] +
                  mat_A[18][18] * mat_B[18][26] +
                  mat_A[18][19] * mat_B[19][26] +
                  mat_A[18][20] * mat_B[20][26] +
                  mat_A[18][21] * mat_B[21][26] +
                  mat_A[18][22] * mat_B[22][26] +
                  mat_A[18][23] * mat_B[23][26] +
                  mat_A[18][24] * mat_B[24][26] +
                  mat_A[18][25] * mat_B[25][26] +
                  mat_A[18][26] * mat_B[26][26] +
                  mat_A[18][27] * mat_B[27][26] +
                  mat_A[18][28] * mat_B[28][26] +
                  mat_A[18][29] * mat_B[29][26] +
                  mat_A[18][30] * mat_B[30][26] +
                  mat_A[18][31] * mat_B[31][26];
    mat_C[18][27] <= 
                  mat_A[18][0] * mat_B[0][27] +
                  mat_A[18][1] * mat_B[1][27] +
                  mat_A[18][2] * mat_B[2][27] +
                  mat_A[18][3] * mat_B[3][27] +
                  mat_A[18][4] * mat_B[4][27] +
                  mat_A[18][5] * mat_B[5][27] +
                  mat_A[18][6] * mat_B[6][27] +
                  mat_A[18][7] * mat_B[7][27] +
                  mat_A[18][8] * mat_B[8][27] +
                  mat_A[18][9] * mat_B[9][27] +
                  mat_A[18][10] * mat_B[10][27] +
                  mat_A[18][11] * mat_B[11][27] +
                  mat_A[18][12] * mat_B[12][27] +
                  mat_A[18][13] * mat_B[13][27] +
                  mat_A[18][14] * mat_B[14][27] +
                  mat_A[18][15] * mat_B[15][27] +
                  mat_A[18][16] * mat_B[16][27] +
                  mat_A[18][17] * mat_B[17][27] +
                  mat_A[18][18] * mat_B[18][27] +
                  mat_A[18][19] * mat_B[19][27] +
                  mat_A[18][20] * mat_B[20][27] +
                  mat_A[18][21] * mat_B[21][27] +
                  mat_A[18][22] * mat_B[22][27] +
                  mat_A[18][23] * mat_B[23][27] +
                  mat_A[18][24] * mat_B[24][27] +
                  mat_A[18][25] * mat_B[25][27] +
                  mat_A[18][26] * mat_B[26][27] +
                  mat_A[18][27] * mat_B[27][27] +
                  mat_A[18][28] * mat_B[28][27] +
                  mat_A[18][29] * mat_B[29][27] +
                  mat_A[18][30] * mat_B[30][27] +
                  mat_A[18][31] * mat_B[31][27];
    mat_C[18][28] <= 
                  mat_A[18][0] * mat_B[0][28] +
                  mat_A[18][1] * mat_B[1][28] +
                  mat_A[18][2] * mat_B[2][28] +
                  mat_A[18][3] * mat_B[3][28] +
                  mat_A[18][4] * mat_B[4][28] +
                  mat_A[18][5] * mat_B[5][28] +
                  mat_A[18][6] * mat_B[6][28] +
                  mat_A[18][7] * mat_B[7][28] +
                  mat_A[18][8] * mat_B[8][28] +
                  mat_A[18][9] * mat_B[9][28] +
                  mat_A[18][10] * mat_B[10][28] +
                  mat_A[18][11] * mat_B[11][28] +
                  mat_A[18][12] * mat_B[12][28] +
                  mat_A[18][13] * mat_B[13][28] +
                  mat_A[18][14] * mat_B[14][28] +
                  mat_A[18][15] * mat_B[15][28] +
                  mat_A[18][16] * mat_B[16][28] +
                  mat_A[18][17] * mat_B[17][28] +
                  mat_A[18][18] * mat_B[18][28] +
                  mat_A[18][19] * mat_B[19][28] +
                  mat_A[18][20] * mat_B[20][28] +
                  mat_A[18][21] * mat_B[21][28] +
                  mat_A[18][22] * mat_B[22][28] +
                  mat_A[18][23] * mat_B[23][28] +
                  mat_A[18][24] * mat_B[24][28] +
                  mat_A[18][25] * mat_B[25][28] +
                  mat_A[18][26] * mat_B[26][28] +
                  mat_A[18][27] * mat_B[27][28] +
                  mat_A[18][28] * mat_B[28][28] +
                  mat_A[18][29] * mat_B[29][28] +
                  mat_A[18][30] * mat_B[30][28] +
                  mat_A[18][31] * mat_B[31][28];
    mat_C[18][29] <= 
                  mat_A[18][0] * mat_B[0][29] +
                  mat_A[18][1] * mat_B[1][29] +
                  mat_A[18][2] * mat_B[2][29] +
                  mat_A[18][3] * mat_B[3][29] +
                  mat_A[18][4] * mat_B[4][29] +
                  mat_A[18][5] * mat_B[5][29] +
                  mat_A[18][6] * mat_B[6][29] +
                  mat_A[18][7] * mat_B[7][29] +
                  mat_A[18][8] * mat_B[8][29] +
                  mat_A[18][9] * mat_B[9][29] +
                  mat_A[18][10] * mat_B[10][29] +
                  mat_A[18][11] * mat_B[11][29] +
                  mat_A[18][12] * mat_B[12][29] +
                  mat_A[18][13] * mat_B[13][29] +
                  mat_A[18][14] * mat_B[14][29] +
                  mat_A[18][15] * mat_B[15][29] +
                  mat_A[18][16] * mat_B[16][29] +
                  mat_A[18][17] * mat_B[17][29] +
                  mat_A[18][18] * mat_B[18][29] +
                  mat_A[18][19] * mat_B[19][29] +
                  mat_A[18][20] * mat_B[20][29] +
                  mat_A[18][21] * mat_B[21][29] +
                  mat_A[18][22] * mat_B[22][29] +
                  mat_A[18][23] * mat_B[23][29] +
                  mat_A[18][24] * mat_B[24][29] +
                  mat_A[18][25] * mat_B[25][29] +
                  mat_A[18][26] * mat_B[26][29] +
                  mat_A[18][27] * mat_B[27][29] +
                  mat_A[18][28] * mat_B[28][29] +
                  mat_A[18][29] * mat_B[29][29] +
                  mat_A[18][30] * mat_B[30][29] +
                  mat_A[18][31] * mat_B[31][29];
    mat_C[18][30] <= 
                  mat_A[18][0] * mat_B[0][30] +
                  mat_A[18][1] * mat_B[1][30] +
                  mat_A[18][2] * mat_B[2][30] +
                  mat_A[18][3] * mat_B[3][30] +
                  mat_A[18][4] * mat_B[4][30] +
                  mat_A[18][5] * mat_B[5][30] +
                  mat_A[18][6] * mat_B[6][30] +
                  mat_A[18][7] * mat_B[7][30] +
                  mat_A[18][8] * mat_B[8][30] +
                  mat_A[18][9] * mat_B[9][30] +
                  mat_A[18][10] * mat_B[10][30] +
                  mat_A[18][11] * mat_B[11][30] +
                  mat_A[18][12] * mat_B[12][30] +
                  mat_A[18][13] * mat_B[13][30] +
                  mat_A[18][14] * mat_B[14][30] +
                  mat_A[18][15] * mat_B[15][30] +
                  mat_A[18][16] * mat_B[16][30] +
                  mat_A[18][17] * mat_B[17][30] +
                  mat_A[18][18] * mat_B[18][30] +
                  mat_A[18][19] * mat_B[19][30] +
                  mat_A[18][20] * mat_B[20][30] +
                  mat_A[18][21] * mat_B[21][30] +
                  mat_A[18][22] * mat_B[22][30] +
                  mat_A[18][23] * mat_B[23][30] +
                  mat_A[18][24] * mat_B[24][30] +
                  mat_A[18][25] * mat_B[25][30] +
                  mat_A[18][26] * mat_B[26][30] +
                  mat_A[18][27] * mat_B[27][30] +
                  mat_A[18][28] * mat_B[28][30] +
                  mat_A[18][29] * mat_B[29][30] +
                  mat_A[18][30] * mat_B[30][30] +
                  mat_A[18][31] * mat_B[31][30];
    mat_C[18][31] <= 
                  mat_A[18][0] * mat_B[0][31] +
                  mat_A[18][1] * mat_B[1][31] +
                  mat_A[18][2] * mat_B[2][31] +
                  mat_A[18][3] * mat_B[3][31] +
                  mat_A[18][4] * mat_B[4][31] +
                  mat_A[18][5] * mat_B[5][31] +
                  mat_A[18][6] * mat_B[6][31] +
                  mat_A[18][7] * mat_B[7][31] +
                  mat_A[18][8] * mat_B[8][31] +
                  mat_A[18][9] * mat_B[9][31] +
                  mat_A[18][10] * mat_B[10][31] +
                  mat_A[18][11] * mat_B[11][31] +
                  mat_A[18][12] * mat_B[12][31] +
                  mat_A[18][13] * mat_B[13][31] +
                  mat_A[18][14] * mat_B[14][31] +
                  mat_A[18][15] * mat_B[15][31] +
                  mat_A[18][16] * mat_B[16][31] +
                  mat_A[18][17] * mat_B[17][31] +
                  mat_A[18][18] * mat_B[18][31] +
                  mat_A[18][19] * mat_B[19][31] +
                  mat_A[18][20] * mat_B[20][31] +
                  mat_A[18][21] * mat_B[21][31] +
                  mat_A[18][22] * mat_B[22][31] +
                  mat_A[18][23] * mat_B[23][31] +
                  mat_A[18][24] * mat_B[24][31] +
                  mat_A[18][25] * mat_B[25][31] +
                  mat_A[18][26] * mat_B[26][31] +
                  mat_A[18][27] * mat_B[27][31] +
                  mat_A[18][28] * mat_B[28][31] +
                  mat_A[18][29] * mat_B[29][31] +
                  mat_A[18][30] * mat_B[30][31] +
                  mat_A[18][31] * mat_B[31][31];
    mat_C[19][0] <= 
                  mat_A[19][0] * mat_B[0][0] +
                  mat_A[19][1] * mat_B[1][0] +
                  mat_A[19][2] * mat_B[2][0] +
                  mat_A[19][3] * mat_B[3][0] +
                  mat_A[19][4] * mat_B[4][0] +
                  mat_A[19][5] * mat_B[5][0] +
                  mat_A[19][6] * mat_B[6][0] +
                  mat_A[19][7] * mat_B[7][0] +
                  mat_A[19][8] * mat_B[8][0] +
                  mat_A[19][9] * mat_B[9][0] +
                  mat_A[19][10] * mat_B[10][0] +
                  mat_A[19][11] * mat_B[11][0] +
                  mat_A[19][12] * mat_B[12][0] +
                  mat_A[19][13] * mat_B[13][0] +
                  mat_A[19][14] * mat_B[14][0] +
                  mat_A[19][15] * mat_B[15][0] +
                  mat_A[19][16] * mat_B[16][0] +
                  mat_A[19][17] * mat_B[17][0] +
                  mat_A[19][18] * mat_B[18][0] +
                  mat_A[19][19] * mat_B[19][0] +
                  mat_A[19][20] * mat_B[20][0] +
                  mat_A[19][21] * mat_B[21][0] +
                  mat_A[19][22] * mat_B[22][0] +
                  mat_A[19][23] * mat_B[23][0] +
                  mat_A[19][24] * mat_B[24][0] +
                  mat_A[19][25] * mat_B[25][0] +
                  mat_A[19][26] * mat_B[26][0] +
                  mat_A[19][27] * mat_B[27][0] +
                  mat_A[19][28] * mat_B[28][0] +
                  mat_A[19][29] * mat_B[29][0] +
                  mat_A[19][30] * mat_B[30][0] +
                  mat_A[19][31] * mat_B[31][0];
    mat_C[19][1] <= 
                  mat_A[19][0] * mat_B[0][1] +
                  mat_A[19][1] * mat_B[1][1] +
                  mat_A[19][2] * mat_B[2][1] +
                  mat_A[19][3] * mat_B[3][1] +
                  mat_A[19][4] * mat_B[4][1] +
                  mat_A[19][5] * mat_B[5][1] +
                  mat_A[19][6] * mat_B[6][1] +
                  mat_A[19][7] * mat_B[7][1] +
                  mat_A[19][8] * mat_B[8][1] +
                  mat_A[19][9] * mat_B[9][1] +
                  mat_A[19][10] * mat_B[10][1] +
                  mat_A[19][11] * mat_B[11][1] +
                  mat_A[19][12] * mat_B[12][1] +
                  mat_A[19][13] * mat_B[13][1] +
                  mat_A[19][14] * mat_B[14][1] +
                  mat_A[19][15] * mat_B[15][1] +
                  mat_A[19][16] * mat_B[16][1] +
                  mat_A[19][17] * mat_B[17][1] +
                  mat_A[19][18] * mat_B[18][1] +
                  mat_A[19][19] * mat_B[19][1] +
                  mat_A[19][20] * mat_B[20][1] +
                  mat_A[19][21] * mat_B[21][1] +
                  mat_A[19][22] * mat_B[22][1] +
                  mat_A[19][23] * mat_B[23][1] +
                  mat_A[19][24] * mat_B[24][1] +
                  mat_A[19][25] * mat_B[25][1] +
                  mat_A[19][26] * mat_B[26][1] +
                  mat_A[19][27] * mat_B[27][1] +
                  mat_A[19][28] * mat_B[28][1] +
                  mat_A[19][29] * mat_B[29][1] +
                  mat_A[19][30] * mat_B[30][1] +
                  mat_A[19][31] * mat_B[31][1];
    mat_C[19][2] <= 
                  mat_A[19][0] * mat_B[0][2] +
                  mat_A[19][1] * mat_B[1][2] +
                  mat_A[19][2] * mat_B[2][2] +
                  mat_A[19][3] * mat_B[3][2] +
                  mat_A[19][4] * mat_B[4][2] +
                  mat_A[19][5] * mat_B[5][2] +
                  mat_A[19][6] * mat_B[6][2] +
                  mat_A[19][7] * mat_B[7][2] +
                  mat_A[19][8] * mat_B[8][2] +
                  mat_A[19][9] * mat_B[9][2] +
                  mat_A[19][10] * mat_B[10][2] +
                  mat_A[19][11] * mat_B[11][2] +
                  mat_A[19][12] * mat_B[12][2] +
                  mat_A[19][13] * mat_B[13][2] +
                  mat_A[19][14] * mat_B[14][2] +
                  mat_A[19][15] * mat_B[15][2] +
                  mat_A[19][16] * mat_B[16][2] +
                  mat_A[19][17] * mat_B[17][2] +
                  mat_A[19][18] * mat_B[18][2] +
                  mat_A[19][19] * mat_B[19][2] +
                  mat_A[19][20] * mat_B[20][2] +
                  mat_A[19][21] * mat_B[21][2] +
                  mat_A[19][22] * mat_B[22][2] +
                  mat_A[19][23] * mat_B[23][2] +
                  mat_A[19][24] * mat_B[24][2] +
                  mat_A[19][25] * mat_B[25][2] +
                  mat_A[19][26] * mat_B[26][2] +
                  mat_A[19][27] * mat_B[27][2] +
                  mat_A[19][28] * mat_B[28][2] +
                  mat_A[19][29] * mat_B[29][2] +
                  mat_A[19][30] * mat_B[30][2] +
                  mat_A[19][31] * mat_B[31][2];
    mat_C[19][3] <= 
                  mat_A[19][0] * mat_B[0][3] +
                  mat_A[19][1] * mat_B[1][3] +
                  mat_A[19][2] * mat_B[2][3] +
                  mat_A[19][3] * mat_B[3][3] +
                  mat_A[19][4] * mat_B[4][3] +
                  mat_A[19][5] * mat_B[5][3] +
                  mat_A[19][6] * mat_B[6][3] +
                  mat_A[19][7] * mat_B[7][3] +
                  mat_A[19][8] * mat_B[8][3] +
                  mat_A[19][9] * mat_B[9][3] +
                  mat_A[19][10] * mat_B[10][3] +
                  mat_A[19][11] * mat_B[11][3] +
                  mat_A[19][12] * mat_B[12][3] +
                  mat_A[19][13] * mat_B[13][3] +
                  mat_A[19][14] * mat_B[14][3] +
                  mat_A[19][15] * mat_B[15][3] +
                  mat_A[19][16] * mat_B[16][3] +
                  mat_A[19][17] * mat_B[17][3] +
                  mat_A[19][18] * mat_B[18][3] +
                  mat_A[19][19] * mat_B[19][3] +
                  mat_A[19][20] * mat_B[20][3] +
                  mat_A[19][21] * mat_B[21][3] +
                  mat_A[19][22] * mat_B[22][3] +
                  mat_A[19][23] * mat_B[23][3] +
                  mat_A[19][24] * mat_B[24][3] +
                  mat_A[19][25] * mat_B[25][3] +
                  mat_A[19][26] * mat_B[26][3] +
                  mat_A[19][27] * mat_B[27][3] +
                  mat_A[19][28] * mat_B[28][3] +
                  mat_A[19][29] * mat_B[29][3] +
                  mat_A[19][30] * mat_B[30][3] +
                  mat_A[19][31] * mat_B[31][3];
    mat_C[19][4] <= 
                  mat_A[19][0] * mat_B[0][4] +
                  mat_A[19][1] * mat_B[1][4] +
                  mat_A[19][2] * mat_B[2][4] +
                  mat_A[19][3] * mat_B[3][4] +
                  mat_A[19][4] * mat_B[4][4] +
                  mat_A[19][5] * mat_B[5][4] +
                  mat_A[19][6] * mat_B[6][4] +
                  mat_A[19][7] * mat_B[7][4] +
                  mat_A[19][8] * mat_B[8][4] +
                  mat_A[19][9] * mat_B[9][4] +
                  mat_A[19][10] * mat_B[10][4] +
                  mat_A[19][11] * mat_B[11][4] +
                  mat_A[19][12] * mat_B[12][4] +
                  mat_A[19][13] * mat_B[13][4] +
                  mat_A[19][14] * mat_B[14][4] +
                  mat_A[19][15] * mat_B[15][4] +
                  mat_A[19][16] * mat_B[16][4] +
                  mat_A[19][17] * mat_B[17][4] +
                  mat_A[19][18] * mat_B[18][4] +
                  mat_A[19][19] * mat_B[19][4] +
                  mat_A[19][20] * mat_B[20][4] +
                  mat_A[19][21] * mat_B[21][4] +
                  mat_A[19][22] * mat_B[22][4] +
                  mat_A[19][23] * mat_B[23][4] +
                  mat_A[19][24] * mat_B[24][4] +
                  mat_A[19][25] * mat_B[25][4] +
                  mat_A[19][26] * mat_B[26][4] +
                  mat_A[19][27] * mat_B[27][4] +
                  mat_A[19][28] * mat_B[28][4] +
                  mat_A[19][29] * mat_B[29][4] +
                  mat_A[19][30] * mat_B[30][4] +
                  mat_A[19][31] * mat_B[31][4];
    mat_C[19][5] <= 
                  mat_A[19][0] * mat_B[0][5] +
                  mat_A[19][1] * mat_B[1][5] +
                  mat_A[19][2] * mat_B[2][5] +
                  mat_A[19][3] * mat_B[3][5] +
                  mat_A[19][4] * mat_B[4][5] +
                  mat_A[19][5] * mat_B[5][5] +
                  mat_A[19][6] * mat_B[6][5] +
                  mat_A[19][7] * mat_B[7][5] +
                  mat_A[19][8] * mat_B[8][5] +
                  mat_A[19][9] * mat_B[9][5] +
                  mat_A[19][10] * mat_B[10][5] +
                  mat_A[19][11] * mat_B[11][5] +
                  mat_A[19][12] * mat_B[12][5] +
                  mat_A[19][13] * mat_B[13][5] +
                  mat_A[19][14] * mat_B[14][5] +
                  mat_A[19][15] * mat_B[15][5] +
                  mat_A[19][16] * mat_B[16][5] +
                  mat_A[19][17] * mat_B[17][5] +
                  mat_A[19][18] * mat_B[18][5] +
                  mat_A[19][19] * mat_B[19][5] +
                  mat_A[19][20] * mat_B[20][5] +
                  mat_A[19][21] * mat_B[21][5] +
                  mat_A[19][22] * mat_B[22][5] +
                  mat_A[19][23] * mat_B[23][5] +
                  mat_A[19][24] * mat_B[24][5] +
                  mat_A[19][25] * mat_B[25][5] +
                  mat_A[19][26] * mat_B[26][5] +
                  mat_A[19][27] * mat_B[27][5] +
                  mat_A[19][28] * mat_B[28][5] +
                  mat_A[19][29] * mat_B[29][5] +
                  mat_A[19][30] * mat_B[30][5] +
                  mat_A[19][31] * mat_B[31][5];
    mat_C[19][6] <= 
                  mat_A[19][0] * mat_B[0][6] +
                  mat_A[19][1] * mat_B[1][6] +
                  mat_A[19][2] * mat_B[2][6] +
                  mat_A[19][3] * mat_B[3][6] +
                  mat_A[19][4] * mat_B[4][6] +
                  mat_A[19][5] * mat_B[5][6] +
                  mat_A[19][6] * mat_B[6][6] +
                  mat_A[19][7] * mat_B[7][6] +
                  mat_A[19][8] * mat_B[8][6] +
                  mat_A[19][9] * mat_B[9][6] +
                  mat_A[19][10] * mat_B[10][6] +
                  mat_A[19][11] * mat_B[11][6] +
                  mat_A[19][12] * mat_B[12][6] +
                  mat_A[19][13] * mat_B[13][6] +
                  mat_A[19][14] * mat_B[14][6] +
                  mat_A[19][15] * mat_B[15][6] +
                  mat_A[19][16] * mat_B[16][6] +
                  mat_A[19][17] * mat_B[17][6] +
                  mat_A[19][18] * mat_B[18][6] +
                  mat_A[19][19] * mat_B[19][6] +
                  mat_A[19][20] * mat_B[20][6] +
                  mat_A[19][21] * mat_B[21][6] +
                  mat_A[19][22] * mat_B[22][6] +
                  mat_A[19][23] * mat_B[23][6] +
                  mat_A[19][24] * mat_B[24][6] +
                  mat_A[19][25] * mat_B[25][6] +
                  mat_A[19][26] * mat_B[26][6] +
                  mat_A[19][27] * mat_B[27][6] +
                  mat_A[19][28] * mat_B[28][6] +
                  mat_A[19][29] * mat_B[29][6] +
                  mat_A[19][30] * mat_B[30][6] +
                  mat_A[19][31] * mat_B[31][6];
    mat_C[19][7] <= 
                  mat_A[19][0] * mat_B[0][7] +
                  mat_A[19][1] * mat_B[1][7] +
                  mat_A[19][2] * mat_B[2][7] +
                  mat_A[19][3] * mat_B[3][7] +
                  mat_A[19][4] * mat_B[4][7] +
                  mat_A[19][5] * mat_B[5][7] +
                  mat_A[19][6] * mat_B[6][7] +
                  mat_A[19][7] * mat_B[7][7] +
                  mat_A[19][8] * mat_B[8][7] +
                  mat_A[19][9] * mat_B[9][7] +
                  mat_A[19][10] * mat_B[10][7] +
                  mat_A[19][11] * mat_B[11][7] +
                  mat_A[19][12] * mat_B[12][7] +
                  mat_A[19][13] * mat_B[13][7] +
                  mat_A[19][14] * mat_B[14][7] +
                  mat_A[19][15] * mat_B[15][7] +
                  mat_A[19][16] * mat_B[16][7] +
                  mat_A[19][17] * mat_B[17][7] +
                  mat_A[19][18] * mat_B[18][7] +
                  mat_A[19][19] * mat_B[19][7] +
                  mat_A[19][20] * mat_B[20][7] +
                  mat_A[19][21] * mat_B[21][7] +
                  mat_A[19][22] * mat_B[22][7] +
                  mat_A[19][23] * mat_B[23][7] +
                  mat_A[19][24] * mat_B[24][7] +
                  mat_A[19][25] * mat_B[25][7] +
                  mat_A[19][26] * mat_B[26][7] +
                  mat_A[19][27] * mat_B[27][7] +
                  mat_A[19][28] * mat_B[28][7] +
                  mat_A[19][29] * mat_B[29][7] +
                  mat_A[19][30] * mat_B[30][7] +
                  mat_A[19][31] * mat_B[31][7];
    mat_C[19][8] <= 
                  mat_A[19][0] * mat_B[0][8] +
                  mat_A[19][1] * mat_B[1][8] +
                  mat_A[19][2] * mat_B[2][8] +
                  mat_A[19][3] * mat_B[3][8] +
                  mat_A[19][4] * mat_B[4][8] +
                  mat_A[19][5] * mat_B[5][8] +
                  mat_A[19][6] * mat_B[6][8] +
                  mat_A[19][7] * mat_B[7][8] +
                  mat_A[19][8] * mat_B[8][8] +
                  mat_A[19][9] * mat_B[9][8] +
                  mat_A[19][10] * mat_B[10][8] +
                  mat_A[19][11] * mat_B[11][8] +
                  mat_A[19][12] * mat_B[12][8] +
                  mat_A[19][13] * mat_B[13][8] +
                  mat_A[19][14] * mat_B[14][8] +
                  mat_A[19][15] * mat_B[15][8] +
                  mat_A[19][16] * mat_B[16][8] +
                  mat_A[19][17] * mat_B[17][8] +
                  mat_A[19][18] * mat_B[18][8] +
                  mat_A[19][19] * mat_B[19][8] +
                  mat_A[19][20] * mat_B[20][8] +
                  mat_A[19][21] * mat_B[21][8] +
                  mat_A[19][22] * mat_B[22][8] +
                  mat_A[19][23] * mat_B[23][8] +
                  mat_A[19][24] * mat_B[24][8] +
                  mat_A[19][25] * mat_B[25][8] +
                  mat_A[19][26] * mat_B[26][8] +
                  mat_A[19][27] * mat_B[27][8] +
                  mat_A[19][28] * mat_B[28][8] +
                  mat_A[19][29] * mat_B[29][8] +
                  mat_A[19][30] * mat_B[30][8] +
                  mat_A[19][31] * mat_B[31][8];
    mat_C[19][9] <= 
                  mat_A[19][0] * mat_B[0][9] +
                  mat_A[19][1] * mat_B[1][9] +
                  mat_A[19][2] * mat_B[2][9] +
                  mat_A[19][3] * mat_B[3][9] +
                  mat_A[19][4] * mat_B[4][9] +
                  mat_A[19][5] * mat_B[5][9] +
                  mat_A[19][6] * mat_B[6][9] +
                  mat_A[19][7] * mat_B[7][9] +
                  mat_A[19][8] * mat_B[8][9] +
                  mat_A[19][9] * mat_B[9][9] +
                  mat_A[19][10] * mat_B[10][9] +
                  mat_A[19][11] * mat_B[11][9] +
                  mat_A[19][12] * mat_B[12][9] +
                  mat_A[19][13] * mat_B[13][9] +
                  mat_A[19][14] * mat_B[14][9] +
                  mat_A[19][15] * mat_B[15][9] +
                  mat_A[19][16] * mat_B[16][9] +
                  mat_A[19][17] * mat_B[17][9] +
                  mat_A[19][18] * mat_B[18][9] +
                  mat_A[19][19] * mat_B[19][9] +
                  mat_A[19][20] * mat_B[20][9] +
                  mat_A[19][21] * mat_B[21][9] +
                  mat_A[19][22] * mat_B[22][9] +
                  mat_A[19][23] * mat_B[23][9] +
                  mat_A[19][24] * mat_B[24][9] +
                  mat_A[19][25] * mat_B[25][9] +
                  mat_A[19][26] * mat_B[26][9] +
                  mat_A[19][27] * mat_B[27][9] +
                  mat_A[19][28] * mat_B[28][9] +
                  mat_A[19][29] * mat_B[29][9] +
                  mat_A[19][30] * mat_B[30][9] +
                  mat_A[19][31] * mat_B[31][9];
    mat_C[19][10] <= 
                  mat_A[19][0] * mat_B[0][10] +
                  mat_A[19][1] * mat_B[1][10] +
                  mat_A[19][2] * mat_B[2][10] +
                  mat_A[19][3] * mat_B[3][10] +
                  mat_A[19][4] * mat_B[4][10] +
                  mat_A[19][5] * mat_B[5][10] +
                  mat_A[19][6] * mat_B[6][10] +
                  mat_A[19][7] * mat_B[7][10] +
                  mat_A[19][8] * mat_B[8][10] +
                  mat_A[19][9] * mat_B[9][10] +
                  mat_A[19][10] * mat_B[10][10] +
                  mat_A[19][11] * mat_B[11][10] +
                  mat_A[19][12] * mat_B[12][10] +
                  mat_A[19][13] * mat_B[13][10] +
                  mat_A[19][14] * mat_B[14][10] +
                  mat_A[19][15] * mat_B[15][10] +
                  mat_A[19][16] * mat_B[16][10] +
                  mat_A[19][17] * mat_B[17][10] +
                  mat_A[19][18] * mat_B[18][10] +
                  mat_A[19][19] * mat_B[19][10] +
                  mat_A[19][20] * mat_B[20][10] +
                  mat_A[19][21] * mat_B[21][10] +
                  mat_A[19][22] * mat_B[22][10] +
                  mat_A[19][23] * mat_B[23][10] +
                  mat_A[19][24] * mat_B[24][10] +
                  mat_A[19][25] * mat_B[25][10] +
                  mat_A[19][26] * mat_B[26][10] +
                  mat_A[19][27] * mat_B[27][10] +
                  mat_A[19][28] * mat_B[28][10] +
                  mat_A[19][29] * mat_B[29][10] +
                  mat_A[19][30] * mat_B[30][10] +
                  mat_A[19][31] * mat_B[31][10];
    mat_C[19][11] <= 
                  mat_A[19][0] * mat_B[0][11] +
                  mat_A[19][1] * mat_B[1][11] +
                  mat_A[19][2] * mat_B[2][11] +
                  mat_A[19][3] * mat_B[3][11] +
                  mat_A[19][4] * mat_B[4][11] +
                  mat_A[19][5] * mat_B[5][11] +
                  mat_A[19][6] * mat_B[6][11] +
                  mat_A[19][7] * mat_B[7][11] +
                  mat_A[19][8] * mat_B[8][11] +
                  mat_A[19][9] * mat_B[9][11] +
                  mat_A[19][10] * mat_B[10][11] +
                  mat_A[19][11] * mat_B[11][11] +
                  mat_A[19][12] * mat_B[12][11] +
                  mat_A[19][13] * mat_B[13][11] +
                  mat_A[19][14] * mat_B[14][11] +
                  mat_A[19][15] * mat_B[15][11] +
                  mat_A[19][16] * mat_B[16][11] +
                  mat_A[19][17] * mat_B[17][11] +
                  mat_A[19][18] * mat_B[18][11] +
                  mat_A[19][19] * mat_B[19][11] +
                  mat_A[19][20] * mat_B[20][11] +
                  mat_A[19][21] * mat_B[21][11] +
                  mat_A[19][22] * mat_B[22][11] +
                  mat_A[19][23] * mat_B[23][11] +
                  mat_A[19][24] * mat_B[24][11] +
                  mat_A[19][25] * mat_B[25][11] +
                  mat_A[19][26] * mat_B[26][11] +
                  mat_A[19][27] * mat_B[27][11] +
                  mat_A[19][28] * mat_B[28][11] +
                  mat_A[19][29] * mat_B[29][11] +
                  mat_A[19][30] * mat_B[30][11] +
                  mat_A[19][31] * mat_B[31][11];
    mat_C[19][12] <= 
                  mat_A[19][0] * mat_B[0][12] +
                  mat_A[19][1] * mat_B[1][12] +
                  mat_A[19][2] * mat_B[2][12] +
                  mat_A[19][3] * mat_B[3][12] +
                  mat_A[19][4] * mat_B[4][12] +
                  mat_A[19][5] * mat_B[5][12] +
                  mat_A[19][6] * mat_B[6][12] +
                  mat_A[19][7] * mat_B[7][12] +
                  mat_A[19][8] * mat_B[8][12] +
                  mat_A[19][9] * mat_B[9][12] +
                  mat_A[19][10] * mat_B[10][12] +
                  mat_A[19][11] * mat_B[11][12] +
                  mat_A[19][12] * mat_B[12][12] +
                  mat_A[19][13] * mat_B[13][12] +
                  mat_A[19][14] * mat_B[14][12] +
                  mat_A[19][15] * mat_B[15][12] +
                  mat_A[19][16] * mat_B[16][12] +
                  mat_A[19][17] * mat_B[17][12] +
                  mat_A[19][18] * mat_B[18][12] +
                  mat_A[19][19] * mat_B[19][12] +
                  mat_A[19][20] * mat_B[20][12] +
                  mat_A[19][21] * mat_B[21][12] +
                  mat_A[19][22] * mat_B[22][12] +
                  mat_A[19][23] * mat_B[23][12] +
                  mat_A[19][24] * mat_B[24][12] +
                  mat_A[19][25] * mat_B[25][12] +
                  mat_A[19][26] * mat_B[26][12] +
                  mat_A[19][27] * mat_B[27][12] +
                  mat_A[19][28] * mat_B[28][12] +
                  mat_A[19][29] * mat_B[29][12] +
                  mat_A[19][30] * mat_B[30][12] +
                  mat_A[19][31] * mat_B[31][12];
    mat_C[19][13] <= 
                  mat_A[19][0] * mat_B[0][13] +
                  mat_A[19][1] * mat_B[1][13] +
                  mat_A[19][2] * mat_B[2][13] +
                  mat_A[19][3] * mat_B[3][13] +
                  mat_A[19][4] * mat_B[4][13] +
                  mat_A[19][5] * mat_B[5][13] +
                  mat_A[19][6] * mat_B[6][13] +
                  mat_A[19][7] * mat_B[7][13] +
                  mat_A[19][8] * mat_B[8][13] +
                  mat_A[19][9] * mat_B[9][13] +
                  mat_A[19][10] * mat_B[10][13] +
                  mat_A[19][11] * mat_B[11][13] +
                  mat_A[19][12] * mat_B[12][13] +
                  mat_A[19][13] * mat_B[13][13] +
                  mat_A[19][14] * mat_B[14][13] +
                  mat_A[19][15] * mat_B[15][13] +
                  mat_A[19][16] * mat_B[16][13] +
                  mat_A[19][17] * mat_B[17][13] +
                  mat_A[19][18] * mat_B[18][13] +
                  mat_A[19][19] * mat_B[19][13] +
                  mat_A[19][20] * mat_B[20][13] +
                  mat_A[19][21] * mat_B[21][13] +
                  mat_A[19][22] * mat_B[22][13] +
                  mat_A[19][23] * mat_B[23][13] +
                  mat_A[19][24] * mat_B[24][13] +
                  mat_A[19][25] * mat_B[25][13] +
                  mat_A[19][26] * mat_B[26][13] +
                  mat_A[19][27] * mat_B[27][13] +
                  mat_A[19][28] * mat_B[28][13] +
                  mat_A[19][29] * mat_B[29][13] +
                  mat_A[19][30] * mat_B[30][13] +
                  mat_A[19][31] * mat_B[31][13];
    mat_C[19][14] <= 
                  mat_A[19][0] * mat_B[0][14] +
                  mat_A[19][1] * mat_B[1][14] +
                  mat_A[19][2] * mat_B[2][14] +
                  mat_A[19][3] * mat_B[3][14] +
                  mat_A[19][4] * mat_B[4][14] +
                  mat_A[19][5] * mat_B[5][14] +
                  mat_A[19][6] * mat_B[6][14] +
                  mat_A[19][7] * mat_B[7][14] +
                  mat_A[19][8] * mat_B[8][14] +
                  mat_A[19][9] * mat_B[9][14] +
                  mat_A[19][10] * mat_B[10][14] +
                  mat_A[19][11] * mat_B[11][14] +
                  mat_A[19][12] * mat_B[12][14] +
                  mat_A[19][13] * mat_B[13][14] +
                  mat_A[19][14] * mat_B[14][14] +
                  mat_A[19][15] * mat_B[15][14] +
                  mat_A[19][16] * mat_B[16][14] +
                  mat_A[19][17] * mat_B[17][14] +
                  mat_A[19][18] * mat_B[18][14] +
                  mat_A[19][19] * mat_B[19][14] +
                  mat_A[19][20] * mat_B[20][14] +
                  mat_A[19][21] * mat_B[21][14] +
                  mat_A[19][22] * mat_B[22][14] +
                  mat_A[19][23] * mat_B[23][14] +
                  mat_A[19][24] * mat_B[24][14] +
                  mat_A[19][25] * mat_B[25][14] +
                  mat_A[19][26] * mat_B[26][14] +
                  mat_A[19][27] * mat_B[27][14] +
                  mat_A[19][28] * mat_B[28][14] +
                  mat_A[19][29] * mat_B[29][14] +
                  mat_A[19][30] * mat_B[30][14] +
                  mat_A[19][31] * mat_B[31][14];
    mat_C[19][15] <= 
                  mat_A[19][0] * mat_B[0][15] +
                  mat_A[19][1] * mat_B[1][15] +
                  mat_A[19][2] * mat_B[2][15] +
                  mat_A[19][3] * mat_B[3][15] +
                  mat_A[19][4] * mat_B[4][15] +
                  mat_A[19][5] * mat_B[5][15] +
                  mat_A[19][6] * mat_B[6][15] +
                  mat_A[19][7] * mat_B[7][15] +
                  mat_A[19][8] * mat_B[8][15] +
                  mat_A[19][9] * mat_B[9][15] +
                  mat_A[19][10] * mat_B[10][15] +
                  mat_A[19][11] * mat_B[11][15] +
                  mat_A[19][12] * mat_B[12][15] +
                  mat_A[19][13] * mat_B[13][15] +
                  mat_A[19][14] * mat_B[14][15] +
                  mat_A[19][15] * mat_B[15][15] +
                  mat_A[19][16] * mat_B[16][15] +
                  mat_A[19][17] * mat_B[17][15] +
                  mat_A[19][18] * mat_B[18][15] +
                  mat_A[19][19] * mat_B[19][15] +
                  mat_A[19][20] * mat_B[20][15] +
                  mat_A[19][21] * mat_B[21][15] +
                  mat_A[19][22] * mat_B[22][15] +
                  mat_A[19][23] * mat_B[23][15] +
                  mat_A[19][24] * mat_B[24][15] +
                  mat_A[19][25] * mat_B[25][15] +
                  mat_A[19][26] * mat_B[26][15] +
                  mat_A[19][27] * mat_B[27][15] +
                  mat_A[19][28] * mat_B[28][15] +
                  mat_A[19][29] * mat_B[29][15] +
                  mat_A[19][30] * mat_B[30][15] +
                  mat_A[19][31] * mat_B[31][15];
    mat_C[19][16] <= 
                  mat_A[19][0] * mat_B[0][16] +
                  mat_A[19][1] * mat_B[1][16] +
                  mat_A[19][2] * mat_B[2][16] +
                  mat_A[19][3] * mat_B[3][16] +
                  mat_A[19][4] * mat_B[4][16] +
                  mat_A[19][5] * mat_B[5][16] +
                  mat_A[19][6] * mat_B[6][16] +
                  mat_A[19][7] * mat_B[7][16] +
                  mat_A[19][8] * mat_B[8][16] +
                  mat_A[19][9] * mat_B[9][16] +
                  mat_A[19][10] * mat_B[10][16] +
                  mat_A[19][11] * mat_B[11][16] +
                  mat_A[19][12] * mat_B[12][16] +
                  mat_A[19][13] * mat_B[13][16] +
                  mat_A[19][14] * mat_B[14][16] +
                  mat_A[19][15] * mat_B[15][16] +
                  mat_A[19][16] * mat_B[16][16] +
                  mat_A[19][17] * mat_B[17][16] +
                  mat_A[19][18] * mat_B[18][16] +
                  mat_A[19][19] * mat_B[19][16] +
                  mat_A[19][20] * mat_B[20][16] +
                  mat_A[19][21] * mat_B[21][16] +
                  mat_A[19][22] * mat_B[22][16] +
                  mat_A[19][23] * mat_B[23][16] +
                  mat_A[19][24] * mat_B[24][16] +
                  mat_A[19][25] * mat_B[25][16] +
                  mat_A[19][26] * mat_B[26][16] +
                  mat_A[19][27] * mat_B[27][16] +
                  mat_A[19][28] * mat_B[28][16] +
                  mat_A[19][29] * mat_B[29][16] +
                  mat_A[19][30] * mat_B[30][16] +
                  mat_A[19][31] * mat_B[31][16];
    mat_C[19][17] <= 
                  mat_A[19][0] * mat_B[0][17] +
                  mat_A[19][1] * mat_B[1][17] +
                  mat_A[19][2] * mat_B[2][17] +
                  mat_A[19][3] * mat_B[3][17] +
                  mat_A[19][4] * mat_B[4][17] +
                  mat_A[19][5] * mat_B[5][17] +
                  mat_A[19][6] * mat_B[6][17] +
                  mat_A[19][7] * mat_B[7][17] +
                  mat_A[19][8] * mat_B[8][17] +
                  mat_A[19][9] * mat_B[9][17] +
                  mat_A[19][10] * mat_B[10][17] +
                  mat_A[19][11] * mat_B[11][17] +
                  mat_A[19][12] * mat_B[12][17] +
                  mat_A[19][13] * mat_B[13][17] +
                  mat_A[19][14] * mat_B[14][17] +
                  mat_A[19][15] * mat_B[15][17] +
                  mat_A[19][16] * mat_B[16][17] +
                  mat_A[19][17] * mat_B[17][17] +
                  mat_A[19][18] * mat_B[18][17] +
                  mat_A[19][19] * mat_B[19][17] +
                  mat_A[19][20] * mat_B[20][17] +
                  mat_A[19][21] * mat_B[21][17] +
                  mat_A[19][22] * mat_B[22][17] +
                  mat_A[19][23] * mat_B[23][17] +
                  mat_A[19][24] * mat_B[24][17] +
                  mat_A[19][25] * mat_B[25][17] +
                  mat_A[19][26] * mat_B[26][17] +
                  mat_A[19][27] * mat_B[27][17] +
                  mat_A[19][28] * mat_B[28][17] +
                  mat_A[19][29] * mat_B[29][17] +
                  mat_A[19][30] * mat_B[30][17] +
                  mat_A[19][31] * mat_B[31][17];
    mat_C[19][18] <= 
                  mat_A[19][0] * mat_B[0][18] +
                  mat_A[19][1] * mat_B[1][18] +
                  mat_A[19][2] * mat_B[2][18] +
                  mat_A[19][3] * mat_B[3][18] +
                  mat_A[19][4] * mat_B[4][18] +
                  mat_A[19][5] * mat_B[5][18] +
                  mat_A[19][6] * mat_B[6][18] +
                  mat_A[19][7] * mat_B[7][18] +
                  mat_A[19][8] * mat_B[8][18] +
                  mat_A[19][9] * mat_B[9][18] +
                  mat_A[19][10] * mat_B[10][18] +
                  mat_A[19][11] * mat_B[11][18] +
                  mat_A[19][12] * mat_B[12][18] +
                  mat_A[19][13] * mat_B[13][18] +
                  mat_A[19][14] * mat_B[14][18] +
                  mat_A[19][15] * mat_B[15][18] +
                  mat_A[19][16] * mat_B[16][18] +
                  mat_A[19][17] * mat_B[17][18] +
                  mat_A[19][18] * mat_B[18][18] +
                  mat_A[19][19] * mat_B[19][18] +
                  mat_A[19][20] * mat_B[20][18] +
                  mat_A[19][21] * mat_B[21][18] +
                  mat_A[19][22] * mat_B[22][18] +
                  mat_A[19][23] * mat_B[23][18] +
                  mat_A[19][24] * mat_B[24][18] +
                  mat_A[19][25] * mat_B[25][18] +
                  mat_A[19][26] * mat_B[26][18] +
                  mat_A[19][27] * mat_B[27][18] +
                  mat_A[19][28] * mat_B[28][18] +
                  mat_A[19][29] * mat_B[29][18] +
                  mat_A[19][30] * mat_B[30][18] +
                  mat_A[19][31] * mat_B[31][18];
    mat_C[19][19] <= 
                  mat_A[19][0] * mat_B[0][19] +
                  mat_A[19][1] * mat_B[1][19] +
                  mat_A[19][2] * mat_B[2][19] +
                  mat_A[19][3] * mat_B[3][19] +
                  mat_A[19][4] * mat_B[4][19] +
                  mat_A[19][5] * mat_B[5][19] +
                  mat_A[19][6] * mat_B[6][19] +
                  mat_A[19][7] * mat_B[7][19] +
                  mat_A[19][8] * mat_B[8][19] +
                  mat_A[19][9] * mat_B[9][19] +
                  mat_A[19][10] * mat_B[10][19] +
                  mat_A[19][11] * mat_B[11][19] +
                  mat_A[19][12] * mat_B[12][19] +
                  mat_A[19][13] * mat_B[13][19] +
                  mat_A[19][14] * mat_B[14][19] +
                  mat_A[19][15] * mat_B[15][19] +
                  mat_A[19][16] * mat_B[16][19] +
                  mat_A[19][17] * mat_B[17][19] +
                  mat_A[19][18] * mat_B[18][19] +
                  mat_A[19][19] * mat_B[19][19] +
                  mat_A[19][20] * mat_B[20][19] +
                  mat_A[19][21] * mat_B[21][19] +
                  mat_A[19][22] * mat_B[22][19] +
                  mat_A[19][23] * mat_B[23][19] +
                  mat_A[19][24] * mat_B[24][19] +
                  mat_A[19][25] * mat_B[25][19] +
                  mat_A[19][26] * mat_B[26][19] +
                  mat_A[19][27] * mat_B[27][19] +
                  mat_A[19][28] * mat_B[28][19] +
                  mat_A[19][29] * mat_B[29][19] +
                  mat_A[19][30] * mat_B[30][19] +
                  mat_A[19][31] * mat_B[31][19];
    mat_C[19][20] <= 
                  mat_A[19][0] * mat_B[0][20] +
                  mat_A[19][1] * mat_B[1][20] +
                  mat_A[19][2] * mat_B[2][20] +
                  mat_A[19][3] * mat_B[3][20] +
                  mat_A[19][4] * mat_B[4][20] +
                  mat_A[19][5] * mat_B[5][20] +
                  mat_A[19][6] * mat_B[6][20] +
                  mat_A[19][7] * mat_B[7][20] +
                  mat_A[19][8] * mat_B[8][20] +
                  mat_A[19][9] * mat_B[9][20] +
                  mat_A[19][10] * mat_B[10][20] +
                  mat_A[19][11] * mat_B[11][20] +
                  mat_A[19][12] * mat_B[12][20] +
                  mat_A[19][13] * mat_B[13][20] +
                  mat_A[19][14] * mat_B[14][20] +
                  mat_A[19][15] * mat_B[15][20] +
                  mat_A[19][16] * mat_B[16][20] +
                  mat_A[19][17] * mat_B[17][20] +
                  mat_A[19][18] * mat_B[18][20] +
                  mat_A[19][19] * mat_B[19][20] +
                  mat_A[19][20] * mat_B[20][20] +
                  mat_A[19][21] * mat_B[21][20] +
                  mat_A[19][22] * mat_B[22][20] +
                  mat_A[19][23] * mat_B[23][20] +
                  mat_A[19][24] * mat_B[24][20] +
                  mat_A[19][25] * mat_B[25][20] +
                  mat_A[19][26] * mat_B[26][20] +
                  mat_A[19][27] * mat_B[27][20] +
                  mat_A[19][28] * mat_B[28][20] +
                  mat_A[19][29] * mat_B[29][20] +
                  mat_A[19][30] * mat_B[30][20] +
                  mat_A[19][31] * mat_B[31][20];
    mat_C[19][21] <= 
                  mat_A[19][0] * mat_B[0][21] +
                  mat_A[19][1] * mat_B[1][21] +
                  mat_A[19][2] * mat_B[2][21] +
                  mat_A[19][3] * mat_B[3][21] +
                  mat_A[19][4] * mat_B[4][21] +
                  mat_A[19][5] * mat_B[5][21] +
                  mat_A[19][6] * mat_B[6][21] +
                  mat_A[19][7] * mat_B[7][21] +
                  mat_A[19][8] * mat_B[8][21] +
                  mat_A[19][9] * mat_B[9][21] +
                  mat_A[19][10] * mat_B[10][21] +
                  mat_A[19][11] * mat_B[11][21] +
                  mat_A[19][12] * mat_B[12][21] +
                  mat_A[19][13] * mat_B[13][21] +
                  mat_A[19][14] * mat_B[14][21] +
                  mat_A[19][15] * mat_B[15][21] +
                  mat_A[19][16] * mat_B[16][21] +
                  mat_A[19][17] * mat_B[17][21] +
                  mat_A[19][18] * mat_B[18][21] +
                  mat_A[19][19] * mat_B[19][21] +
                  mat_A[19][20] * mat_B[20][21] +
                  mat_A[19][21] * mat_B[21][21] +
                  mat_A[19][22] * mat_B[22][21] +
                  mat_A[19][23] * mat_B[23][21] +
                  mat_A[19][24] * mat_B[24][21] +
                  mat_A[19][25] * mat_B[25][21] +
                  mat_A[19][26] * mat_B[26][21] +
                  mat_A[19][27] * mat_B[27][21] +
                  mat_A[19][28] * mat_B[28][21] +
                  mat_A[19][29] * mat_B[29][21] +
                  mat_A[19][30] * mat_B[30][21] +
                  mat_A[19][31] * mat_B[31][21];
    mat_C[19][22] <= 
                  mat_A[19][0] * mat_B[0][22] +
                  mat_A[19][1] * mat_B[1][22] +
                  mat_A[19][2] * mat_B[2][22] +
                  mat_A[19][3] * mat_B[3][22] +
                  mat_A[19][4] * mat_B[4][22] +
                  mat_A[19][5] * mat_B[5][22] +
                  mat_A[19][6] * mat_B[6][22] +
                  mat_A[19][7] * mat_B[7][22] +
                  mat_A[19][8] * mat_B[8][22] +
                  mat_A[19][9] * mat_B[9][22] +
                  mat_A[19][10] * mat_B[10][22] +
                  mat_A[19][11] * mat_B[11][22] +
                  mat_A[19][12] * mat_B[12][22] +
                  mat_A[19][13] * mat_B[13][22] +
                  mat_A[19][14] * mat_B[14][22] +
                  mat_A[19][15] * mat_B[15][22] +
                  mat_A[19][16] * mat_B[16][22] +
                  mat_A[19][17] * mat_B[17][22] +
                  mat_A[19][18] * mat_B[18][22] +
                  mat_A[19][19] * mat_B[19][22] +
                  mat_A[19][20] * mat_B[20][22] +
                  mat_A[19][21] * mat_B[21][22] +
                  mat_A[19][22] * mat_B[22][22] +
                  mat_A[19][23] * mat_B[23][22] +
                  mat_A[19][24] * mat_B[24][22] +
                  mat_A[19][25] * mat_B[25][22] +
                  mat_A[19][26] * mat_B[26][22] +
                  mat_A[19][27] * mat_B[27][22] +
                  mat_A[19][28] * mat_B[28][22] +
                  mat_A[19][29] * mat_B[29][22] +
                  mat_A[19][30] * mat_B[30][22] +
                  mat_A[19][31] * mat_B[31][22];
    mat_C[19][23] <= 
                  mat_A[19][0] * mat_B[0][23] +
                  mat_A[19][1] * mat_B[1][23] +
                  mat_A[19][2] * mat_B[2][23] +
                  mat_A[19][3] * mat_B[3][23] +
                  mat_A[19][4] * mat_B[4][23] +
                  mat_A[19][5] * mat_B[5][23] +
                  mat_A[19][6] * mat_B[6][23] +
                  mat_A[19][7] * mat_B[7][23] +
                  mat_A[19][8] * mat_B[8][23] +
                  mat_A[19][9] * mat_B[9][23] +
                  mat_A[19][10] * mat_B[10][23] +
                  mat_A[19][11] * mat_B[11][23] +
                  mat_A[19][12] * mat_B[12][23] +
                  mat_A[19][13] * mat_B[13][23] +
                  mat_A[19][14] * mat_B[14][23] +
                  mat_A[19][15] * mat_B[15][23] +
                  mat_A[19][16] * mat_B[16][23] +
                  mat_A[19][17] * mat_B[17][23] +
                  mat_A[19][18] * mat_B[18][23] +
                  mat_A[19][19] * mat_B[19][23] +
                  mat_A[19][20] * mat_B[20][23] +
                  mat_A[19][21] * mat_B[21][23] +
                  mat_A[19][22] * mat_B[22][23] +
                  mat_A[19][23] * mat_B[23][23] +
                  mat_A[19][24] * mat_B[24][23] +
                  mat_A[19][25] * mat_B[25][23] +
                  mat_A[19][26] * mat_B[26][23] +
                  mat_A[19][27] * mat_B[27][23] +
                  mat_A[19][28] * mat_B[28][23] +
                  mat_A[19][29] * mat_B[29][23] +
                  mat_A[19][30] * mat_B[30][23] +
                  mat_A[19][31] * mat_B[31][23];
    mat_C[19][24] <= 
                  mat_A[19][0] * mat_B[0][24] +
                  mat_A[19][1] * mat_B[1][24] +
                  mat_A[19][2] * mat_B[2][24] +
                  mat_A[19][3] * mat_B[3][24] +
                  mat_A[19][4] * mat_B[4][24] +
                  mat_A[19][5] * mat_B[5][24] +
                  mat_A[19][6] * mat_B[6][24] +
                  mat_A[19][7] * mat_B[7][24] +
                  mat_A[19][8] * mat_B[8][24] +
                  mat_A[19][9] * mat_B[9][24] +
                  mat_A[19][10] * mat_B[10][24] +
                  mat_A[19][11] * mat_B[11][24] +
                  mat_A[19][12] * mat_B[12][24] +
                  mat_A[19][13] * mat_B[13][24] +
                  mat_A[19][14] * mat_B[14][24] +
                  mat_A[19][15] * mat_B[15][24] +
                  mat_A[19][16] * mat_B[16][24] +
                  mat_A[19][17] * mat_B[17][24] +
                  mat_A[19][18] * mat_B[18][24] +
                  mat_A[19][19] * mat_B[19][24] +
                  mat_A[19][20] * mat_B[20][24] +
                  mat_A[19][21] * mat_B[21][24] +
                  mat_A[19][22] * mat_B[22][24] +
                  mat_A[19][23] * mat_B[23][24] +
                  mat_A[19][24] * mat_B[24][24] +
                  mat_A[19][25] * mat_B[25][24] +
                  mat_A[19][26] * mat_B[26][24] +
                  mat_A[19][27] * mat_B[27][24] +
                  mat_A[19][28] * mat_B[28][24] +
                  mat_A[19][29] * mat_B[29][24] +
                  mat_A[19][30] * mat_B[30][24] +
                  mat_A[19][31] * mat_B[31][24];
    mat_C[19][25] <= 
                  mat_A[19][0] * mat_B[0][25] +
                  mat_A[19][1] * mat_B[1][25] +
                  mat_A[19][2] * mat_B[2][25] +
                  mat_A[19][3] * mat_B[3][25] +
                  mat_A[19][4] * mat_B[4][25] +
                  mat_A[19][5] * mat_B[5][25] +
                  mat_A[19][6] * mat_B[6][25] +
                  mat_A[19][7] * mat_B[7][25] +
                  mat_A[19][8] * mat_B[8][25] +
                  mat_A[19][9] * mat_B[9][25] +
                  mat_A[19][10] * mat_B[10][25] +
                  mat_A[19][11] * mat_B[11][25] +
                  mat_A[19][12] * mat_B[12][25] +
                  mat_A[19][13] * mat_B[13][25] +
                  mat_A[19][14] * mat_B[14][25] +
                  mat_A[19][15] * mat_B[15][25] +
                  mat_A[19][16] * mat_B[16][25] +
                  mat_A[19][17] * mat_B[17][25] +
                  mat_A[19][18] * mat_B[18][25] +
                  mat_A[19][19] * mat_B[19][25] +
                  mat_A[19][20] * mat_B[20][25] +
                  mat_A[19][21] * mat_B[21][25] +
                  mat_A[19][22] * mat_B[22][25] +
                  mat_A[19][23] * mat_B[23][25] +
                  mat_A[19][24] * mat_B[24][25] +
                  mat_A[19][25] * mat_B[25][25] +
                  mat_A[19][26] * mat_B[26][25] +
                  mat_A[19][27] * mat_B[27][25] +
                  mat_A[19][28] * mat_B[28][25] +
                  mat_A[19][29] * mat_B[29][25] +
                  mat_A[19][30] * mat_B[30][25] +
                  mat_A[19][31] * mat_B[31][25];
    mat_C[19][26] <= 
                  mat_A[19][0] * mat_B[0][26] +
                  mat_A[19][1] * mat_B[1][26] +
                  mat_A[19][2] * mat_B[2][26] +
                  mat_A[19][3] * mat_B[3][26] +
                  mat_A[19][4] * mat_B[4][26] +
                  mat_A[19][5] * mat_B[5][26] +
                  mat_A[19][6] * mat_B[6][26] +
                  mat_A[19][7] * mat_B[7][26] +
                  mat_A[19][8] * mat_B[8][26] +
                  mat_A[19][9] * mat_B[9][26] +
                  mat_A[19][10] * mat_B[10][26] +
                  mat_A[19][11] * mat_B[11][26] +
                  mat_A[19][12] * mat_B[12][26] +
                  mat_A[19][13] * mat_B[13][26] +
                  mat_A[19][14] * mat_B[14][26] +
                  mat_A[19][15] * mat_B[15][26] +
                  mat_A[19][16] * mat_B[16][26] +
                  mat_A[19][17] * mat_B[17][26] +
                  mat_A[19][18] * mat_B[18][26] +
                  mat_A[19][19] * mat_B[19][26] +
                  mat_A[19][20] * mat_B[20][26] +
                  mat_A[19][21] * mat_B[21][26] +
                  mat_A[19][22] * mat_B[22][26] +
                  mat_A[19][23] * mat_B[23][26] +
                  mat_A[19][24] * mat_B[24][26] +
                  mat_A[19][25] * mat_B[25][26] +
                  mat_A[19][26] * mat_B[26][26] +
                  mat_A[19][27] * mat_B[27][26] +
                  mat_A[19][28] * mat_B[28][26] +
                  mat_A[19][29] * mat_B[29][26] +
                  mat_A[19][30] * mat_B[30][26] +
                  mat_A[19][31] * mat_B[31][26];
    mat_C[19][27] <= 
                  mat_A[19][0] * mat_B[0][27] +
                  mat_A[19][1] * mat_B[1][27] +
                  mat_A[19][2] * mat_B[2][27] +
                  mat_A[19][3] * mat_B[3][27] +
                  mat_A[19][4] * mat_B[4][27] +
                  mat_A[19][5] * mat_B[5][27] +
                  mat_A[19][6] * mat_B[6][27] +
                  mat_A[19][7] * mat_B[7][27] +
                  mat_A[19][8] * mat_B[8][27] +
                  mat_A[19][9] * mat_B[9][27] +
                  mat_A[19][10] * mat_B[10][27] +
                  mat_A[19][11] * mat_B[11][27] +
                  mat_A[19][12] * mat_B[12][27] +
                  mat_A[19][13] * mat_B[13][27] +
                  mat_A[19][14] * mat_B[14][27] +
                  mat_A[19][15] * mat_B[15][27] +
                  mat_A[19][16] * mat_B[16][27] +
                  mat_A[19][17] * mat_B[17][27] +
                  mat_A[19][18] * mat_B[18][27] +
                  mat_A[19][19] * mat_B[19][27] +
                  mat_A[19][20] * mat_B[20][27] +
                  mat_A[19][21] * mat_B[21][27] +
                  mat_A[19][22] * mat_B[22][27] +
                  mat_A[19][23] * mat_B[23][27] +
                  mat_A[19][24] * mat_B[24][27] +
                  mat_A[19][25] * mat_B[25][27] +
                  mat_A[19][26] * mat_B[26][27] +
                  mat_A[19][27] * mat_B[27][27] +
                  mat_A[19][28] * mat_B[28][27] +
                  mat_A[19][29] * mat_B[29][27] +
                  mat_A[19][30] * mat_B[30][27] +
                  mat_A[19][31] * mat_B[31][27];
    mat_C[19][28] <= 
                  mat_A[19][0] * mat_B[0][28] +
                  mat_A[19][1] * mat_B[1][28] +
                  mat_A[19][2] * mat_B[2][28] +
                  mat_A[19][3] * mat_B[3][28] +
                  mat_A[19][4] * mat_B[4][28] +
                  mat_A[19][5] * mat_B[5][28] +
                  mat_A[19][6] * mat_B[6][28] +
                  mat_A[19][7] * mat_B[7][28] +
                  mat_A[19][8] * mat_B[8][28] +
                  mat_A[19][9] * mat_B[9][28] +
                  mat_A[19][10] * mat_B[10][28] +
                  mat_A[19][11] * mat_B[11][28] +
                  mat_A[19][12] * mat_B[12][28] +
                  mat_A[19][13] * mat_B[13][28] +
                  mat_A[19][14] * mat_B[14][28] +
                  mat_A[19][15] * mat_B[15][28] +
                  mat_A[19][16] * mat_B[16][28] +
                  mat_A[19][17] * mat_B[17][28] +
                  mat_A[19][18] * mat_B[18][28] +
                  mat_A[19][19] * mat_B[19][28] +
                  mat_A[19][20] * mat_B[20][28] +
                  mat_A[19][21] * mat_B[21][28] +
                  mat_A[19][22] * mat_B[22][28] +
                  mat_A[19][23] * mat_B[23][28] +
                  mat_A[19][24] * mat_B[24][28] +
                  mat_A[19][25] * mat_B[25][28] +
                  mat_A[19][26] * mat_B[26][28] +
                  mat_A[19][27] * mat_B[27][28] +
                  mat_A[19][28] * mat_B[28][28] +
                  mat_A[19][29] * mat_B[29][28] +
                  mat_A[19][30] * mat_B[30][28] +
                  mat_A[19][31] * mat_B[31][28];
    mat_C[19][29] <= 
                  mat_A[19][0] * mat_B[0][29] +
                  mat_A[19][1] * mat_B[1][29] +
                  mat_A[19][2] * mat_B[2][29] +
                  mat_A[19][3] * mat_B[3][29] +
                  mat_A[19][4] * mat_B[4][29] +
                  mat_A[19][5] * mat_B[5][29] +
                  mat_A[19][6] * mat_B[6][29] +
                  mat_A[19][7] * mat_B[7][29] +
                  mat_A[19][8] * mat_B[8][29] +
                  mat_A[19][9] * mat_B[9][29] +
                  mat_A[19][10] * mat_B[10][29] +
                  mat_A[19][11] * mat_B[11][29] +
                  mat_A[19][12] * mat_B[12][29] +
                  mat_A[19][13] * mat_B[13][29] +
                  mat_A[19][14] * mat_B[14][29] +
                  mat_A[19][15] * mat_B[15][29] +
                  mat_A[19][16] * mat_B[16][29] +
                  mat_A[19][17] * mat_B[17][29] +
                  mat_A[19][18] * mat_B[18][29] +
                  mat_A[19][19] * mat_B[19][29] +
                  mat_A[19][20] * mat_B[20][29] +
                  mat_A[19][21] * mat_B[21][29] +
                  mat_A[19][22] * mat_B[22][29] +
                  mat_A[19][23] * mat_B[23][29] +
                  mat_A[19][24] * mat_B[24][29] +
                  mat_A[19][25] * mat_B[25][29] +
                  mat_A[19][26] * mat_B[26][29] +
                  mat_A[19][27] * mat_B[27][29] +
                  mat_A[19][28] * mat_B[28][29] +
                  mat_A[19][29] * mat_B[29][29] +
                  mat_A[19][30] * mat_B[30][29] +
                  mat_A[19][31] * mat_B[31][29];
    mat_C[19][30] <= 
                  mat_A[19][0] * mat_B[0][30] +
                  mat_A[19][1] * mat_B[1][30] +
                  mat_A[19][2] * mat_B[2][30] +
                  mat_A[19][3] * mat_B[3][30] +
                  mat_A[19][4] * mat_B[4][30] +
                  mat_A[19][5] * mat_B[5][30] +
                  mat_A[19][6] * mat_B[6][30] +
                  mat_A[19][7] * mat_B[7][30] +
                  mat_A[19][8] * mat_B[8][30] +
                  mat_A[19][9] * mat_B[9][30] +
                  mat_A[19][10] * mat_B[10][30] +
                  mat_A[19][11] * mat_B[11][30] +
                  mat_A[19][12] * mat_B[12][30] +
                  mat_A[19][13] * mat_B[13][30] +
                  mat_A[19][14] * mat_B[14][30] +
                  mat_A[19][15] * mat_B[15][30] +
                  mat_A[19][16] * mat_B[16][30] +
                  mat_A[19][17] * mat_B[17][30] +
                  mat_A[19][18] * mat_B[18][30] +
                  mat_A[19][19] * mat_B[19][30] +
                  mat_A[19][20] * mat_B[20][30] +
                  mat_A[19][21] * mat_B[21][30] +
                  mat_A[19][22] * mat_B[22][30] +
                  mat_A[19][23] * mat_B[23][30] +
                  mat_A[19][24] * mat_B[24][30] +
                  mat_A[19][25] * mat_B[25][30] +
                  mat_A[19][26] * mat_B[26][30] +
                  mat_A[19][27] * mat_B[27][30] +
                  mat_A[19][28] * mat_B[28][30] +
                  mat_A[19][29] * mat_B[29][30] +
                  mat_A[19][30] * mat_B[30][30] +
                  mat_A[19][31] * mat_B[31][30];
    mat_C[19][31] <= 
                  mat_A[19][0] * mat_B[0][31] +
                  mat_A[19][1] * mat_B[1][31] +
                  mat_A[19][2] * mat_B[2][31] +
                  mat_A[19][3] * mat_B[3][31] +
                  mat_A[19][4] * mat_B[4][31] +
                  mat_A[19][5] * mat_B[5][31] +
                  mat_A[19][6] * mat_B[6][31] +
                  mat_A[19][7] * mat_B[7][31] +
                  mat_A[19][8] * mat_B[8][31] +
                  mat_A[19][9] * mat_B[9][31] +
                  mat_A[19][10] * mat_B[10][31] +
                  mat_A[19][11] * mat_B[11][31] +
                  mat_A[19][12] * mat_B[12][31] +
                  mat_A[19][13] * mat_B[13][31] +
                  mat_A[19][14] * mat_B[14][31] +
                  mat_A[19][15] * mat_B[15][31] +
                  mat_A[19][16] * mat_B[16][31] +
                  mat_A[19][17] * mat_B[17][31] +
                  mat_A[19][18] * mat_B[18][31] +
                  mat_A[19][19] * mat_B[19][31] +
                  mat_A[19][20] * mat_B[20][31] +
                  mat_A[19][21] * mat_B[21][31] +
                  mat_A[19][22] * mat_B[22][31] +
                  mat_A[19][23] * mat_B[23][31] +
                  mat_A[19][24] * mat_B[24][31] +
                  mat_A[19][25] * mat_B[25][31] +
                  mat_A[19][26] * mat_B[26][31] +
                  mat_A[19][27] * mat_B[27][31] +
                  mat_A[19][28] * mat_B[28][31] +
                  mat_A[19][29] * mat_B[29][31] +
                  mat_A[19][30] * mat_B[30][31] +
                  mat_A[19][31] * mat_B[31][31];
    mat_C[20][0] <= 
                  mat_A[20][0] * mat_B[0][0] +
                  mat_A[20][1] * mat_B[1][0] +
                  mat_A[20][2] * mat_B[2][0] +
                  mat_A[20][3] * mat_B[3][0] +
                  mat_A[20][4] * mat_B[4][0] +
                  mat_A[20][5] * mat_B[5][0] +
                  mat_A[20][6] * mat_B[6][0] +
                  mat_A[20][7] * mat_B[7][0] +
                  mat_A[20][8] * mat_B[8][0] +
                  mat_A[20][9] * mat_B[9][0] +
                  mat_A[20][10] * mat_B[10][0] +
                  mat_A[20][11] * mat_B[11][0] +
                  mat_A[20][12] * mat_B[12][0] +
                  mat_A[20][13] * mat_B[13][0] +
                  mat_A[20][14] * mat_B[14][0] +
                  mat_A[20][15] * mat_B[15][0] +
                  mat_A[20][16] * mat_B[16][0] +
                  mat_A[20][17] * mat_B[17][0] +
                  mat_A[20][18] * mat_B[18][0] +
                  mat_A[20][19] * mat_B[19][0] +
                  mat_A[20][20] * mat_B[20][0] +
                  mat_A[20][21] * mat_B[21][0] +
                  mat_A[20][22] * mat_B[22][0] +
                  mat_A[20][23] * mat_B[23][0] +
                  mat_A[20][24] * mat_B[24][0] +
                  mat_A[20][25] * mat_B[25][0] +
                  mat_A[20][26] * mat_B[26][0] +
                  mat_A[20][27] * mat_B[27][0] +
                  mat_A[20][28] * mat_B[28][0] +
                  mat_A[20][29] * mat_B[29][0] +
                  mat_A[20][30] * mat_B[30][0] +
                  mat_A[20][31] * mat_B[31][0];
    mat_C[20][1] <= 
                  mat_A[20][0] * mat_B[0][1] +
                  mat_A[20][1] * mat_B[1][1] +
                  mat_A[20][2] * mat_B[2][1] +
                  mat_A[20][3] * mat_B[3][1] +
                  mat_A[20][4] * mat_B[4][1] +
                  mat_A[20][5] * mat_B[5][1] +
                  mat_A[20][6] * mat_B[6][1] +
                  mat_A[20][7] * mat_B[7][1] +
                  mat_A[20][8] * mat_B[8][1] +
                  mat_A[20][9] * mat_B[9][1] +
                  mat_A[20][10] * mat_B[10][1] +
                  mat_A[20][11] * mat_B[11][1] +
                  mat_A[20][12] * mat_B[12][1] +
                  mat_A[20][13] * mat_B[13][1] +
                  mat_A[20][14] * mat_B[14][1] +
                  mat_A[20][15] * mat_B[15][1] +
                  mat_A[20][16] * mat_B[16][1] +
                  mat_A[20][17] * mat_B[17][1] +
                  mat_A[20][18] * mat_B[18][1] +
                  mat_A[20][19] * mat_B[19][1] +
                  mat_A[20][20] * mat_B[20][1] +
                  mat_A[20][21] * mat_B[21][1] +
                  mat_A[20][22] * mat_B[22][1] +
                  mat_A[20][23] * mat_B[23][1] +
                  mat_A[20][24] * mat_B[24][1] +
                  mat_A[20][25] * mat_B[25][1] +
                  mat_A[20][26] * mat_B[26][1] +
                  mat_A[20][27] * mat_B[27][1] +
                  mat_A[20][28] * mat_B[28][1] +
                  mat_A[20][29] * mat_B[29][1] +
                  mat_A[20][30] * mat_B[30][1] +
                  mat_A[20][31] * mat_B[31][1];
    mat_C[20][2] <= 
                  mat_A[20][0] * mat_B[0][2] +
                  mat_A[20][1] * mat_B[1][2] +
                  mat_A[20][2] * mat_B[2][2] +
                  mat_A[20][3] * mat_B[3][2] +
                  mat_A[20][4] * mat_B[4][2] +
                  mat_A[20][5] * mat_B[5][2] +
                  mat_A[20][6] * mat_B[6][2] +
                  mat_A[20][7] * mat_B[7][2] +
                  mat_A[20][8] * mat_B[8][2] +
                  mat_A[20][9] * mat_B[9][2] +
                  mat_A[20][10] * mat_B[10][2] +
                  mat_A[20][11] * mat_B[11][2] +
                  mat_A[20][12] * mat_B[12][2] +
                  mat_A[20][13] * mat_B[13][2] +
                  mat_A[20][14] * mat_B[14][2] +
                  mat_A[20][15] * mat_B[15][2] +
                  mat_A[20][16] * mat_B[16][2] +
                  mat_A[20][17] * mat_B[17][2] +
                  mat_A[20][18] * mat_B[18][2] +
                  mat_A[20][19] * mat_B[19][2] +
                  mat_A[20][20] * mat_B[20][2] +
                  mat_A[20][21] * mat_B[21][2] +
                  mat_A[20][22] * mat_B[22][2] +
                  mat_A[20][23] * mat_B[23][2] +
                  mat_A[20][24] * mat_B[24][2] +
                  mat_A[20][25] * mat_B[25][2] +
                  mat_A[20][26] * mat_B[26][2] +
                  mat_A[20][27] * mat_B[27][2] +
                  mat_A[20][28] * mat_B[28][2] +
                  mat_A[20][29] * mat_B[29][2] +
                  mat_A[20][30] * mat_B[30][2] +
                  mat_A[20][31] * mat_B[31][2];
    mat_C[20][3] <= 
                  mat_A[20][0] * mat_B[0][3] +
                  mat_A[20][1] * mat_B[1][3] +
                  mat_A[20][2] * mat_B[2][3] +
                  mat_A[20][3] * mat_B[3][3] +
                  mat_A[20][4] * mat_B[4][3] +
                  mat_A[20][5] * mat_B[5][3] +
                  mat_A[20][6] * mat_B[6][3] +
                  mat_A[20][7] * mat_B[7][3] +
                  mat_A[20][8] * mat_B[8][3] +
                  mat_A[20][9] * mat_B[9][3] +
                  mat_A[20][10] * mat_B[10][3] +
                  mat_A[20][11] * mat_B[11][3] +
                  mat_A[20][12] * mat_B[12][3] +
                  mat_A[20][13] * mat_B[13][3] +
                  mat_A[20][14] * mat_B[14][3] +
                  mat_A[20][15] * mat_B[15][3] +
                  mat_A[20][16] * mat_B[16][3] +
                  mat_A[20][17] * mat_B[17][3] +
                  mat_A[20][18] * mat_B[18][3] +
                  mat_A[20][19] * mat_B[19][3] +
                  mat_A[20][20] * mat_B[20][3] +
                  mat_A[20][21] * mat_B[21][3] +
                  mat_A[20][22] * mat_B[22][3] +
                  mat_A[20][23] * mat_B[23][3] +
                  mat_A[20][24] * mat_B[24][3] +
                  mat_A[20][25] * mat_B[25][3] +
                  mat_A[20][26] * mat_B[26][3] +
                  mat_A[20][27] * mat_B[27][3] +
                  mat_A[20][28] * mat_B[28][3] +
                  mat_A[20][29] * mat_B[29][3] +
                  mat_A[20][30] * mat_B[30][3] +
                  mat_A[20][31] * mat_B[31][3];
    mat_C[20][4] <= 
                  mat_A[20][0] * mat_B[0][4] +
                  mat_A[20][1] * mat_B[1][4] +
                  mat_A[20][2] * mat_B[2][4] +
                  mat_A[20][3] * mat_B[3][4] +
                  mat_A[20][4] * mat_B[4][4] +
                  mat_A[20][5] * mat_B[5][4] +
                  mat_A[20][6] * mat_B[6][4] +
                  mat_A[20][7] * mat_B[7][4] +
                  mat_A[20][8] * mat_B[8][4] +
                  mat_A[20][9] * mat_B[9][4] +
                  mat_A[20][10] * mat_B[10][4] +
                  mat_A[20][11] * mat_B[11][4] +
                  mat_A[20][12] * mat_B[12][4] +
                  mat_A[20][13] * mat_B[13][4] +
                  mat_A[20][14] * mat_B[14][4] +
                  mat_A[20][15] * mat_B[15][4] +
                  mat_A[20][16] * mat_B[16][4] +
                  mat_A[20][17] * mat_B[17][4] +
                  mat_A[20][18] * mat_B[18][4] +
                  mat_A[20][19] * mat_B[19][4] +
                  mat_A[20][20] * mat_B[20][4] +
                  mat_A[20][21] * mat_B[21][4] +
                  mat_A[20][22] * mat_B[22][4] +
                  mat_A[20][23] * mat_B[23][4] +
                  mat_A[20][24] * mat_B[24][4] +
                  mat_A[20][25] * mat_B[25][4] +
                  mat_A[20][26] * mat_B[26][4] +
                  mat_A[20][27] * mat_B[27][4] +
                  mat_A[20][28] * mat_B[28][4] +
                  mat_A[20][29] * mat_B[29][4] +
                  mat_A[20][30] * mat_B[30][4] +
                  mat_A[20][31] * mat_B[31][4];
    mat_C[20][5] <= 
                  mat_A[20][0] * mat_B[0][5] +
                  mat_A[20][1] * mat_B[1][5] +
                  mat_A[20][2] * mat_B[2][5] +
                  mat_A[20][3] * mat_B[3][5] +
                  mat_A[20][4] * mat_B[4][5] +
                  mat_A[20][5] * mat_B[5][5] +
                  mat_A[20][6] * mat_B[6][5] +
                  mat_A[20][7] * mat_B[7][5] +
                  mat_A[20][8] * mat_B[8][5] +
                  mat_A[20][9] * mat_B[9][5] +
                  mat_A[20][10] * mat_B[10][5] +
                  mat_A[20][11] * mat_B[11][5] +
                  mat_A[20][12] * mat_B[12][5] +
                  mat_A[20][13] * mat_B[13][5] +
                  mat_A[20][14] * mat_B[14][5] +
                  mat_A[20][15] * mat_B[15][5] +
                  mat_A[20][16] * mat_B[16][5] +
                  mat_A[20][17] * mat_B[17][5] +
                  mat_A[20][18] * mat_B[18][5] +
                  mat_A[20][19] * mat_B[19][5] +
                  mat_A[20][20] * mat_B[20][5] +
                  mat_A[20][21] * mat_B[21][5] +
                  mat_A[20][22] * mat_B[22][5] +
                  mat_A[20][23] * mat_B[23][5] +
                  mat_A[20][24] * mat_B[24][5] +
                  mat_A[20][25] * mat_B[25][5] +
                  mat_A[20][26] * mat_B[26][5] +
                  mat_A[20][27] * mat_B[27][5] +
                  mat_A[20][28] * mat_B[28][5] +
                  mat_A[20][29] * mat_B[29][5] +
                  mat_A[20][30] * mat_B[30][5] +
                  mat_A[20][31] * mat_B[31][5];
    mat_C[20][6] <= 
                  mat_A[20][0] * mat_B[0][6] +
                  mat_A[20][1] * mat_B[1][6] +
                  mat_A[20][2] * mat_B[2][6] +
                  mat_A[20][3] * mat_B[3][6] +
                  mat_A[20][4] * mat_B[4][6] +
                  mat_A[20][5] * mat_B[5][6] +
                  mat_A[20][6] * mat_B[6][6] +
                  mat_A[20][7] * mat_B[7][6] +
                  mat_A[20][8] * mat_B[8][6] +
                  mat_A[20][9] * mat_B[9][6] +
                  mat_A[20][10] * mat_B[10][6] +
                  mat_A[20][11] * mat_B[11][6] +
                  mat_A[20][12] * mat_B[12][6] +
                  mat_A[20][13] * mat_B[13][6] +
                  mat_A[20][14] * mat_B[14][6] +
                  mat_A[20][15] * mat_B[15][6] +
                  mat_A[20][16] * mat_B[16][6] +
                  mat_A[20][17] * mat_B[17][6] +
                  mat_A[20][18] * mat_B[18][6] +
                  mat_A[20][19] * mat_B[19][6] +
                  mat_A[20][20] * mat_B[20][6] +
                  mat_A[20][21] * mat_B[21][6] +
                  mat_A[20][22] * mat_B[22][6] +
                  mat_A[20][23] * mat_B[23][6] +
                  mat_A[20][24] * mat_B[24][6] +
                  mat_A[20][25] * mat_B[25][6] +
                  mat_A[20][26] * mat_B[26][6] +
                  mat_A[20][27] * mat_B[27][6] +
                  mat_A[20][28] * mat_B[28][6] +
                  mat_A[20][29] * mat_B[29][6] +
                  mat_A[20][30] * mat_B[30][6] +
                  mat_A[20][31] * mat_B[31][6];
    mat_C[20][7] <= 
                  mat_A[20][0] * mat_B[0][7] +
                  mat_A[20][1] * mat_B[1][7] +
                  mat_A[20][2] * mat_B[2][7] +
                  mat_A[20][3] * mat_B[3][7] +
                  mat_A[20][4] * mat_B[4][7] +
                  mat_A[20][5] * mat_B[5][7] +
                  mat_A[20][6] * mat_B[6][7] +
                  mat_A[20][7] * mat_B[7][7] +
                  mat_A[20][8] * mat_B[8][7] +
                  mat_A[20][9] * mat_B[9][7] +
                  mat_A[20][10] * mat_B[10][7] +
                  mat_A[20][11] * mat_B[11][7] +
                  mat_A[20][12] * mat_B[12][7] +
                  mat_A[20][13] * mat_B[13][7] +
                  mat_A[20][14] * mat_B[14][7] +
                  mat_A[20][15] * mat_B[15][7] +
                  mat_A[20][16] * mat_B[16][7] +
                  mat_A[20][17] * mat_B[17][7] +
                  mat_A[20][18] * mat_B[18][7] +
                  mat_A[20][19] * mat_B[19][7] +
                  mat_A[20][20] * mat_B[20][7] +
                  mat_A[20][21] * mat_B[21][7] +
                  mat_A[20][22] * mat_B[22][7] +
                  mat_A[20][23] * mat_B[23][7] +
                  mat_A[20][24] * mat_B[24][7] +
                  mat_A[20][25] * mat_B[25][7] +
                  mat_A[20][26] * mat_B[26][7] +
                  mat_A[20][27] * mat_B[27][7] +
                  mat_A[20][28] * mat_B[28][7] +
                  mat_A[20][29] * mat_B[29][7] +
                  mat_A[20][30] * mat_B[30][7] +
                  mat_A[20][31] * mat_B[31][7];
    mat_C[20][8] <= 
                  mat_A[20][0] * mat_B[0][8] +
                  mat_A[20][1] * mat_B[1][8] +
                  mat_A[20][2] * mat_B[2][8] +
                  mat_A[20][3] * mat_B[3][8] +
                  mat_A[20][4] * mat_B[4][8] +
                  mat_A[20][5] * mat_B[5][8] +
                  mat_A[20][6] * mat_B[6][8] +
                  mat_A[20][7] * mat_B[7][8] +
                  mat_A[20][8] * mat_B[8][8] +
                  mat_A[20][9] * mat_B[9][8] +
                  mat_A[20][10] * mat_B[10][8] +
                  mat_A[20][11] * mat_B[11][8] +
                  mat_A[20][12] * mat_B[12][8] +
                  mat_A[20][13] * mat_B[13][8] +
                  mat_A[20][14] * mat_B[14][8] +
                  mat_A[20][15] * mat_B[15][8] +
                  mat_A[20][16] * mat_B[16][8] +
                  mat_A[20][17] * mat_B[17][8] +
                  mat_A[20][18] * mat_B[18][8] +
                  mat_A[20][19] * mat_B[19][8] +
                  mat_A[20][20] * mat_B[20][8] +
                  mat_A[20][21] * mat_B[21][8] +
                  mat_A[20][22] * mat_B[22][8] +
                  mat_A[20][23] * mat_B[23][8] +
                  mat_A[20][24] * mat_B[24][8] +
                  mat_A[20][25] * mat_B[25][8] +
                  mat_A[20][26] * mat_B[26][8] +
                  mat_A[20][27] * mat_B[27][8] +
                  mat_A[20][28] * mat_B[28][8] +
                  mat_A[20][29] * mat_B[29][8] +
                  mat_A[20][30] * mat_B[30][8] +
                  mat_A[20][31] * mat_B[31][8];
    mat_C[20][9] <= 
                  mat_A[20][0] * mat_B[0][9] +
                  mat_A[20][1] * mat_B[1][9] +
                  mat_A[20][2] * mat_B[2][9] +
                  mat_A[20][3] * mat_B[3][9] +
                  mat_A[20][4] * mat_B[4][9] +
                  mat_A[20][5] * mat_B[5][9] +
                  mat_A[20][6] * mat_B[6][9] +
                  mat_A[20][7] * mat_B[7][9] +
                  mat_A[20][8] * mat_B[8][9] +
                  mat_A[20][9] * mat_B[9][9] +
                  mat_A[20][10] * mat_B[10][9] +
                  mat_A[20][11] * mat_B[11][9] +
                  mat_A[20][12] * mat_B[12][9] +
                  mat_A[20][13] * mat_B[13][9] +
                  mat_A[20][14] * mat_B[14][9] +
                  mat_A[20][15] * mat_B[15][9] +
                  mat_A[20][16] * mat_B[16][9] +
                  mat_A[20][17] * mat_B[17][9] +
                  mat_A[20][18] * mat_B[18][9] +
                  mat_A[20][19] * mat_B[19][9] +
                  mat_A[20][20] * mat_B[20][9] +
                  mat_A[20][21] * mat_B[21][9] +
                  mat_A[20][22] * mat_B[22][9] +
                  mat_A[20][23] * mat_B[23][9] +
                  mat_A[20][24] * mat_B[24][9] +
                  mat_A[20][25] * mat_B[25][9] +
                  mat_A[20][26] * mat_B[26][9] +
                  mat_A[20][27] * mat_B[27][9] +
                  mat_A[20][28] * mat_B[28][9] +
                  mat_A[20][29] * mat_B[29][9] +
                  mat_A[20][30] * mat_B[30][9] +
                  mat_A[20][31] * mat_B[31][9];
    mat_C[20][10] <= 
                  mat_A[20][0] * mat_B[0][10] +
                  mat_A[20][1] * mat_B[1][10] +
                  mat_A[20][2] * mat_B[2][10] +
                  mat_A[20][3] * mat_B[3][10] +
                  mat_A[20][4] * mat_B[4][10] +
                  mat_A[20][5] * mat_B[5][10] +
                  mat_A[20][6] * mat_B[6][10] +
                  mat_A[20][7] * mat_B[7][10] +
                  mat_A[20][8] * mat_B[8][10] +
                  mat_A[20][9] * mat_B[9][10] +
                  mat_A[20][10] * mat_B[10][10] +
                  mat_A[20][11] * mat_B[11][10] +
                  mat_A[20][12] * mat_B[12][10] +
                  mat_A[20][13] * mat_B[13][10] +
                  mat_A[20][14] * mat_B[14][10] +
                  mat_A[20][15] * mat_B[15][10] +
                  mat_A[20][16] * mat_B[16][10] +
                  mat_A[20][17] * mat_B[17][10] +
                  mat_A[20][18] * mat_B[18][10] +
                  mat_A[20][19] * mat_B[19][10] +
                  mat_A[20][20] * mat_B[20][10] +
                  mat_A[20][21] * mat_B[21][10] +
                  mat_A[20][22] * mat_B[22][10] +
                  mat_A[20][23] * mat_B[23][10] +
                  mat_A[20][24] * mat_B[24][10] +
                  mat_A[20][25] * mat_B[25][10] +
                  mat_A[20][26] * mat_B[26][10] +
                  mat_A[20][27] * mat_B[27][10] +
                  mat_A[20][28] * mat_B[28][10] +
                  mat_A[20][29] * mat_B[29][10] +
                  mat_A[20][30] * mat_B[30][10] +
                  mat_A[20][31] * mat_B[31][10];
    mat_C[20][11] <= 
                  mat_A[20][0] * mat_B[0][11] +
                  mat_A[20][1] * mat_B[1][11] +
                  mat_A[20][2] * mat_B[2][11] +
                  mat_A[20][3] * mat_B[3][11] +
                  mat_A[20][4] * mat_B[4][11] +
                  mat_A[20][5] * mat_B[5][11] +
                  mat_A[20][6] * mat_B[6][11] +
                  mat_A[20][7] * mat_B[7][11] +
                  mat_A[20][8] * mat_B[8][11] +
                  mat_A[20][9] * mat_B[9][11] +
                  mat_A[20][10] * mat_B[10][11] +
                  mat_A[20][11] * mat_B[11][11] +
                  mat_A[20][12] * mat_B[12][11] +
                  mat_A[20][13] * mat_B[13][11] +
                  mat_A[20][14] * mat_B[14][11] +
                  mat_A[20][15] * mat_B[15][11] +
                  mat_A[20][16] * mat_B[16][11] +
                  mat_A[20][17] * mat_B[17][11] +
                  mat_A[20][18] * mat_B[18][11] +
                  mat_A[20][19] * mat_B[19][11] +
                  mat_A[20][20] * mat_B[20][11] +
                  mat_A[20][21] * mat_B[21][11] +
                  mat_A[20][22] * mat_B[22][11] +
                  mat_A[20][23] * mat_B[23][11] +
                  mat_A[20][24] * mat_B[24][11] +
                  mat_A[20][25] * mat_B[25][11] +
                  mat_A[20][26] * mat_B[26][11] +
                  mat_A[20][27] * mat_B[27][11] +
                  mat_A[20][28] * mat_B[28][11] +
                  mat_A[20][29] * mat_B[29][11] +
                  mat_A[20][30] * mat_B[30][11] +
                  mat_A[20][31] * mat_B[31][11];
    mat_C[20][12] <= 
                  mat_A[20][0] * mat_B[0][12] +
                  mat_A[20][1] * mat_B[1][12] +
                  mat_A[20][2] * mat_B[2][12] +
                  mat_A[20][3] * mat_B[3][12] +
                  mat_A[20][4] * mat_B[4][12] +
                  mat_A[20][5] * mat_B[5][12] +
                  mat_A[20][6] * mat_B[6][12] +
                  mat_A[20][7] * mat_B[7][12] +
                  mat_A[20][8] * mat_B[8][12] +
                  mat_A[20][9] * mat_B[9][12] +
                  mat_A[20][10] * mat_B[10][12] +
                  mat_A[20][11] * mat_B[11][12] +
                  mat_A[20][12] * mat_B[12][12] +
                  mat_A[20][13] * mat_B[13][12] +
                  mat_A[20][14] * mat_B[14][12] +
                  mat_A[20][15] * mat_B[15][12] +
                  mat_A[20][16] * mat_B[16][12] +
                  mat_A[20][17] * mat_B[17][12] +
                  mat_A[20][18] * mat_B[18][12] +
                  mat_A[20][19] * mat_B[19][12] +
                  mat_A[20][20] * mat_B[20][12] +
                  mat_A[20][21] * mat_B[21][12] +
                  mat_A[20][22] * mat_B[22][12] +
                  mat_A[20][23] * mat_B[23][12] +
                  mat_A[20][24] * mat_B[24][12] +
                  mat_A[20][25] * mat_B[25][12] +
                  mat_A[20][26] * mat_B[26][12] +
                  mat_A[20][27] * mat_B[27][12] +
                  mat_A[20][28] * mat_B[28][12] +
                  mat_A[20][29] * mat_B[29][12] +
                  mat_A[20][30] * mat_B[30][12] +
                  mat_A[20][31] * mat_B[31][12];
    mat_C[20][13] <= 
                  mat_A[20][0] * mat_B[0][13] +
                  mat_A[20][1] * mat_B[1][13] +
                  mat_A[20][2] * mat_B[2][13] +
                  mat_A[20][3] * mat_B[3][13] +
                  mat_A[20][4] * mat_B[4][13] +
                  mat_A[20][5] * mat_B[5][13] +
                  mat_A[20][6] * mat_B[6][13] +
                  mat_A[20][7] * mat_B[7][13] +
                  mat_A[20][8] * mat_B[8][13] +
                  mat_A[20][9] * mat_B[9][13] +
                  mat_A[20][10] * mat_B[10][13] +
                  mat_A[20][11] * mat_B[11][13] +
                  mat_A[20][12] * mat_B[12][13] +
                  mat_A[20][13] * mat_B[13][13] +
                  mat_A[20][14] * mat_B[14][13] +
                  mat_A[20][15] * mat_B[15][13] +
                  mat_A[20][16] * mat_B[16][13] +
                  mat_A[20][17] * mat_B[17][13] +
                  mat_A[20][18] * mat_B[18][13] +
                  mat_A[20][19] * mat_B[19][13] +
                  mat_A[20][20] * mat_B[20][13] +
                  mat_A[20][21] * mat_B[21][13] +
                  mat_A[20][22] * mat_B[22][13] +
                  mat_A[20][23] * mat_B[23][13] +
                  mat_A[20][24] * mat_B[24][13] +
                  mat_A[20][25] * mat_B[25][13] +
                  mat_A[20][26] * mat_B[26][13] +
                  mat_A[20][27] * mat_B[27][13] +
                  mat_A[20][28] * mat_B[28][13] +
                  mat_A[20][29] * mat_B[29][13] +
                  mat_A[20][30] * mat_B[30][13] +
                  mat_A[20][31] * mat_B[31][13];
    mat_C[20][14] <= 
                  mat_A[20][0] * mat_B[0][14] +
                  mat_A[20][1] * mat_B[1][14] +
                  mat_A[20][2] * mat_B[2][14] +
                  mat_A[20][3] * mat_B[3][14] +
                  mat_A[20][4] * mat_B[4][14] +
                  mat_A[20][5] * mat_B[5][14] +
                  mat_A[20][6] * mat_B[6][14] +
                  mat_A[20][7] * mat_B[7][14] +
                  mat_A[20][8] * mat_B[8][14] +
                  mat_A[20][9] * mat_B[9][14] +
                  mat_A[20][10] * mat_B[10][14] +
                  mat_A[20][11] * mat_B[11][14] +
                  mat_A[20][12] * mat_B[12][14] +
                  mat_A[20][13] * mat_B[13][14] +
                  mat_A[20][14] * mat_B[14][14] +
                  mat_A[20][15] * mat_B[15][14] +
                  mat_A[20][16] * mat_B[16][14] +
                  mat_A[20][17] * mat_B[17][14] +
                  mat_A[20][18] * mat_B[18][14] +
                  mat_A[20][19] * mat_B[19][14] +
                  mat_A[20][20] * mat_B[20][14] +
                  mat_A[20][21] * mat_B[21][14] +
                  mat_A[20][22] * mat_B[22][14] +
                  mat_A[20][23] * mat_B[23][14] +
                  mat_A[20][24] * mat_B[24][14] +
                  mat_A[20][25] * mat_B[25][14] +
                  mat_A[20][26] * mat_B[26][14] +
                  mat_A[20][27] * mat_B[27][14] +
                  mat_A[20][28] * mat_B[28][14] +
                  mat_A[20][29] * mat_B[29][14] +
                  mat_A[20][30] * mat_B[30][14] +
                  mat_A[20][31] * mat_B[31][14];
    mat_C[20][15] <= 
                  mat_A[20][0] * mat_B[0][15] +
                  mat_A[20][1] * mat_B[1][15] +
                  mat_A[20][2] * mat_B[2][15] +
                  mat_A[20][3] * mat_B[3][15] +
                  mat_A[20][4] * mat_B[4][15] +
                  mat_A[20][5] * mat_B[5][15] +
                  mat_A[20][6] * mat_B[6][15] +
                  mat_A[20][7] * mat_B[7][15] +
                  mat_A[20][8] * mat_B[8][15] +
                  mat_A[20][9] * mat_B[9][15] +
                  mat_A[20][10] * mat_B[10][15] +
                  mat_A[20][11] * mat_B[11][15] +
                  mat_A[20][12] * mat_B[12][15] +
                  mat_A[20][13] * mat_B[13][15] +
                  mat_A[20][14] * mat_B[14][15] +
                  mat_A[20][15] * mat_B[15][15] +
                  mat_A[20][16] * mat_B[16][15] +
                  mat_A[20][17] * mat_B[17][15] +
                  mat_A[20][18] * mat_B[18][15] +
                  mat_A[20][19] * mat_B[19][15] +
                  mat_A[20][20] * mat_B[20][15] +
                  mat_A[20][21] * mat_B[21][15] +
                  mat_A[20][22] * mat_B[22][15] +
                  mat_A[20][23] * mat_B[23][15] +
                  mat_A[20][24] * mat_B[24][15] +
                  mat_A[20][25] * mat_B[25][15] +
                  mat_A[20][26] * mat_B[26][15] +
                  mat_A[20][27] * mat_B[27][15] +
                  mat_A[20][28] * mat_B[28][15] +
                  mat_A[20][29] * mat_B[29][15] +
                  mat_A[20][30] * mat_B[30][15] +
                  mat_A[20][31] * mat_B[31][15];
    mat_C[20][16] <= 
                  mat_A[20][0] * mat_B[0][16] +
                  mat_A[20][1] * mat_B[1][16] +
                  mat_A[20][2] * mat_B[2][16] +
                  mat_A[20][3] * mat_B[3][16] +
                  mat_A[20][4] * mat_B[4][16] +
                  mat_A[20][5] * mat_B[5][16] +
                  mat_A[20][6] * mat_B[6][16] +
                  mat_A[20][7] * mat_B[7][16] +
                  mat_A[20][8] * mat_B[8][16] +
                  mat_A[20][9] * mat_B[9][16] +
                  mat_A[20][10] * mat_B[10][16] +
                  mat_A[20][11] * mat_B[11][16] +
                  mat_A[20][12] * mat_B[12][16] +
                  mat_A[20][13] * mat_B[13][16] +
                  mat_A[20][14] * mat_B[14][16] +
                  mat_A[20][15] * mat_B[15][16] +
                  mat_A[20][16] * mat_B[16][16] +
                  mat_A[20][17] * mat_B[17][16] +
                  mat_A[20][18] * mat_B[18][16] +
                  mat_A[20][19] * mat_B[19][16] +
                  mat_A[20][20] * mat_B[20][16] +
                  mat_A[20][21] * mat_B[21][16] +
                  mat_A[20][22] * mat_B[22][16] +
                  mat_A[20][23] * mat_B[23][16] +
                  mat_A[20][24] * mat_B[24][16] +
                  mat_A[20][25] * mat_B[25][16] +
                  mat_A[20][26] * mat_B[26][16] +
                  mat_A[20][27] * mat_B[27][16] +
                  mat_A[20][28] * mat_B[28][16] +
                  mat_A[20][29] * mat_B[29][16] +
                  mat_A[20][30] * mat_B[30][16] +
                  mat_A[20][31] * mat_B[31][16];
    mat_C[20][17] <= 
                  mat_A[20][0] * mat_B[0][17] +
                  mat_A[20][1] * mat_B[1][17] +
                  mat_A[20][2] * mat_B[2][17] +
                  mat_A[20][3] * mat_B[3][17] +
                  mat_A[20][4] * mat_B[4][17] +
                  mat_A[20][5] * mat_B[5][17] +
                  mat_A[20][6] * mat_B[6][17] +
                  mat_A[20][7] * mat_B[7][17] +
                  mat_A[20][8] * mat_B[8][17] +
                  mat_A[20][9] * mat_B[9][17] +
                  mat_A[20][10] * mat_B[10][17] +
                  mat_A[20][11] * mat_B[11][17] +
                  mat_A[20][12] * mat_B[12][17] +
                  mat_A[20][13] * mat_B[13][17] +
                  mat_A[20][14] * mat_B[14][17] +
                  mat_A[20][15] * mat_B[15][17] +
                  mat_A[20][16] * mat_B[16][17] +
                  mat_A[20][17] * mat_B[17][17] +
                  mat_A[20][18] * mat_B[18][17] +
                  mat_A[20][19] * mat_B[19][17] +
                  mat_A[20][20] * mat_B[20][17] +
                  mat_A[20][21] * mat_B[21][17] +
                  mat_A[20][22] * mat_B[22][17] +
                  mat_A[20][23] * mat_B[23][17] +
                  mat_A[20][24] * mat_B[24][17] +
                  mat_A[20][25] * mat_B[25][17] +
                  mat_A[20][26] * mat_B[26][17] +
                  mat_A[20][27] * mat_B[27][17] +
                  mat_A[20][28] * mat_B[28][17] +
                  mat_A[20][29] * mat_B[29][17] +
                  mat_A[20][30] * mat_B[30][17] +
                  mat_A[20][31] * mat_B[31][17];
    mat_C[20][18] <= 
                  mat_A[20][0] * mat_B[0][18] +
                  mat_A[20][1] * mat_B[1][18] +
                  mat_A[20][2] * mat_B[2][18] +
                  mat_A[20][3] * mat_B[3][18] +
                  mat_A[20][4] * mat_B[4][18] +
                  mat_A[20][5] * mat_B[5][18] +
                  mat_A[20][6] * mat_B[6][18] +
                  mat_A[20][7] * mat_B[7][18] +
                  mat_A[20][8] * mat_B[8][18] +
                  mat_A[20][9] * mat_B[9][18] +
                  mat_A[20][10] * mat_B[10][18] +
                  mat_A[20][11] * mat_B[11][18] +
                  mat_A[20][12] * mat_B[12][18] +
                  mat_A[20][13] * mat_B[13][18] +
                  mat_A[20][14] * mat_B[14][18] +
                  mat_A[20][15] * mat_B[15][18] +
                  mat_A[20][16] * mat_B[16][18] +
                  mat_A[20][17] * mat_B[17][18] +
                  mat_A[20][18] * mat_B[18][18] +
                  mat_A[20][19] * mat_B[19][18] +
                  mat_A[20][20] * mat_B[20][18] +
                  mat_A[20][21] * mat_B[21][18] +
                  mat_A[20][22] * mat_B[22][18] +
                  mat_A[20][23] * mat_B[23][18] +
                  mat_A[20][24] * mat_B[24][18] +
                  mat_A[20][25] * mat_B[25][18] +
                  mat_A[20][26] * mat_B[26][18] +
                  mat_A[20][27] * mat_B[27][18] +
                  mat_A[20][28] * mat_B[28][18] +
                  mat_A[20][29] * mat_B[29][18] +
                  mat_A[20][30] * mat_B[30][18] +
                  mat_A[20][31] * mat_B[31][18];
    mat_C[20][19] <= 
                  mat_A[20][0] * mat_B[0][19] +
                  mat_A[20][1] * mat_B[1][19] +
                  mat_A[20][2] * mat_B[2][19] +
                  mat_A[20][3] * mat_B[3][19] +
                  mat_A[20][4] * mat_B[4][19] +
                  mat_A[20][5] * mat_B[5][19] +
                  mat_A[20][6] * mat_B[6][19] +
                  mat_A[20][7] * mat_B[7][19] +
                  mat_A[20][8] * mat_B[8][19] +
                  mat_A[20][9] * mat_B[9][19] +
                  mat_A[20][10] * mat_B[10][19] +
                  mat_A[20][11] * mat_B[11][19] +
                  mat_A[20][12] * mat_B[12][19] +
                  mat_A[20][13] * mat_B[13][19] +
                  mat_A[20][14] * mat_B[14][19] +
                  mat_A[20][15] * mat_B[15][19] +
                  mat_A[20][16] * mat_B[16][19] +
                  mat_A[20][17] * mat_B[17][19] +
                  mat_A[20][18] * mat_B[18][19] +
                  mat_A[20][19] * mat_B[19][19] +
                  mat_A[20][20] * mat_B[20][19] +
                  mat_A[20][21] * mat_B[21][19] +
                  mat_A[20][22] * mat_B[22][19] +
                  mat_A[20][23] * mat_B[23][19] +
                  mat_A[20][24] * mat_B[24][19] +
                  mat_A[20][25] * mat_B[25][19] +
                  mat_A[20][26] * mat_B[26][19] +
                  mat_A[20][27] * mat_B[27][19] +
                  mat_A[20][28] * mat_B[28][19] +
                  mat_A[20][29] * mat_B[29][19] +
                  mat_A[20][30] * mat_B[30][19] +
                  mat_A[20][31] * mat_B[31][19];
    mat_C[20][20] <= 
                  mat_A[20][0] * mat_B[0][20] +
                  mat_A[20][1] * mat_B[1][20] +
                  mat_A[20][2] * mat_B[2][20] +
                  mat_A[20][3] * mat_B[3][20] +
                  mat_A[20][4] * mat_B[4][20] +
                  mat_A[20][5] * mat_B[5][20] +
                  mat_A[20][6] * mat_B[6][20] +
                  mat_A[20][7] * mat_B[7][20] +
                  mat_A[20][8] * mat_B[8][20] +
                  mat_A[20][9] * mat_B[9][20] +
                  mat_A[20][10] * mat_B[10][20] +
                  mat_A[20][11] * mat_B[11][20] +
                  mat_A[20][12] * mat_B[12][20] +
                  mat_A[20][13] * mat_B[13][20] +
                  mat_A[20][14] * mat_B[14][20] +
                  mat_A[20][15] * mat_B[15][20] +
                  mat_A[20][16] * mat_B[16][20] +
                  mat_A[20][17] * mat_B[17][20] +
                  mat_A[20][18] * mat_B[18][20] +
                  mat_A[20][19] * mat_B[19][20] +
                  mat_A[20][20] * mat_B[20][20] +
                  mat_A[20][21] * mat_B[21][20] +
                  mat_A[20][22] * mat_B[22][20] +
                  mat_A[20][23] * mat_B[23][20] +
                  mat_A[20][24] * mat_B[24][20] +
                  mat_A[20][25] * mat_B[25][20] +
                  mat_A[20][26] * mat_B[26][20] +
                  mat_A[20][27] * mat_B[27][20] +
                  mat_A[20][28] * mat_B[28][20] +
                  mat_A[20][29] * mat_B[29][20] +
                  mat_A[20][30] * mat_B[30][20] +
                  mat_A[20][31] * mat_B[31][20];
    mat_C[20][21] <= 
                  mat_A[20][0] * mat_B[0][21] +
                  mat_A[20][1] * mat_B[1][21] +
                  mat_A[20][2] * mat_B[2][21] +
                  mat_A[20][3] * mat_B[3][21] +
                  mat_A[20][4] * mat_B[4][21] +
                  mat_A[20][5] * mat_B[5][21] +
                  mat_A[20][6] * mat_B[6][21] +
                  mat_A[20][7] * mat_B[7][21] +
                  mat_A[20][8] * mat_B[8][21] +
                  mat_A[20][9] * mat_B[9][21] +
                  mat_A[20][10] * mat_B[10][21] +
                  mat_A[20][11] * mat_B[11][21] +
                  mat_A[20][12] * mat_B[12][21] +
                  mat_A[20][13] * mat_B[13][21] +
                  mat_A[20][14] * mat_B[14][21] +
                  mat_A[20][15] * mat_B[15][21] +
                  mat_A[20][16] * mat_B[16][21] +
                  mat_A[20][17] * mat_B[17][21] +
                  mat_A[20][18] * mat_B[18][21] +
                  mat_A[20][19] * mat_B[19][21] +
                  mat_A[20][20] * mat_B[20][21] +
                  mat_A[20][21] * mat_B[21][21] +
                  mat_A[20][22] * mat_B[22][21] +
                  mat_A[20][23] * mat_B[23][21] +
                  mat_A[20][24] * mat_B[24][21] +
                  mat_A[20][25] * mat_B[25][21] +
                  mat_A[20][26] * mat_B[26][21] +
                  mat_A[20][27] * mat_B[27][21] +
                  mat_A[20][28] * mat_B[28][21] +
                  mat_A[20][29] * mat_B[29][21] +
                  mat_A[20][30] * mat_B[30][21] +
                  mat_A[20][31] * mat_B[31][21];
    mat_C[20][22] <= 
                  mat_A[20][0] * mat_B[0][22] +
                  mat_A[20][1] * mat_B[1][22] +
                  mat_A[20][2] * mat_B[2][22] +
                  mat_A[20][3] * mat_B[3][22] +
                  mat_A[20][4] * mat_B[4][22] +
                  mat_A[20][5] * mat_B[5][22] +
                  mat_A[20][6] * mat_B[6][22] +
                  mat_A[20][7] * mat_B[7][22] +
                  mat_A[20][8] * mat_B[8][22] +
                  mat_A[20][9] * mat_B[9][22] +
                  mat_A[20][10] * mat_B[10][22] +
                  mat_A[20][11] * mat_B[11][22] +
                  mat_A[20][12] * mat_B[12][22] +
                  mat_A[20][13] * mat_B[13][22] +
                  mat_A[20][14] * mat_B[14][22] +
                  mat_A[20][15] * mat_B[15][22] +
                  mat_A[20][16] * mat_B[16][22] +
                  mat_A[20][17] * mat_B[17][22] +
                  mat_A[20][18] * mat_B[18][22] +
                  mat_A[20][19] * mat_B[19][22] +
                  mat_A[20][20] * mat_B[20][22] +
                  mat_A[20][21] * mat_B[21][22] +
                  mat_A[20][22] * mat_B[22][22] +
                  mat_A[20][23] * mat_B[23][22] +
                  mat_A[20][24] * mat_B[24][22] +
                  mat_A[20][25] * mat_B[25][22] +
                  mat_A[20][26] * mat_B[26][22] +
                  mat_A[20][27] * mat_B[27][22] +
                  mat_A[20][28] * mat_B[28][22] +
                  mat_A[20][29] * mat_B[29][22] +
                  mat_A[20][30] * mat_B[30][22] +
                  mat_A[20][31] * mat_B[31][22];
    mat_C[20][23] <= 
                  mat_A[20][0] * mat_B[0][23] +
                  mat_A[20][1] * mat_B[1][23] +
                  mat_A[20][2] * mat_B[2][23] +
                  mat_A[20][3] * mat_B[3][23] +
                  mat_A[20][4] * mat_B[4][23] +
                  mat_A[20][5] * mat_B[5][23] +
                  mat_A[20][6] * mat_B[6][23] +
                  mat_A[20][7] * mat_B[7][23] +
                  mat_A[20][8] * mat_B[8][23] +
                  mat_A[20][9] * mat_B[9][23] +
                  mat_A[20][10] * mat_B[10][23] +
                  mat_A[20][11] * mat_B[11][23] +
                  mat_A[20][12] * mat_B[12][23] +
                  mat_A[20][13] * mat_B[13][23] +
                  mat_A[20][14] * mat_B[14][23] +
                  mat_A[20][15] * mat_B[15][23] +
                  mat_A[20][16] * mat_B[16][23] +
                  mat_A[20][17] * mat_B[17][23] +
                  mat_A[20][18] * mat_B[18][23] +
                  mat_A[20][19] * mat_B[19][23] +
                  mat_A[20][20] * mat_B[20][23] +
                  mat_A[20][21] * mat_B[21][23] +
                  mat_A[20][22] * mat_B[22][23] +
                  mat_A[20][23] * mat_B[23][23] +
                  mat_A[20][24] * mat_B[24][23] +
                  mat_A[20][25] * mat_B[25][23] +
                  mat_A[20][26] * mat_B[26][23] +
                  mat_A[20][27] * mat_B[27][23] +
                  mat_A[20][28] * mat_B[28][23] +
                  mat_A[20][29] * mat_B[29][23] +
                  mat_A[20][30] * mat_B[30][23] +
                  mat_A[20][31] * mat_B[31][23];
    mat_C[20][24] <= 
                  mat_A[20][0] * mat_B[0][24] +
                  mat_A[20][1] * mat_B[1][24] +
                  mat_A[20][2] * mat_B[2][24] +
                  mat_A[20][3] * mat_B[3][24] +
                  mat_A[20][4] * mat_B[4][24] +
                  mat_A[20][5] * mat_B[5][24] +
                  mat_A[20][6] * mat_B[6][24] +
                  mat_A[20][7] * mat_B[7][24] +
                  mat_A[20][8] * mat_B[8][24] +
                  mat_A[20][9] * mat_B[9][24] +
                  mat_A[20][10] * mat_B[10][24] +
                  mat_A[20][11] * mat_B[11][24] +
                  mat_A[20][12] * mat_B[12][24] +
                  mat_A[20][13] * mat_B[13][24] +
                  mat_A[20][14] * mat_B[14][24] +
                  mat_A[20][15] * mat_B[15][24] +
                  mat_A[20][16] * mat_B[16][24] +
                  mat_A[20][17] * mat_B[17][24] +
                  mat_A[20][18] * mat_B[18][24] +
                  mat_A[20][19] * mat_B[19][24] +
                  mat_A[20][20] * mat_B[20][24] +
                  mat_A[20][21] * mat_B[21][24] +
                  mat_A[20][22] * mat_B[22][24] +
                  mat_A[20][23] * mat_B[23][24] +
                  mat_A[20][24] * mat_B[24][24] +
                  mat_A[20][25] * mat_B[25][24] +
                  mat_A[20][26] * mat_B[26][24] +
                  mat_A[20][27] * mat_B[27][24] +
                  mat_A[20][28] * mat_B[28][24] +
                  mat_A[20][29] * mat_B[29][24] +
                  mat_A[20][30] * mat_B[30][24] +
                  mat_A[20][31] * mat_B[31][24];
    mat_C[20][25] <= 
                  mat_A[20][0] * mat_B[0][25] +
                  mat_A[20][1] * mat_B[1][25] +
                  mat_A[20][2] * mat_B[2][25] +
                  mat_A[20][3] * mat_B[3][25] +
                  mat_A[20][4] * mat_B[4][25] +
                  mat_A[20][5] * mat_B[5][25] +
                  mat_A[20][6] * mat_B[6][25] +
                  mat_A[20][7] * mat_B[7][25] +
                  mat_A[20][8] * mat_B[8][25] +
                  mat_A[20][9] * mat_B[9][25] +
                  mat_A[20][10] * mat_B[10][25] +
                  mat_A[20][11] * mat_B[11][25] +
                  mat_A[20][12] * mat_B[12][25] +
                  mat_A[20][13] * mat_B[13][25] +
                  mat_A[20][14] * mat_B[14][25] +
                  mat_A[20][15] * mat_B[15][25] +
                  mat_A[20][16] * mat_B[16][25] +
                  mat_A[20][17] * mat_B[17][25] +
                  mat_A[20][18] * mat_B[18][25] +
                  mat_A[20][19] * mat_B[19][25] +
                  mat_A[20][20] * mat_B[20][25] +
                  mat_A[20][21] * mat_B[21][25] +
                  mat_A[20][22] * mat_B[22][25] +
                  mat_A[20][23] * mat_B[23][25] +
                  mat_A[20][24] * mat_B[24][25] +
                  mat_A[20][25] * mat_B[25][25] +
                  mat_A[20][26] * mat_B[26][25] +
                  mat_A[20][27] * mat_B[27][25] +
                  mat_A[20][28] * mat_B[28][25] +
                  mat_A[20][29] * mat_B[29][25] +
                  mat_A[20][30] * mat_B[30][25] +
                  mat_A[20][31] * mat_B[31][25];
    mat_C[20][26] <= 
                  mat_A[20][0] * mat_B[0][26] +
                  mat_A[20][1] * mat_B[1][26] +
                  mat_A[20][2] * mat_B[2][26] +
                  mat_A[20][3] * mat_B[3][26] +
                  mat_A[20][4] * mat_B[4][26] +
                  mat_A[20][5] * mat_B[5][26] +
                  mat_A[20][6] * mat_B[6][26] +
                  mat_A[20][7] * mat_B[7][26] +
                  mat_A[20][8] * mat_B[8][26] +
                  mat_A[20][9] * mat_B[9][26] +
                  mat_A[20][10] * mat_B[10][26] +
                  mat_A[20][11] * mat_B[11][26] +
                  mat_A[20][12] * mat_B[12][26] +
                  mat_A[20][13] * mat_B[13][26] +
                  mat_A[20][14] * mat_B[14][26] +
                  mat_A[20][15] * mat_B[15][26] +
                  mat_A[20][16] * mat_B[16][26] +
                  mat_A[20][17] * mat_B[17][26] +
                  mat_A[20][18] * mat_B[18][26] +
                  mat_A[20][19] * mat_B[19][26] +
                  mat_A[20][20] * mat_B[20][26] +
                  mat_A[20][21] * mat_B[21][26] +
                  mat_A[20][22] * mat_B[22][26] +
                  mat_A[20][23] * mat_B[23][26] +
                  mat_A[20][24] * mat_B[24][26] +
                  mat_A[20][25] * mat_B[25][26] +
                  mat_A[20][26] * mat_B[26][26] +
                  mat_A[20][27] * mat_B[27][26] +
                  mat_A[20][28] * mat_B[28][26] +
                  mat_A[20][29] * mat_B[29][26] +
                  mat_A[20][30] * mat_B[30][26] +
                  mat_A[20][31] * mat_B[31][26];
    mat_C[20][27] <= 
                  mat_A[20][0] * mat_B[0][27] +
                  mat_A[20][1] * mat_B[1][27] +
                  mat_A[20][2] * mat_B[2][27] +
                  mat_A[20][3] * mat_B[3][27] +
                  mat_A[20][4] * mat_B[4][27] +
                  mat_A[20][5] * mat_B[5][27] +
                  mat_A[20][6] * mat_B[6][27] +
                  mat_A[20][7] * mat_B[7][27] +
                  mat_A[20][8] * mat_B[8][27] +
                  mat_A[20][9] * mat_B[9][27] +
                  mat_A[20][10] * mat_B[10][27] +
                  mat_A[20][11] * mat_B[11][27] +
                  mat_A[20][12] * mat_B[12][27] +
                  mat_A[20][13] * mat_B[13][27] +
                  mat_A[20][14] * mat_B[14][27] +
                  mat_A[20][15] * mat_B[15][27] +
                  mat_A[20][16] * mat_B[16][27] +
                  mat_A[20][17] * mat_B[17][27] +
                  mat_A[20][18] * mat_B[18][27] +
                  mat_A[20][19] * mat_B[19][27] +
                  mat_A[20][20] * mat_B[20][27] +
                  mat_A[20][21] * mat_B[21][27] +
                  mat_A[20][22] * mat_B[22][27] +
                  mat_A[20][23] * mat_B[23][27] +
                  mat_A[20][24] * mat_B[24][27] +
                  mat_A[20][25] * mat_B[25][27] +
                  mat_A[20][26] * mat_B[26][27] +
                  mat_A[20][27] * mat_B[27][27] +
                  mat_A[20][28] * mat_B[28][27] +
                  mat_A[20][29] * mat_B[29][27] +
                  mat_A[20][30] * mat_B[30][27] +
                  mat_A[20][31] * mat_B[31][27];
    mat_C[20][28] <= 
                  mat_A[20][0] * mat_B[0][28] +
                  mat_A[20][1] * mat_B[1][28] +
                  mat_A[20][2] * mat_B[2][28] +
                  mat_A[20][3] * mat_B[3][28] +
                  mat_A[20][4] * mat_B[4][28] +
                  mat_A[20][5] * mat_B[5][28] +
                  mat_A[20][6] * mat_B[6][28] +
                  mat_A[20][7] * mat_B[7][28] +
                  mat_A[20][8] * mat_B[8][28] +
                  mat_A[20][9] * mat_B[9][28] +
                  mat_A[20][10] * mat_B[10][28] +
                  mat_A[20][11] * mat_B[11][28] +
                  mat_A[20][12] * mat_B[12][28] +
                  mat_A[20][13] * mat_B[13][28] +
                  mat_A[20][14] * mat_B[14][28] +
                  mat_A[20][15] * mat_B[15][28] +
                  mat_A[20][16] * mat_B[16][28] +
                  mat_A[20][17] * mat_B[17][28] +
                  mat_A[20][18] * mat_B[18][28] +
                  mat_A[20][19] * mat_B[19][28] +
                  mat_A[20][20] * mat_B[20][28] +
                  mat_A[20][21] * mat_B[21][28] +
                  mat_A[20][22] * mat_B[22][28] +
                  mat_A[20][23] * mat_B[23][28] +
                  mat_A[20][24] * mat_B[24][28] +
                  mat_A[20][25] * mat_B[25][28] +
                  mat_A[20][26] * mat_B[26][28] +
                  mat_A[20][27] * mat_B[27][28] +
                  mat_A[20][28] * mat_B[28][28] +
                  mat_A[20][29] * mat_B[29][28] +
                  mat_A[20][30] * mat_B[30][28] +
                  mat_A[20][31] * mat_B[31][28];
    mat_C[20][29] <= 
                  mat_A[20][0] * mat_B[0][29] +
                  mat_A[20][1] * mat_B[1][29] +
                  mat_A[20][2] * mat_B[2][29] +
                  mat_A[20][3] * mat_B[3][29] +
                  mat_A[20][4] * mat_B[4][29] +
                  mat_A[20][5] * mat_B[5][29] +
                  mat_A[20][6] * mat_B[6][29] +
                  mat_A[20][7] * mat_B[7][29] +
                  mat_A[20][8] * mat_B[8][29] +
                  mat_A[20][9] * mat_B[9][29] +
                  mat_A[20][10] * mat_B[10][29] +
                  mat_A[20][11] * mat_B[11][29] +
                  mat_A[20][12] * mat_B[12][29] +
                  mat_A[20][13] * mat_B[13][29] +
                  mat_A[20][14] * mat_B[14][29] +
                  mat_A[20][15] * mat_B[15][29] +
                  mat_A[20][16] * mat_B[16][29] +
                  mat_A[20][17] * mat_B[17][29] +
                  mat_A[20][18] * mat_B[18][29] +
                  mat_A[20][19] * mat_B[19][29] +
                  mat_A[20][20] * mat_B[20][29] +
                  mat_A[20][21] * mat_B[21][29] +
                  mat_A[20][22] * mat_B[22][29] +
                  mat_A[20][23] * mat_B[23][29] +
                  mat_A[20][24] * mat_B[24][29] +
                  mat_A[20][25] * mat_B[25][29] +
                  mat_A[20][26] * mat_B[26][29] +
                  mat_A[20][27] * mat_B[27][29] +
                  mat_A[20][28] * mat_B[28][29] +
                  mat_A[20][29] * mat_B[29][29] +
                  mat_A[20][30] * mat_B[30][29] +
                  mat_A[20][31] * mat_B[31][29];
    mat_C[20][30] <= 
                  mat_A[20][0] * mat_B[0][30] +
                  mat_A[20][1] * mat_B[1][30] +
                  mat_A[20][2] * mat_B[2][30] +
                  mat_A[20][3] * mat_B[3][30] +
                  mat_A[20][4] * mat_B[4][30] +
                  mat_A[20][5] * mat_B[5][30] +
                  mat_A[20][6] * mat_B[6][30] +
                  mat_A[20][7] * mat_B[7][30] +
                  mat_A[20][8] * mat_B[8][30] +
                  mat_A[20][9] * mat_B[9][30] +
                  mat_A[20][10] * mat_B[10][30] +
                  mat_A[20][11] * mat_B[11][30] +
                  mat_A[20][12] * mat_B[12][30] +
                  mat_A[20][13] * mat_B[13][30] +
                  mat_A[20][14] * mat_B[14][30] +
                  mat_A[20][15] * mat_B[15][30] +
                  mat_A[20][16] * mat_B[16][30] +
                  mat_A[20][17] * mat_B[17][30] +
                  mat_A[20][18] * mat_B[18][30] +
                  mat_A[20][19] * mat_B[19][30] +
                  mat_A[20][20] * mat_B[20][30] +
                  mat_A[20][21] * mat_B[21][30] +
                  mat_A[20][22] * mat_B[22][30] +
                  mat_A[20][23] * mat_B[23][30] +
                  mat_A[20][24] * mat_B[24][30] +
                  mat_A[20][25] * mat_B[25][30] +
                  mat_A[20][26] * mat_B[26][30] +
                  mat_A[20][27] * mat_B[27][30] +
                  mat_A[20][28] * mat_B[28][30] +
                  mat_A[20][29] * mat_B[29][30] +
                  mat_A[20][30] * mat_B[30][30] +
                  mat_A[20][31] * mat_B[31][30];
    mat_C[20][31] <= 
                  mat_A[20][0] * mat_B[0][31] +
                  mat_A[20][1] * mat_B[1][31] +
                  mat_A[20][2] * mat_B[2][31] +
                  mat_A[20][3] * mat_B[3][31] +
                  mat_A[20][4] * mat_B[4][31] +
                  mat_A[20][5] * mat_B[5][31] +
                  mat_A[20][6] * mat_B[6][31] +
                  mat_A[20][7] * mat_B[7][31] +
                  mat_A[20][8] * mat_B[8][31] +
                  mat_A[20][9] * mat_B[9][31] +
                  mat_A[20][10] * mat_B[10][31] +
                  mat_A[20][11] * mat_B[11][31] +
                  mat_A[20][12] * mat_B[12][31] +
                  mat_A[20][13] * mat_B[13][31] +
                  mat_A[20][14] * mat_B[14][31] +
                  mat_A[20][15] * mat_B[15][31] +
                  mat_A[20][16] * mat_B[16][31] +
                  mat_A[20][17] * mat_B[17][31] +
                  mat_A[20][18] * mat_B[18][31] +
                  mat_A[20][19] * mat_B[19][31] +
                  mat_A[20][20] * mat_B[20][31] +
                  mat_A[20][21] * mat_B[21][31] +
                  mat_A[20][22] * mat_B[22][31] +
                  mat_A[20][23] * mat_B[23][31] +
                  mat_A[20][24] * mat_B[24][31] +
                  mat_A[20][25] * mat_B[25][31] +
                  mat_A[20][26] * mat_B[26][31] +
                  mat_A[20][27] * mat_B[27][31] +
                  mat_A[20][28] * mat_B[28][31] +
                  mat_A[20][29] * mat_B[29][31] +
                  mat_A[20][30] * mat_B[30][31] +
                  mat_A[20][31] * mat_B[31][31];
    mat_C[21][0] <= 
                  mat_A[21][0] * mat_B[0][0] +
                  mat_A[21][1] * mat_B[1][0] +
                  mat_A[21][2] * mat_B[2][0] +
                  mat_A[21][3] * mat_B[3][0] +
                  mat_A[21][4] * mat_B[4][0] +
                  mat_A[21][5] * mat_B[5][0] +
                  mat_A[21][6] * mat_B[6][0] +
                  mat_A[21][7] * mat_B[7][0] +
                  mat_A[21][8] * mat_B[8][0] +
                  mat_A[21][9] * mat_B[9][0] +
                  mat_A[21][10] * mat_B[10][0] +
                  mat_A[21][11] * mat_B[11][0] +
                  mat_A[21][12] * mat_B[12][0] +
                  mat_A[21][13] * mat_B[13][0] +
                  mat_A[21][14] * mat_B[14][0] +
                  mat_A[21][15] * mat_B[15][0] +
                  mat_A[21][16] * mat_B[16][0] +
                  mat_A[21][17] * mat_B[17][0] +
                  mat_A[21][18] * mat_B[18][0] +
                  mat_A[21][19] * mat_B[19][0] +
                  mat_A[21][20] * mat_B[20][0] +
                  mat_A[21][21] * mat_B[21][0] +
                  mat_A[21][22] * mat_B[22][0] +
                  mat_A[21][23] * mat_B[23][0] +
                  mat_A[21][24] * mat_B[24][0] +
                  mat_A[21][25] * mat_B[25][0] +
                  mat_A[21][26] * mat_B[26][0] +
                  mat_A[21][27] * mat_B[27][0] +
                  mat_A[21][28] * mat_B[28][0] +
                  mat_A[21][29] * mat_B[29][0] +
                  mat_A[21][30] * mat_B[30][0] +
                  mat_A[21][31] * mat_B[31][0];
    mat_C[21][1] <= 
                  mat_A[21][0] * mat_B[0][1] +
                  mat_A[21][1] * mat_B[1][1] +
                  mat_A[21][2] * mat_B[2][1] +
                  mat_A[21][3] * mat_B[3][1] +
                  mat_A[21][4] * mat_B[4][1] +
                  mat_A[21][5] * mat_B[5][1] +
                  mat_A[21][6] * mat_B[6][1] +
                  mat_A[21][7] * mat_B[7][1] +
                  mat_A[21][8] * mat_B[8][1] +
                  mat_A[21][9] * mat_B[9][1] +
                  mat_A[21][10] * mat_B[10][1] +
                  mat_A[21][11] * mat_B[11][1] +
                  mat_A[21][12] * mat_B[12][1] +
                  mat_A[21][13] * mat_B[13][1] +
                  mat_A[21][14] * mat_B[14][1] +
                  mat_A[21][15] * mat_B[15][1] +
                  mat_A[21][16] * mat_B[16][1] +
                  mat_A[21][17] * mat_B[17][1] +
                  mat_A[21][18] * mat_B[18][1] +
                  mat_A[21][19] * mat_B[19][1] +
                  mat_A[21][20] * mat_B[20][1] +
                  mat_A[21][21] * mat_B[21][1] +
                  mat_A[21][22] * mat_B[22][1] +
                  mat_A[21][23] * mat_B[23][1] +
                  mat_A[21][24] * mat_B[24][1] +
                  mat_A[21][25] * mat_B[25][1] +
                  mat_A[21][26] * mat_B[26][1] +
                  mat_A[21][27] * mat_B[27][1] +
                  mat_A[21][28] * mat_B[28][1] +
                  mat_A[21][29] * mat_B[29][1] +
                  mat_A[21][30] * mat_B[30][1] +
                  mat_A[21][31] * mat_B[31][1];
    mat_C[21][2] <= 
                  mat_A[21][0] * mat_B[0][2] +
                  mat_A[21][1] * mat_B[1][2] +
                  mat_A[21][2] * mat_B[2][2] +
                  mat_A[21][3] * mat_B[3][2] +
                  mat_A[21][4] * mat_B[4][2] +
                  mat_A[21][5] * mat_B[5][2] +
                  mat_A[21][6] * mat_B[6][2] +
                  mat_A[21][7] * mat_B[7][2] +
                  mat_A[21][8] * mat_B[8][2] +
                  mat_A[21][9] * mat_B[9][2] +
                  mat_A[21][10] * mat_B[10][2] +
                  mat_A[21][11] * mat_B[11][2] +
                  mat_A[21][12] * mat_B[12][2] +
                  mat_A[21][13] * mat_B[13][2] +
                  mat_A[21][14] * mat_B[14][2] +
                  mat_A[21][15] * mat_B[15][2] +
                  mat_A[21][16] * mat_B[16][2] +
                  mat_A[21][17] * mat_B[17][2] +
                  mat_A[21][18] * mat_B[18][2] +
                  mat_A[21][19] * mat_B[19][2] +
                  mat_A[21][20] * mat_B[20][2] +
                  mat_A[21][21] * mat_B[21][2] +
                  mat_A[21][22] * mat_B[22][2] +
                  mat_A[21][23] * mat_B[23][2] +
                  mat_A[21][24] * mat_B[24][2] +
                  mat_A[21][25] * mat_B[25][2] +
                  mat_A[21][26] * mat_B[26][2] +
                  mat_A[21][27] * mat_B[27][2] +
                  mat_A[21][28] * mat_B[28][2] +
                  mat_A[21][29] * mat_B[29][2] +
                  mat_A[21][30] * mat_B[30][2] +
                  mat_A[21][31] * mat_B[31][2];
    mat_C[21][3] <= 
                  mat_A[21][0] * mat_B[0][3] +
                  mat_A[21][1] * mat_B[1][3] +
                  mat_A[21][2] * mat_B[2][3] +
                  mat_A[21][3] * mat_B[3][3] +
                  mat_A[21][4] * mat_B[4][3] +
                  mat_A[21][5] * mat_B[5][3] +
                  mat_A[21][6] * mat_B[6][3] +
                  mat_A[21][7] * mat_B[7][3] +
                  mat_A[21][8] * mat_B[8][3] +
                  mat_A[21][9] * mat_B[9][3] +
                  mat_A[21][10] * mat_B[10][3] +
                  mat_A[21][11] * mat_B[11][3] +
                  mat_A[21][12] * mat_B[12][3] +
                  mat_A[21][13] * mat_B[13][3] +
                  mat_A[21][14] * mat_B[14][3] +
                  mat_A[21][15] * mat_B[15][3] +
                  mat_A[21][16] * mat_B[16][3] +
                  mat_A[21][17] * mat_B[17][3] +
                  mat_A[21][18] * mat_B[18][3] +
                  mat_A[21][19] * mat_B[19][3] +
                  mat_A[21][20] * mat_B[20][3] +
                  mat_A[21][21] * mat_B[21][3] +
                  mat_A[21][22] * mat_B[22][3] +
                  mat_A[21][23] * mat_B[23][3] +
                  mat_A[21][24] * mat_B[24][3] +
                  mat_A[21][25] * mat_B[25][3] +
                  mat_A[21][26] * mat_B[26][3] +
                  mat_A[21][27] * mat_B[27][3] +
                  mat_A[21][28] * mat_B[28][3] +
                  mat_A[21][29] * mat_B[29][3] +
                  mat_A[21][30] * mat_B[30][3] +
                  mat_A[21][31] * mat_B[31][3];
    mat_C[21][4] <= 
                  mat_A[21][0] * mat_B[0][4] +
                  mat_A[21][1] * mat_B[1][4] +
                  mat_A[21][2] * mat_B[2][4] +
                  mat_A[21][3] * mat_B[3][4] +
                  mat_A[21][4] * mat_B[4][4] +
                  mat_A[21][5] * mat_B[5][4] +
                  mat_A[21][6] * mat_B[6][4] +
                  mat_A[21][7] * mat_B[7][4] +
                  mat_A[21][8] * mat_B[8][4] +
                  mat_A[21][9] * mat_B[9][4] +
                  mat_A[21][10] * mat_B[10][4] +
                  mat_A[21][11] * mat_B[11][4] +
                  mat_A[21][12] * mat_B[12][4] +
                  mat_A[21][13] * mat_B[13][4] +
                  mat_A[21][14] * mat_B[14][4] +
                  mat_A[21][15] * mat_B[15][4] +
                  mat_A[21][16] * mat_B[16][4] +
                  mat_A[21][17] * mat_B[17][4] +
                  mat_A[21][18] * mat_B[18][4] +
                  mat_A[21][19] * mat_B[19][4] +
                  mat_A[21][20] * mat_B[20][4] +
                  mat_A[21][21] * mat_B[21][4] +
                  mat_A[21][22] * mat_B[22][4] +
                  mat_A[21][23] * mat_B[23][4] +
                  mat_A[21][24] * mat_B[24][4] +
                  mat_A[21][25] * mat_B[25][4] +
                  mat_A[21][26] * mat_B[26][4] +
                  mat_A[21][27] * mat_B[27][4] +
                  mat_A[21][28] * mat_B[28][4] +
                  mat_A[21][29] * mat_B[29][4] +
                  mat_A[21][30] * mat_B[30][4] +
                  mat_A[21][31] * mat_B[31][4];
    mat_C[21][5] <= 
                  mat_A[21][0] * mat_B[0][5] +
                  mat_A[21][1] * mat_B[1][5] +
                  mat_A[21][2] * mat_B[2][5] +
                  mat_A[21][3] * mat_B[3][5] +
                  mat_A[21][4] * mat_B[4][5] +
                  mat_A[21][5] * mat_B[5][5] +
                  mat_A[21][6] * mat_B[6][5] +
                  mat_A[21][7] * mat_B[7][5] +
                  mat_A[21][8] * mat_B[8][5] +
                  mat_A[21][9] * mat_B[9][5] +
                  mat_A[21][10] * mat_B[10][5] +
                  mat_A[21][11] * mat_B[11][5] +
                  mat_A[21][12] * mat_B[12][5] +
                  mat_A[21][13] * mat_B[13][5] +
                  mat_A[21][14] * mat_B[14][5] +
                  mat_A[21][15] * mat_B[15][5] +
                  mat_A[21][16] * mat_B[16][5] +
                  mat_A[21][17] * mat_B[17][5] +
                  mat_A[21][18] * mat_B[18][5] +
                  mat_A[21][19] * mat_B[19][5] +
                  mat_A[21][20] * mat_B[20][5] +
                  mat_A[21][21] * mat_B[21][5] +
                  mat_A[21][22] * mat_B[22][5] +
                  mat_A[21][23] * mat_B[23][5] +
                  mat_A[21][24] * mat_B[24][5] +
                  mat_A[21][25] * mat_B[25][5] +
                  mat_A[21][26] * mat_B[26][5] +
                  mat_A[21][27] * mat_B[27][5] +
                  mat_A[21][28] * mat_B[28][5] +
                  mat_A[21][29] * mat_B[29][5] +
                  mat_A[21][30] * mat_B[30][5] +
                  mat_A[21][31] * mat_B[31][5];
    mat_C[21][6] <= 
                  mat_A[21][0] * mat_B[0][6] +
                  mat_A[21][1] * mat_B[1][6] +
                  mat_A[21][2] * mat_B[2][6] +
                  mat_A[21][3] * mat_B[3][6] +
                  mat_A[21][4] * mat_B[4][6] +
                  mat_A[21][5] * mat_B[5][6] +
                  mat_A[21][6] * mat_B[6][6] +
                  mat_A[21][7] * mat_B[7][6] +
                  mat_A[21][8] * mat_B[8][6] +
                  mat_A[21][9] * mat_B[9][6] +
                  mat_A[21][10] * mat_B[10][6] +
                  mat_A[21][11] * mat_B[11][6] +
                  mat_A[21][12] * mat_B[12][6] +
                  mat_A[21][13] * mat_B[13][6] +
                  mat_A[21][14] * mat_B[14][6] +
                  mat_A[21][15] * mat_B[15][6] +
                  mat_A[21][16] * mat_B[16][6] +
                  mat_A[21][17] * mat_B[17][6] +
                  mat_A[21][18] * mat_B[18][6] +
                  mat_A[21][19] * mat_B[19][6] +
                  mat_A[21][20] * mat_B[20][6] +
                  mat_A[21][21] * mat_B[21][6] +
                  mat_A[21][22] * mat_B[22][6] +
                  mat_A[21][23] * mat_B[23][6] +
                  mat_A[21][24] * mat_B[24][6] +
                  mat_A[21][25] * mat_B[25][6] +
                  mat_A[21][26] * mat_B[26][6] +
                  mat_A[21][27] * mat_B[27][6] +
                  mat_A[21][28] * mat_B[28][6] +
                  mat_A[21][29] * mat_B[29][6] +
                  mat_A[21][30] * mat_B[30][6] +
                  mat_A[21][31] * mat_B[31][6];
    mat_C[21][7] <= 
                  mat_A[21][0] * mat_B[0][7] +
                  mat_A[21][1] * mat_B[1][7] +
                  mat_A[21][2] * mat_B[2][7] +
                  mat_A[21][3] * mat_B[3][7] +
                  mat_A[21][4] * mat_B[4][7] +
                  mat_A[21][5] * mat_B[5][7] +
                  mat_A[21][6] * mat_B[6][7] +
                  mat_A[21][7] * mat_B[7][7] +
                  mat_A[21][8] * mat_B[8][7] +
                  mat_A[21][9] * mat_B[9][7] +
                  mat_A[21][10] * mat_B[10][7] +
                  mat_A[21][11] * mat_B[11][7] +
                  mat_A[21][12] * mat_B[12][7] +
                  mat_A[21][13] * mat_B[13][7] +
                  mat_A[21][14] * mat_B[14][7] +
                  mat_A[21][15] * mat_B[15][7] +
                  mat_A[21][16] * mat_B[16][7] +
                  mat_A[21][17] * mat_B[17][7] +
                  mat_A[21][18] * mat_B[18][7] +
                  mat_A[21][19] * mat_B[19][7] +
                  mat_A[21][20] * mat_B[20][7] +
                  mat_A[21][21] * mat_B[21][7] +
                  mat_A[21][22] * mat_B[22][7] +
                  mat_A[21][23] * mat_B[23][7] +
                  mat_A[21][24] * mat_B[24][7] +
                  mat_A[21][25] * mat_B[25][7] +
                  mat_A[21][26] * mat_B[26][7] +
                  mat_A[21][27] * mat_B[27][7] +
                  mat_A[21][28] * mat_B[28][7] +
                  mat_A[21][29] * mat_B[29][7] +
                  mat_A[21][30] * mat_B[30][7] +
                  mat_A[21][31] * mat_B[31][7];
    mat_C[21][8] <= 
                  mat_A[21][0] * mat_B[0][8] +
                  mat_A[21][1] * mat_B[1][8] +
                  mat_A[21][2] * mat_B[2][8] +
                  mat_A[21][3] * mat_B[3][8] +
                  mat_A[21][4] * mat_B[4][8] +
                  mat_A[21][5] * mat_B[5][8] +
                  mat_A[21][6] * mat_B[6][8] +
                  mat_A[21][7] * mat_B[7][8] +
                  mat_A[21][8] * mat_B[8][8] +
                  mat_A[21][9] * mat_B[9][8] +
                  mat_A[21][10] * mat_B[10][8] +
                  mat_A[21][11] * mat_B[11][8] +
                  mat_A[21][12] * mat_B[12][8] +
                  mat_A[21][13] * mat_B[13][8] +
                  mat_A[21][14] * mat_B[14][8] +
                  mat_A[21][15] * mat_B[15][8] +
                  mat_A[21][16] * mat_B[16][8] +
                  mat_A[21][17] * mat_B[17][8] +
                  mat_A[21][18] * mat_B[18][8] +
                  mat_A[21][19] * mat_B[19][8] +
                  mat_A[21][20] * mat_B[20][8] +
                  mat_A[21][21] * mat_B[21][8] +
                  mat_A[21][22] * mat_B[22][8] +
                  mat_A[21][23] * mat_B[23][8] +
                  mat_A[21][24] * mat_B[24][8] +
                  mat_A[21][25] * mat_B[25][8] +
                  mat_A[21][26] * mat_B[26][8] +
                  mat_A[21][27] * mat_B[27][8] +
                  mat_A[21][28] * mat_B[28][8] +
                  mat_A[21][29] * mat_B[29][8] +
                  mat_A[21][30] * mat_B[30][8] +
                  mat_A[21][31] * mat_B[31][8];
    mat_C[21][9] <= 
                  mat_A[21][0] * mat_B[0][9] +
                  mat_A[21][1] * mat_B[1][9] +
                  mat_A[21][2] * mat_B[2][9] +
                  mat_A[21][3] * mat_B[3][9] +
                  mat_A[21][4] * mat_B[4][9] +
                  mat_A[21][5] * mat_B[5][9] +
                  mat_A[21][6] * mat_B[6][9] +
                  mat_A[21][7] * mat_B[7][9] +
                  mat_A[21][8] * mat_B[8][9] +
                  mat_A[21][9] * mat_B[9][9] +
                  mat_A[21][10] * mat_B[10][9] +
                  mat_A[21][11] * mat_B[11][9] +
                  mat_A[21][12] * mat_B[12][9] +
                  mat_A[21][13] * mat_B[13][9] +
                  mat_A[21][14] * mat_B[14][9] +
                  mat_A[21][15] * mat_B[15][9] +
                  mat_A[21][16] * mat_B[16][9] +
                  mat_A[21][17] * mat_B[17][9] +
                  mat_A[21][18] * mat_B[18][9] +
                  mat_A[21][19] * mat_B[19][9] +
                  mat_A[21][20] * mat_B[20][9] +
                  mat_A[21][21] * mat_B[21][9] +
                  mat_A[21][22] * mat_B[22][9] +
                  mat_A[21][23] * mat_B[23][9] +
                  mat_A[21][24] * mat_B[24][9] +
                  mat_A[21][25] * mat_B[25][9] +
                  mat_A[21][26] * mat_B[26][9] +
                  mat_A[21][27] * mat_B[27][9] +
                  mat_A[21][28] * mat_B[28][9] +
                  mat_A[21][29] * mat_B[29][9] +
                  mat_A[21][30] * mat_B[30][9] +
                  mat_A[21][31] * mat_B[31][9];
    mat_C[21][10] <= 
                  mat_A[21][0] * mat_B[0][10] +
                  mat_A[21][1] * mat_B[1][10] +
                  mat_A[21][2] * mat_B[2][10] +
                  mat_A[21][3] * mat_B[3][10] +
                  mat_A[21][4] * mat_B[4][10] +
                  mat_A[21][5] * mat_B[5][10] +
                  mat_A[21][6] * mat_B[6][10] +
                  mat_A[21][7] * mat_B[7][10] +
                  mat_A[21][8] * mat_B[8][10] +
                  mat_A[21][9] * mat_B[9][10] +
                  mat_A[21][10] * mat_B[10][10] +
                  mat_A[21][11] * mat_B[11][10] +
                  mat_A[21][12] * mat_B[12][10] +
                  mat_A[21][13] * mat_B[13][10] +
                  mat_A[21][14] * mat_B[14][10] +
                  mat_A[21][15] * mat_B[15][10] +
                  mat_A[21][16] * mat_B[16][10] +
                  mat_A[21][17] * mat_B[17][10] +
                  mat_A[21][18] * mat_B[18][10] +
                  mat_A[21][19] * mat_B[19][10] +
                  mat_A[21][20] * mat_B[20][10] +
                  mat_A[21][21] * mat_B[21][10] +
                  mat_A[21][22] * mat_B[22][10] +
                  mat_A[21][23] * mat_B[23][10] +
                  mat_A[21][24] * mat_B[24][10] +
                  mat_A[21][25] * mat_B[25][10] +
                  mat_A[21][26] * mat_B[26][10] +
                  mat_A[21][27] * mat_B[27][10] +
                  mat_A[21][28] * mat_B[28][10] +
                  mat_A[21][29] * mat_B[29][10] +
                  mat_A[21][30] * mat_B[30][10] +
                  mat_A[21][31] * mat_B[31][10];
    mat_C[21][11] <= 
                  mat_A[21][0] * mat_B[0][11] +
                  mat_A[21][1] * mat_B[1][11] +
                  mat_A[21][2] * mat_B[2][11] +
                  mat_A[21][3] * mat_B[3][11] +
                  mat_A[21][4] * mat_B[4][11] +
                  mat_A[21][5] * mat_B[5][11] +
                  mat_A[21][6] * mat_B[6][11] +
                  mat_A[21][7] * mat_B[7][11] +
                  mat_A[21][8] * mat_B[8][11] +
                  mat_A[21][9] * mat_B[9][11] +
                  mat_A[21][10] * mat_B[10][11] +
                  mat_A[21][11] * mat_B[11][11] +
                  mat_A[21][12] * mat_B[12][11] +
                  mat_A[21][13] * mat_B[13][11] +
                  mat_A[21][14] * mat_B[14][11] +
                  mat_A[21][15] * mat_B[15][11] +
                  mat_A[21][16] * mat_B[16][11] +
                  mat_A[21][17] * mat_B[17][11] +
                  mat_A[21][18] * mat_B[18][11] +
                  mat_A[21][19] * mat_B[19][11] +
                  mat_A[21][20] * mat_B[20][11] +
                  mat_A[21][21] * mat_B[21][11] +
                  mat_A[21][22] * mat_B[22][11] +
                  mat_A[21][23] * mat_B[23][11] +
                  mat_A[21][24] * mat_B[24][11] +
                  mat_A[21][25] * mat_B[25][11] +
                  mat_A[21][26] * mat_B[26][11] +
                  mat_A[21][27] * mat_B[27][11] +
                  mat_A[21][28] * mat_B[28][11] +
                  mat_A[21][29] * mat_B[29][11] +
                  mat_A[21][30] * mat_B[30][11] +
                  mat_A[21][31] * mat_B[31][11];
    mat_C[21][12] <= 
                  mat_A[21][0] * mat_B[0][12] +
                  mat_A[21][1] * mat_B[1][12] +
                  mat_A[21][2] * mat_B[2][12] +
                  mat_A[21][3] * mat_B[3][12] +
                  mat_A[21][4] * mat_B[4][12] +
                  mat_A[21][5] * mat_B[5][12] +
                  mat_A[21][6] * mat_B[6][12] +
                  mat_A[21][7] * mat_B[7][12] +
                  mat_A[21][8] * mat_B[8][12] +
                  mat_A[21][9] * mat_B[9][12] +
                  mat_A[21][10] * mat_B[10][12] +
                  mat_A[21][11] * mat_B[11][12] +
                  mat_A[21][12] * mat_B[12][12] +
                  mat_A[21][13] * mat_B[13][12] +
                  mat_A[21][14] * mat_B[14][12] +
                  mat_A[21][15] * mat_B[15][12] +
                  mat_A[21][16] * mat_B[16][12] +
                  mat_A[21][17] * mat_B[17][12] +
                  mat_A[21][18] * mat_B[18][12] +
                  mat_A[21][19] * mat_B[19][12] +
                  mat_A[21][20] * mat_B[20][12] +
                  mat_A[21][21] * mat_B[21][12] +
                  mat_A[21][22] * mat_B[22][12] +
                  mat_A[21][23] * mat_B[23][12] +
                  mat_A[21][24] * mat_B[24][12] +
                  mat_A[21][25] * mat_B[25][12] +
                  mat_A[21][26] * mat_B[26][12] +
                  mat_A[21][27] * mat_B[27][12] +
                  mat_A[21][28] * mat_B[28][12] +
                  mat_A[21][29] * mat_B[29][12] +
                  mat_A[21][30] * mat_B[30][12] +
                  mat_A[21][31] * mat_B[31][12];
    mat_C[21][13] <= 
                  mat_A[21][0] * mat_B[0][13] +
                  mat_A[21][1] * mat_B[1][13] +
                  mat_A[21][2] * mat_B[2][13] +
                  mat_A[21][3] * mat_B[3][13] +
                  mat_A[21][4] * mat_B[4][13] +
                  mat_A[21][5] * mat_B[5][13] +
                  mat_A[21][6] * mat_B[6][13] +
                  mat_A[21][7] * mat_B[7][13] +
                  mat_A[21][8] * mat_B[8][13] +
                  mat_A[21][9] * mat_B[9][13] +
                  mat_A[21][10] * mat_B[10][13] +
                  mat_A[21][11] * mat_B[11][13] +
                  mat_A[21][12] * mat_B[12][13] +
                  mat_A[21][13] * mat_B[13][13] +
                  mat_A[21][14] * mat_B[14][13] +
                  mat_A[21][15] * mat_B[15][13] +
                  mat_A[21][16] * mat_B[16][13] +
                  mat_A[21][17] * mat_B[17][13] +
                  mat_A[21][18] * mat_B[18][13] +
                  mat_A[21][19] * mat_B[19][13] +
                  mat_A[21][20] * mat_B[20][13] +
                  mat_A[21][21] * mat_B[21][13] +
                  mat_A[21][22] * mat_B[22][13] +
                  mat_A[21][23] * mat_B[23][13] +
                  mat_A[21][24] * mat_B[24][13] +
                  mat_A[21][25] * mat_B[25][13] +
                  mat_A[21][26] * mat_B[26][13] +
                  mat_A[21][27] * mat_B[27][13] +
                  mat_A[21][28] * mat_B[28][13] +
                  mat_A[21][29] * mat_B[29][13] +
                  mat_A[21][30] * mat_B[30][13] +
                  mat_A[21][31] * mat_B[31][13];
    mat_C[21][14] <= 
                  mat_A[21][0] * mat_B[0][14] +
                  mat_A[21][1] * mat_B[1][14] +
                  mat_A[21][2] * mat_B[2][14] +
                  mat_A[21][3] * mat_B[3][14] +
                  mat_A[21][4] * mat_B[4][14] +
                  mat_A[21][5] * mat_B[5][14] +
                  mat_A[21][6] * mat_B[6][14] +
                  mat_A[21][7] * mat_B[7][14] +
                  mat_A[21][8] * mat_B[8][14] +
                  mat_A[21][9] * mat_B[9][14] +
                  mat_A[21][10] * mat_B[10][14] +
                  mat_A[21][11] * mat_B[11][14] +
                  mat_A[21][12] * mat_B[12][14] +
                  mat_A[21][13] * mat_B[13][14] +
                  mat_A[21][14] * mat_B[14][14] +
                  mat_A[21][15] * mat_B[15][14] +
                  mat_A[21][16] * mat_B[16][14] +
                  mat_A[21][17] * mat_B[17][14] +
                  mat_A[21][18] * mat_B[18][14] +
                  mat_A[21][19] * mat_B[19][14] +
                  mat_A[21][20] * mat_B[20][14] +
                  mat_A[21][21] * mat_B[21][14] +
                  mat_A[21][22] * mat_B[22][14] +
                  mat_A[21][23] * mat_B[23][14] +
                  mat_A[21][24] * mat_B[24][14] +
                  mat_A[21][25] * mat_B[25][14] +
                  mat_A[21][26] * mat_B[26][14] +
                  mat_A[21][27] * mat_B[27][14] +
                  mat_A[21][28] * mat_B[28][14] +
                  mat_A[21][29] * mat_B[29][14] +
                  mat_A[21][30] * mat_B[30][14] +
                  mat_A[21][31] * mat_B[31][14];
    mat_C[21][15] <= 
                  mat_A[21][0] * mat_B[0][15] +
                  mat_A[21][1] * mat_B[1][15] +
                  mat_A[21][2] * mat_B[2][15] +
                  mat_A[21][3] * mat_B[3][15] +
                  mat_A[21][4] * mat_B[4][15] +
                  mat_A[21][5] * mat_B[5][15] +
                  mat_A[21][6] * mat_B[6][15] +
                  mat_A[21][7] * mat_B[7][15] +
                  mat_A[21][8] * mat_B[8][15] +
                  mat_A[21][9] * mat_B[9][15] +
                  mat_A[21][10] * mat_B[10][15] +
                  mat_A[21][11] * mat_B[11][15] +
                  mat_A[21][12] * mat_B[12][15] +
                  mat_A[21][13] * mat_B[13][15] +
                  mat_A[21][14] * mat_B[14][15] +
                  mat_A[21][15] * mat_B[15][15] +
                  mat_A[21][16] * mat_B[16][15] +
                  mat_A[21][17] * mat_B[17][15] +
                  mat_A[21][18] * mat_B[18][15] +
                  mat_A[21][19] * mat_B[19][15] +
                  mat_A[21][20] * mat_B[20][15] +
                  mat_A[21][21] * mat_B[21][15] +
                  mat_A[21][22] * mat_B[22][15] +
                  mat_A[21][23] * mat_B[23][15] +
                  mat_A[21][24] * mat_B[24][15] +
                  mat_A[21][25] * mat_B[25][15] +
                  mat_A[21][26] * mat_B[26][15] +
                  mat_A[21][27] * mat_B[27][15] +
                  mat_A[21][28] * mat_B[28][15] +
                  mat_A[21][29] * mat_B[29][15] +
                  mat_A[21][30] * mat_B[30][15] +
                  mat_A[21][31] * mat_B[31][15];
    mat_C[21][16] <= 
                  mat_A[21][0] * mat_B[0][16] +
                  mat_A[21][1] * mat_B[1][16] +
                  mat_A[21][2] * mat_B[2][16] +
                  mat_A[21][3] * mat_B[3][16] +
                  mat_A[21][4] * mat_B[4][16] +
                  mat_A[21][5] * mat_B[5][16] +
                  mat_A[21][6] * mat_B[6][16] +
                  mat_A[21][7] * mat_B[7][16] +
                  mat_A[21][8] * mat_B[8][16] +
                  mat_A[21][9] * mat_B[9][16] +
                  mat_A[21][10] * mat_B[10][16] +
                  mat_A[21][11] * mat_B[11][16] +
                  mat_A[21][12] * mat_B[12][16] +
                  mat_A[21][13] * mat_B[13][16] +
                  mat_A[21][14] * mat_B[14][16] +
                  mat_A[21][15] * mat_B[15][16] +
                  mat_A[21][16] * mat_B[16][16] +
                  mat_A[21][17] * mat_B[17][16] +
                  mat_A[21][18] * mat_B[18][16] +
                  mat_A[21][19] * mat_B[19][16] +
                  mat_A[21][20] * mat_B[20][16] +
                  mat_A[21][21] * mat_B[21][16] +
                  mat_A[21][22] * mat_B[22][16] +
                  mat_A[21][23] * mat_B[23][16] +
                  mat_A[21][24] * mat_B[24][16] +
                  mat_A[21][25] * mat_B[25][16] +
                  mat_A[21][26] * mat_B[26][16] +
                  mat_A[21][27] * mat_B[27][16] +
                  mat_A[21][28] * mat_B[28][16] +
                  mat_A[21][29] * mat_B[29][16] +
                  mat_A[21][30] * mat_B[30][16] +
                  mat_A[21][31] * mat_B[31][16];
    mat_C[21][17] <= 
                  mat_A[21][0] * mat_B[0][17] +
                  mat_A[21][1] * mat_B[1][17] +
                  mat_A[21][2] * mat_B[2][17] +
                  mat_A[21][3] * mat_B[3][17] +
                  mat_A[21][4] * mat_B[4][17] +
                  mat_A[21][5] * mat_B[5][17] +
                  mat_A[21][6] * mat_B[6][17] +
                  mat_A[21][7] * mat_B[7][17] +
                  mat_A[21][8] * mat_B[8][17] +
                  mat_A[21][9] * mat_B[9][17] +
                  mat_A[21][10] * mat_B[10][17] +
                  mat_A[21][11] * mat_B[11][17] +
                  mat_A[21][12] * mat_B[12][17] +
                  mat_A[21][13] * mat_B[13][17] +
                  mat_A[21][14] * mat_B[14][17] +
                  mat_A[21][15] * mat_B[15][17] +
                  mat_A[21][16] * mat_B[16][17] +
                  mat_A[21][17] * mat_B[17][17] +
                  mat_A[21][18] * mat_B[18][17] +
                  mat_A[21][19] * mat_B[19][17] +
                  mat_A[21][20] * mat_B[20][17] +
                  mat_A[21][21] * mat_B[21][17] +
                  mat_A[21][22] * mat_B[22][17] +
                  mat_A[21][23] * mat_B[23][17] +
                  mat_A[21][24] * mat_B[24][17] +
                  mat_A[21][25] * mat_B[25][17] +
                  mat_A[21][26] * mat_B[26][17] +
                  mat_A[21][27] * mat_B[27][17] +
                  mat_A[21][28] * mat_B[28][17] +
                  mat_A[21][29] * mat_B[29][17] +
                  mat_A[21][30] * mat_B[30][17] +
                  mat_A[21][31] * mat_B[31][17];
    mat_C[21][18] <= 
                  mat_A[21][0] * mat_B[0][18] +
                  mat_A[21][1] * mat_B[1][18] +
                  mat_A[21][2] * mat_B[2][18] +
                  mat_A[21][3] * mat_B[3][18] +
                  mat_A[21][4] * mat_B[4][18] +
                  mat_A[21][5] * mat_B[5][18] +
                  mat_A[21][6] * mat_B[6][18] +
                  mat_A[21][7] * mat_B[7][18] +
                  mat_A[21][8] * mat_B[8][18] +
                  mat_A[21][9] * mat_B[9][18] +
                  mat_A[21][10] * mat_B[10][18] +
                  mat_A[21][11] * mat_B[11][18] +
                  mat_A[21][12] * mat_B[12][18] +
                  mat_A[21][13] * mat_B[13][18] +
                  mat_A[21][14] * mat_B[14][18] +
                  mat_A[21][15] * mat_B[15][18] +
                  mat_A[21][16] * mat_B[16][18] +
                  mat_A[21][17] * mat_B[17][18] +
                  mat_A[21][18] * mat_B[18][18] +
                  mat_A[21][19] * mat_B[19][18] +
                  mat_A[21][20] * mat_B[20][18] +
                  mat_A[21][21] * mat_B[21][18] +
                  mat_A[21][22] * mat_B[22][18] +
                  mat_A[21][23] * mat_B[23][18] +
                  mat_A[21][24] * mat_B[24][18] +
                  mat_A[21][25] * mat_B[25][18] +
                  mat_A[21][26] * mat_B[26][18] +
                  mat_A[21][27] * mat_B[27][18] +
                  mat_A[21][28] * mat_B[28][18] +
                  mat_A[21][29] * mat_B[29][18] +
                  mat_A[21][30] * mat_B[30][18] +
                  mat_A[21][31] * mat_B[31][18];
    mat_C[21][19] <= 
                  mat_A[21][0] * mat_B[0][19] +
                  mat_A[21][1] * mat_B[1][19] +
                  mat_A[21][2] * mat_B[2][19] +
                  mat_A[21][3] * mat_B[3][19] +
                  mat_A[21][4] * mat_B[4][19] +
                  mat_A[21][5] * mat_B[5][19] +
                  mat_A[21][6] * mat_B[6][19] +
                  mat_A[21][7] * mat_B[7][19] +
                  mat_A[21][8] * mat_B[8][19] +
                  mat_A[21][9] * mat_B[9][19] +
                  mat_A[21][10] * mat_B[10][19] +
                  mat_A[21][11] * mat_B[11][19] +
                  mat_A[21][12] * mat_B[12][19] +
                  mat_A[21][13] * mat_B[13][19] +
                  mat_A[21][14] * mat_B[14][19] +
                  mat_A[21][15] * mat_B[15][19] +
                  mat_A[21][16] * mat_B[16][19] +
                  mat_A[21][17] * mat_B[17][19] +
                  mat_A[21][18] * mat_B[18][19] +
                  mat_A[21][19] * mat_B[19][19] +
                  mat_A[21][20] * mat_B[20][19] +
                  mat_A[21][21] * mat_B[21][19] +
                  mat_A[21][22] * mat_B[22][19] +
                  mat_A[21][23] * mat_B[23][19] +
                  mat_A[21][24] * mat_B[24][19] +
                  mat_A[21][25] * mat_B[25][19] +
                  mat_A[21][26] * mat_B[26][19] +
                  mat_A[21][27] * mat_B[27][19] +
                  mat_A[21][28] * mat_B[28][19] +
                  mat_A[21][29] * mat_B[29][19] +
                  mat_A[21][30] * mat_B[30][19] +
                  mat_A[21][31] * mat_B[31][19];
    mat_C[21][20] <= 
                  mat_A[21][0] * mat_B[0][20] +
                  mat_A[21][1] * mat_B[1][20] +
                  mat_A[21][2] * mat_B[2][20] +
                  mat_A[21][3] * mat_B[3][20] +
                  mat_A[21][4] * mat_B[4][20] +
                  mat_A[21][5] * mat_B[5][20] +
                  mat_A[21][6] * mat_B[6][20] +
                  mat_A[21][7] * mat_B[7][20] +
                  mat_A[21][8] * mat_B[8][20] +
                  mat_A[21][9] * mat_B[9][20] +
                  mat_A[21][10] * mat_B[10][20] +
                  mat_A[21][11] * mat_B[11][20] +
                  mat_A[21][12] * mat_B[12][20] +
                  mat_A[21][13] * mat_B[13][20] +
                  mat_A[21][14] * mat_B[14][20] +
                  mat_A[21][15] * mat_B[15][20] +
                  mat_A[21][16] * mat_B[16][20] +
                  mat_A[21][17] * mat_B[17][20] +
                  mat_A[21][18] * mat_B[18][20] +
                  mat_A[21][19] * mat_B[19][20] +
                  mat_A[21][20] * mat_B[20][20] +
                  mat_A[21][21] * mat_B[21][20] +
                  mat_A[21][22] * mat_B[22][20] +
                  mat_A[21][23] * mat_B[23][20] +
                  mat_A[21][24] * mat_B[24][20] +
                  mat_A[21][25] * mat_B[25][20] +
                  mat_A[21][26] * mat_B[26][20] +
                  mat_A[21][27] * mat_B[27][20] +
                  mat_A[21][28] * mat_B[28][20] +
                  mat_A[21][29] * mat_B[29][20] +
                  mat_A[21][30] * mat_B[30][20] +
                  mat_A[21][31] * mat_B[31][20];
    mat_C[21][21] <= 
                  mat_A[21][0] * mat_B[0][21] +
                  mat_A[21][1] * mat_B[1][21] +
                  mat_A[21][2] * mat_B[2][21] +
                  mat_A[21][3] * mat_B[3][21] +
                  mat_A[21][4] * mat_B[4][21] +
                  mat_A[21][5] * mat_B[5][21] +
                  mat_A[21][6] * mat_B[6][21] +
                  mat_A[21][7] * mat_B[7][21] +
                  mat_A[21][8] * mat_B[8][21] +
                  mat_A[21][9] * mat_B[9][21] +
                  mat_A[21][10] * mat_B[10][21] +
                  mat_A[21][11] * mat_B[11][21] +
                  mat_A[21][12] * mat_B[12][21] +
                  mat_A[21][13] * mat_B[13][21] +
                  mat_A[21][14] * mat_B[14][21] +
                  mat_A[21][15] * mat_B[15][21] +
                  mat_A[21][16] * mat_B[16][21] +
                  mat_A[21][17] * mat_B[17][21] +
                  mat_A[21][18] * mat_B[18][21] +
                  mat_A[21][19] * mat_B[19][21] +
                  mat_A[21][20] * mat_B[20][21] +
                  mat_A[21][21] * mat_B[21][21] +
                  mat_A[21][22] * mat_B[22][21] +
                  mat_A[21][23] * mat_B[23][21] +
                  mat_A[21][24] * mat_B[24][21] +
                  mat_A[21][25] * mat_B[25][21] +
                  mat_A[21][26] * mat_B[26][21] +
                  mat_A[21][27] * mat_B[27][21] +
                  mat_A[21][28] * mat_B[28][21] +
                  mat_A[21][29] * mat_B[29][21] +
                  mat_A[21][30] * mat_B[30][21] +
                  mat_A[21][31] * mat_B[31][21];
    mat_C[21][22] <= 
                  mat_A[21][0] * mat_B[0][22] +
                  mat_A[21][1] * mat_B[1][22] +
                  mat_A[21][2] * mat_B[2][22] +
                  mat_A[21][3] * mat_B[3][22] +
                  mat_A[21][4] * mat_B[4][22] +
                  mat_A[21][5] * mat_B[5][22] +
                  mat_A[21][6] * mat_B[6][22] +
                  mat_A[21][7] * mat_B[7][22] +
                  mat_A[21][8] * mat_B[8][22] +
                  mat_A[21][9] * mat_B[9][22] +
                  mat_A[21][10] * mat_B[10][22] +
                  mat_A[21][11] * mat_B[11][22] +
                  mat_A[21][12] * mat_B[12][22] +
                  mat_A[21][13] * mat_B[13][22] +
                  mat_A[21][14] * mat_B[14][22] +
                  mat_A[21][15] * mat_B[15][22] +
                  mat_A[21][16] * mat_B[16][22] +
                  mat_A[21][17] * mat_B[17][22] +
                  mat_A[21][18] * mat_B[18][22] +
                  mat_A[21][19] * mat_B[19][22] +
                  mat_A[21][20] * mat_B[20][22] +
                  mat_A[21][21] * mat_B[21][22] +
                  mat_A[21][22] * mat_B[22][22] +
                  mat_A[21][23] * mat_B[23][22] +
                  mat_A[21][24] * mat_B[24][22] +
                  mat_A[21][25] * mat_B[25][22] +
                  mat_A[21][26] * mat_B[26][22] +
                  mat_A[21][27] * mat_B[27][22] +
                  mat_A[21][28] * mat_B[28][22] +
                  mat_A[21][29] * mat_B[29][22] +
                  mat_A[21][30] * mat_B[30][22] +
                  mat_A[21][31] * mat_B[31][22];
    mat_C[21][23] <= 
                  mat_A[21][0] * mat_B[0][23] +
                  mat_A[21][1] * mat_B[1][23] +
                  mat_A[21][2] * mat_B[2][23] +
                  mat_A[21][3] * mat_B[3][23] +
                  mat_A[21][4] * mat_B[4][23] +
                  mat_A[21][5] * mat_B[5][23] +
                  mat_A[21][6] * mat_B[6][23] +
                  mat_A[21][7] * mat_B[7][23] +
                  mat_A[21][8] * mat_B[8][23] +
                  mat_A[21][9] * mat_B[9][23] +
                  mat_A[21][10] * mat_B[10][23] +
                  mat_A[21][11] * mat_B[11][23] +
                  mat_A[21][12] * mat_B[12][23] +
                  mat_A[21][13] * mat_B[13][23] +
                  mat_A[21][14] * mat_B[14][23] +
                  mat_A[21][15] * mat_B[15][23] +
                  mat_A[21][16] * mat_B[16][23] +
                  mat_A[21][17] * mat_B[17][23] +
                  mat_A[21][18] * mat_B[18][23] +
                  mat_A[21][19] * mat_B[19][23] +
                  mat_A[21][20] * mat_B[20][23] +
                  mat_A[21][21] * mat_B[21][23] +
                  mat_A[21][22] * mat_B[22][23] +
                  mat_A[21][23] * mat_B[23][23] +
                  mat_A[21][24] * mat_B[24][23] +
                  mat_A[21][25] * mat_B[25][23] +
                  mat_A[21][26] * mat_B[26][23] +
                  mat_A[21][27] * mat_B[27][23] +
                  mat_A[21][28] * mat_B[28][23] +
                  mat_A[21][29] * mat_B[29][23] +
                  mat_A[21][30] * mat_B[30][23] +
                  mat_A[21][31] * mat_B[31][23];
    mat_C[21][24] <= 
                  mat_A[21][0] * mat_B[0][24] +
                  mat_A[21][1] * mat_B[1][24] +
                  mat_A[21][2] * mat_B[2][24] +
                  mat_A[21][3] * mat_B[3][24] +
                  mat_A[21][4] * mat_B[4][24] +
                  mat_A[21][5] * mat_B[5][24] +
                  mat_A[21][6] * mat_B[6][24] +
                  mat_A[21][7] * mat_B[7][24] +
                  mat_A[21][8] * mat_B[8][24] +
                  mat_A[21][9] * mat_B[9][24] +
                  mat_A[21][10] * mat_B[10][24] +
                  mat_A[21][11] * mat_B[11][24] +
                  mat_A[21][12] * mat_B[12][24] +
                  mat_A[21][13] * mat_B[13][24] +
                  mat_A[21][14] * mat_B[14][24] +
                  mat_A[21][15] * mat_B[15][24] +
                  mat_A[21][16] * mat_B[16][24] +
                  mat_A[21][17] * mat_B[17][24] +
                  mat_A[21][18] * mat_B[18][24] +
                  mat_A[21][19] * mat_B[19][24] +
                  mat_A[21][20] * mat_B[20][24] +
                  mat_A[21][21] * mat_B[21][24] +
                  mat_A[21][22] * mat_B[22][24] +
                  mat_A[21][23] * mat_B[23][24] +
                  mat_A[21][24] * mat_B[24][24] +
                  mat_A[21][25] * mat_B[25][24] +
                  mat_A[21][26] * mat_B[26][24] +
                  mat_A[21][27] * mat_B[27][24] +
                  mat_A[21][28] * mat_B[28][24] +
                  mat_A[21][29] * mat_B[29][24] +
                  mat_A[21][30] * mat_B[30][24] +
                  mat_A[21][31] * mat_B[31][24];
    mat_C[21][25] <= 
                  mat_A[21][0] * mat_B[0][25] +
                  mat_A[21][1] * mat_B[1][25] +
                  mat_A[21][2] * mat_B[2][25] +
                  mat_A[21][3] * mat_B[3][25] +
                  mat_A[21][4] * mat_B[4][25] +
                  mat_A[21][5] * mat_B[5][25] +
                  mat_A[21][6] * mat_B[6][25] +
                  mat_A[21][7] * mat_B[7][25] +
                  mat_A[21][8] * mat_B[8][25] +
                  mat_A[21][9] * mat_B[9][25] +
                  mat_A[21][10] * mat_B[10][25] +
                  mat_A[21][11] * mat_B[11][25] +
                  mat_A[21][12] * mat_B[12][25] +
                  mat_A[21][13] * mat_B[13][25] +
                  mat_A[21][14] * mat_B[14][25] +
                  mat_A[21][15] * mat_B[15][25] +
                  mat_A[21][16] * mat_B[16][25] +
                  mat_A[21][17] * mat_B[17][25] +
                  mat_A[21][18] * mat_B[18][25] +
                  mat_A[21][19] * mat_B[19][25] +
                  mat_A[21][20] * mat_B[20][25] +
                  mat_A[21][21] * mat_B[21][25] +
                  mat_A[21][22] * mat_B[22][25] +
                  mat_A[21][23] * mat_B[23][25] +
                  mat_A[21][24] * mat_B[24][25] +
                  mat_A[21][25] * mat_B[25][25] +
                  mat_A[21][26] * mat_B[26][25] +
                  mat_A[21][27] * mat_B[27][25] +
                  mat_A[21][28] * mat_B[28][25] +
                  mat_A[21][29] * mat_B[29][25] +
                  mat_A[21][30] * mat_B[30][25] +
                  mat_A[21][31] * mat_B[31][25];
    mat_C[21][26] <= 
                  mat_A[21][0] * mat_B[0][26] +
                  mat_A[21][1] * mat_B[1][26] +
                  mat_A[21][2] * mat_B[2][26] +
                  mat_A[21][3] * mat_B[3][26] +
                  mat_A[21][4] * mat_B[4][26] +
                  mat_A[21][5] * mat_B[5][26] +
                  mat_A[21][6] * mat_B[6][26] +
                  mat_A[21][7] * mat_B[7][26] +
                  mat_A[21][8] * mat_B[8][26] +
                  mat_A[21][9] * mat_B[9][26] +
                  mat_A[21][10] * mat_B[10][26] +
                  mat_A[21][11] * mat_B[11][26] +
                  mat_A[21][12] * mat_B[12][26] +
                  mat_A[21][13] * mat_B[13][26] +
                  mat_A[21][14] * mat_B[14][26] +
                  mat_A[21][15] * mat_B[15][26] +
                  mat_A[21][16] * mat_B[16][26] +
                  mat_A[21][17] * mat_B[17][26] +
                  mat_A[21][18] * mat_B[18][26] +
                  mat_A[21][19] * mat_B[19][26] +
                  mat_A[21][20] * mat_B[20][26] +
                  mat_A[21][21] * mat_B[21][26] +
                  mat_A[21][22] * mat_B[22][26] +
                  mat_A[21][23] * mat_B[23][26] +
                  mat_A[21][24] * mat_B[24][26] +
                  mat_A[21][25] * mat_B[25][26] +
                  mat_A[21][26] * mat_B[26][26] +
                  mat_A[21][27] * mat_B[27][26] +
                  mat_A[21][28] * mat_B[28][26] +
                  mat_A[21][29] * mat_B[29][26] +
                  mat_A[21][30] * mat_B[30][26] +
                  mat_A[21][31] * mat_B[31][26];
    mat_C[21][27] <= 
                  mat_A[21][0] * mat_B[0][27] +
                  mat_A[21][1] * mat_B[1][27] +
                  mat_A[21][2] * mat_B[2][27] +
                  mat_A[21][3] * mat_B[3][27] +
                  mat_A[21][4] * mat_B[4][27] +
                  mat_A[21][5] * mat_B[5][27] +
                  mat_A[21][6] * mat_B[6][27] +
                  mat_A[21][7] * mat_B[7][27] +
                  mat_A[21][8] * mat_B[8][27] +
                  mat_A[21][9] * mat_B[9][27] +
                  mat_A[21][10] * mat_B[10][27] +
                  mat_A[21][11] * mat_B[11][27] +
                  mat_A[21][12] * mat_B[12][27] +
                  mat_A[21][13] * mat_B[13][27] +
                  mat_A[21][14] * mat_B[14][27] +
                  mat_A[21][15] * mat_B[15][27] +
                  mat_A[21][16] * mat_B[16][27] +
                  mat_A[21][17] * mat_B[17][27] +
                  mat_A[21][18] * mat_B[18][27] +
                  mat_A[21][19] * mat_B[19][27] +
                  mat_A[21][20] * mat_B[20][27] +
                  mat_A[21][21] * mat_B[21][27] +
                  mat_A[21][22] * mat_B[22][27] +
                  mat_A[21][23] * mat_B[23][27] +
                  mat_A[21][24] * mat_B[24][27] +
                  mat_A[21][25] * mat_B[25][27] +
                  mat_A[21][26] * mat_B[26][27] +
                  mat_A[21][27] * mat_B[27][27] +
                  mat_A[21][28] * mat_B[28][27] +
                  mat_A[21][29] * mat_B[29][27] +
                  mat_A[21][30] * mat_B[30][27] +
                  mat_A[21][31] * mat_B[31][27];
    mat_C[21][28] <= 
                  mat_A[21][0] * mat_B[0][28] +
                  mat_A[21][1] * mat_B[1][28] +
                  mat_A[21][2] * mat_B[2][28] +
                  mat_A[21][3] * mat_B[3][28] +
                  mat_A[21][4] * mat_B[4][28] +
                  mat_A[21][5] * mat_B[5][28] +
                  mat_A[21][6] * mat_B[6][28] +
                  mat_A[21][7] * mat_B[7][28] +
                  mat_A[21][8] * mat_B[8][28] +
                  mat_A[21][9] * mat_B[9][28] +
                  mat_A[21][10] * mat_B[10][28] +
                  mat_A[21][11] * mat_B[11][28] +
                  mat_A[21][12] * mat_B[12][28] +
                  mat_A[21][13] * mat_B[13][28] +
                  mat_A[21][14] * mat_B[14][28] +
                  mat_A[21][15] * mat_B[15][28] +
                  mat_A[21][16] * mat_B[16][28] +
                  mat_A[21][17] * mat_B[17][28] +
                  mat_A[21][18] * mat_B[18][28] +
                  mat_A[21][19] * mat_B[19][28] +
                  mat_A[21][20] * mat_B[20][28] +
                  mat_A[21][21] * mat_B[21][28] +
                  mat_A[21][22] * mat_B[22][28] +
                  mat_A[21][23] * mat_B[23][28] +
                  mat_A[21][24] * mat_B[24][28] +
                  mat_A[21][25] * mat_B[25][28] +
                  mat_A[21][26] * mat_B[26][28] +
                  mat_A[21][27] * mat_B[27][28] +
                  mat_A[21][28] * mat_B[28][28] +
                  mat_A[21][29] * mat_B[29][28] +
                  mat_A[21][30] * mat_B[30][28] +
                  mat_A[21][31] * mat_B[31][28];
    mat_C[21][29] <= 
                  mat_A[21][0] * mat_B[0][29] +
                  mat_A[21][1] * mat_B[1][29] +
                  mat_A[21][2] * mat_B[2][29] +
                  mat_A[21][3] * mat_B[3][29] +
                  mat_A[21][4] * mat_B[4][29] +
                  mat_A[21][5] * mat_B[5][29] +
                  mat_A[21][6] * mat_B[6][29] +
                  mat_A[21][7] * mat_B[7][29] +
                  mat_A[21][8] * mat_B[8][29] +
                  mat_A[21][9] * mat_B[9][29] +
                  mat_A[21][10] * mat_B[10][29] +
                  mat_A[21][11] * mat_B[11][29] +
                  mat_A[21][12] * mat_B[12][29] +
                  mat_A[21][13] * mat_B[13][29] +
                  mat_A[21][14] * mat_B[14][29] +
                  mat_A[21][15] * mat_B[15][29] +
                  mat_A[21][16] * mat_B[16][29] +
                  mat_A[21][17] * mat_B[17][29] +
                  mat_A[21][18] * mat_B[18][29] +
                  mat_A[21][19] * mat_B[19][29] +
                  mat_A[21][20] * mat_B[20][29] +
                  mat_A[21][21] * mat_B[21][29] +
                  mat_A[21][22] * mat_B[22][29] +
                  mat_A[21][23] * mat_B[23][29] +
                  mat_A[21][24] * mat_B[24][29] +
                  mat_A[21][25] * mat_B[25][29] +
                  mat_A[21][26] * mat_B[26][29] +
                  mat_A[21][27] * mat_B[27][29] +
                  mat_A[21][28] * mat_B[28][29] +
                  mat_A[21][29] * mat_B[29][29] +
                  mat_A[21][30] * mat_B[30][29] +
                  mat_A[21][31] * mat_B[31][29];
    mat_C[21][30] <= 
                  mat_A[21][0] * mat_B[0][30] +
                  mat_A[21][1] * mat_B[1][30] +
                  mat_A[21][2] * mat_B[2][30] +
                  mat_A[21][3] * mat_B[3][30] +
                  mat_A[21][4] * mat_B[4][30] +
                  mat_A[21][5] * mat_B[5][30] +
                  mat_A[21][6] * mat_B[6][30] +
                  mat_A[21][7] * mat_B[7][30] +
                  mat_A[21][8] * mat_B[8][30] +
                  mat_A[21][9] * mat_B[9][30] +
                  mat_A[21][10] * mat_B[10][30] +
                  mat_A[21][11] * mat_B[11][30] +
                  mat_A[21][12] * mat_B[12][30] +
                  mat_A[21][13] * mat_B[13][30] +
                  mat_A[21][14] * mat_B[14][30] +
                  mat_A[21][15] * mat_B[15][30] +
                  mat_A[21][16] * mat_B[16][30] +
                  mat_A[21][17] * mat_B[17][30] +
                  mat_A[21][18] * mat_B[18][30] +
                  mat_A[21][19] * mat_B[19][30] +
                  mat_A[21][20] * mat_B[20][30] +
                  mat_A[21][21] * mat_B[21][30] +
                  mat_A[21][22] * mat_B[22][30] +
                  mat_A[21][23] * mat_B[23][30] +
                  mat_A[21][24] * mat_B[24][30] +
                  mat_A[21][25] * mat_B[25][30] +
                  mat_A[21][26] * mat_B[26][30] +
                  mat_A[21][27] * mat_B[27][30] +
                  mat_A[21][28] * mat_B[28][30] +
                  mat_A[21][29] * mat_B[29][30] +
                  mat_A[21][30] * mat_B[30][30] +
                  mat_A[21][31] * mat_B[31][30];
    mat_C[21][31] <= 
                  mat_A[21][0] * mat_B[0][31] +
                  mat_A[21][1] * mat_B[1][31] +
                  mat_A[21][2] * mat_B[2][31] +
                  mat_A[21][3] * mat_B[3][31] +
                  mat_A[21][4] * mat_B[4][31] +
                  mat_A[21][5] * mat_B[5][31] +
                  mat_A[21][6] * mat_B[6][31] +
                  mat_A[21][7] * mat_B[7][31] +
                  mat_A[21][8] * mat_B[8][31] +
                  mat_A[21][9] * mat_B[9][31] +
                  mat_A[21][10] * mat_B[10][31] +
                  mat_A[21][11] * mat_B[11][31] +
                  mat_A[21][12] * mat_B[12][31] +
                  mat_A[21][13] * mat_B[13][31] +
                  mat_A[21][14] * mat_B[14][31] +
                  mat_A[21][15] * mat_B[15][31] +
                  mat_A[21][16] * mat_B[16][31] +
                  mat_A[21][17] * mat_B[17][31] +
                  mat_A[21][18] * mat_B[18][31] +
                  mat_A[21][19] * mat_B[19][31] +
                  mat_A[21][20] * mat_B[20][31] +
                  mat_A[21][21] * mat_B[21][31] +
                  mat_A[21][22] * mat_B[22][31] +
                  mat_A[21][23] * mat_B[23][31] +
                  mat_A[21][24] * mat_B[24][31] +
                  mat_A[21][25] * mat_B[25][31] +
                  mat_A[21][26] * mat_B[26][31] +
                  mat_A[21][27] * mat_B[27][31] +
                  mat_A[21][28] * mat_B[28][31] +
                  mat_A[21][29] * mat_B[29][31] +
                  mat_A[21][30] * mat_B[30][31] +
                  mat_A[21][31] * mat_B[31][31];
    mat_C[22][0] <= 
                  mat_A[22][0] * mat_B[0][0] +
                  mat_A[22][1] * mat_B[1][0] +
                  mat_A[22][2] * mat_B[2][0] +
                  mat_A[22][3] * mat_B[3][0] +
                  mat_A[22][4] * mat_B[4][0] +
                  mat_A[22][5] * mat_B[5][0] +
                  mat_A[22][6] * mat_B[6][0] +
                  mat_A[22][7] * mat_B[7][0] +
                  mat_A[22][8] * mat_B[8][0] +
                  mat_A[22][9] * mat_B[9][0] +
                  mat_A[22][10] * mat_B[10][0] +
                  mat_A[22][11] * mat_B[11][0] +
                  mat_A[22][12] * mat_B[12][0] +
                  mat_A[22][13] * mat_B[13][0] +
                  mat_A[22][14] * mat_B[14][0] +
                  mat_A[22][15] * mat_B[15][0] +
                  mat_A[22][16] * mat_B[16][0] +
                  mat_A[22][17] * mat_B[17][0] +
                  mat_A[22][18] * mat_B[18][0] +
                  mat_A[22][19] * mat_B[19][0] +
                  mat_A[22][20] * mat_B[20][0] +
                  mat_A[22][21] * mat_B[21][0] +
                  mat_A[22][22] * mat_B[22][0] +
                  mat_A[22][23] * mat_B[23][0] +
                  mat_A[22][24] * mat_B[24][0] +
                  mat_A[22][25] * mat_B[25][0] +
                  mat_A[22][26] * mat_B[26][0] +
                  mat_A[22][27] * mat_B[27][0] +
                  mat_A[22][28] * mat_B[28][0] +
                  mat_A[22][29] * mat_B[29][0] +
                  mat_A[22][30] * mat_B[30][0] +
                  mat_A[22][31] * mat_B[31][0];
    mat_C[22][1] <= 
                  mat_A[22][0] * mat_B[0][1] +
                  mat_A[22][1] * mat_B[1][1] +
                  mat_A[22][2] * mat_B[2][1] +
                  mat_A[22][3] * mat_B[3][1] +
                  mat_A[22][4] * mat_B[4][1] +
                  mat_A[22][5] * mat_B[5][1] +
                  mat_A[22][6] * mat_B[6][1] +
                  mat_A[22][7] * mat_B[7][1] +
                  mat_A[22][8] * mat_B[8][1] +
                  mat_A[22][9] * mat_B[9][1] +
                  mat_A[22][10] * mat_B[10][1] +
                  mat_A[22][11] * mat_B[11][1] +
                  mat_A[22][12] * mat_B[12][1] +
                  mat_A[22][13] * mat_B[13][1] +
                  mat_A[22][14] * mat_B[14][1] +
                  mat_A[22][15] * mat_B[15][1] +
                  mat_A[22][16] * mat_B[16][1] +
                  mat_A[22][17] * mat_B[17][1] +
                  mat_A[22][18] * mat_B[18][1] +
                  mat_A[22][19] * mat_B[19][1] +
                  mat_A[22][20] * mat_B[20][1] +
                  mat_A[22][21] * mat_B[21][1] +
                  mat_A[22][22] * mat_B[22][1] +
                  mat_A[22][23] * mat_B[23][1] +
                  mat_A[22][24] * mat_B[24][1] +
                  mat_A[22][25] * mat_B[25][1] +
                  mat_A[22][26] * mat_B[26][1] +
                  mat_A[22][27] * mat_B[27][1] +
                  mat_A[22][28] * mat_B[28][1] +
                  mat_A[22][29] * mat_B[29][1] +
                  mat_A[22][30] * mat_B[30][1] +
                  mat_A[22][31] * mat_B[31][1];
    mat_C[22][2] <= 
                  mat_A[22][0] * mat_B[0][2] +
                  mat_A[22][1] * mat_B[1][2] +
                  mat_A[22][2] * mat_B[2][2] +
                  mat_A[22][3] * mat_B[3][2] +
                  mat_A[22][4] * mat_B[4][2] +
                  mat_A[22][5] * mat_B[5][2] +
                  mat_A[22][6] * mat_B[6][2] +
                  mat_A[22][7] * mat_B[7][2] +
                  mat_A[22][8] * mat_B[8][2] +
                  mat_A[22][9] * mat_B[9][2] +
                  mat_A[22][10] * mat_B[10][2] +
                  mat_A[22][11] * mat_B[11][2] +
                  mat_A[22][12] * mat_B[12][2] +
                  mat_A[22][13] * mat_B[13][2] +
                  mat_A[22][14] * mat_B[14][2] +
                  mat_A[22][15] * mat_B[15][2] +
                  mat_A[22][16] * mat_B[16][2] +
                  mat_A[22][17] * mat_B[17][2] +
                  mat_A[22][18] * mat_B[18][2] +
                  mat_A[22][19] * mat_B[19][2] +
                  mat_A[22][20] * mat_B[20][2] +
                  mat_A[22][21] * mat_B[21][2] +
                  mat_A[22][22] * mat_B[22][2] +
                  mat_A[22][23] * mat_B[23][2] +
                  mat_A[22][24] * mat_B[24][2] +
                  mat_A[22][25] * mat_B[25][2] +
                  mat_A[22][26] * mat_B[26][2] +
                  mat_A[22][27] * mat_B[27][2] +
                  mat_A[22][28] * mat_B[28][2] +
                  mat_A[22][29] * mat_B[29][2] +
                  mat_A[22][30] * mat_B[30][2] +
                  mat_A[22][31] * mat_B[31][2];
    mat_C[22][3] <= 
                  mat_A[22][0] * mat_B[0][3] +
                  mat_A[22][1] * mat_B[1][3] +
                  mat_A[22][2] * mat_B[2][3] +
                  mat_A[22][3] * mat_B[3][3] +
                  mat_A[22][4] * mat_B[4][3] +
                  mat_A[22][5] * mat_B[5][3] +
                  mat_A[22][6] * mat_B[6][3] +
                  mat_A[22][7] * mat_B[7][3] +
                  mat_A[22][8] * mat_B[8][3] +
                  mat_A[22][9] * mat_B[9][3] +
                  mat_A[22][10] * mat_B[10][3] +
                  mat_A[22][11] * mat_B[11][3] +
                  mat_A[22][12] * mat_B[12][3] +
                  mat_A[22][13] * mat_B[13][3] +
                  mat_A[22][14] * mat_B[14][3] +
                  mat_A[22][15] * mat_B[15][3] +
                  mat_A[22][16] * mat_B[16][3] +
                  mat_A[22][17] * mat_B[17][3] +
                  mat_A[22][18] * mat_B[18][3] +
                  mat_A[22][19] * mat_B[19][3] +
                  mat_A[22][20] * mat_B[20][3] +
                  mat_A[22][21] * mat_B[21][3] +
                  mat_A[22][22] * mat_B[22][3] +
                  mat_A[22][23] * mat_B[23][3] +
                  mat_A[22][24] * mat_B[24][3] +
                  mat_A[22][25] * mat_B[25][3] +
                  mat_A[22][26] * mat_B[26][3] +
                  mat_A[22][27] * mat_B[27][3] +
                  mat_A[22][28] * mat_B[28][3] +
                  mat_A[22][29] * mat_B[29][3] +
                  mat_A[22][30] * mat_B[30][3] +
                  mat_A[22][31] * mat_B[31][3];
    mat_C[22][4] <= 
                  mat_A[22][0] * mat_B[0][4] +
                  mat_A[22][1] * mat_B[1][4] +
                  mat_A[22][2] * mat_B[2][4] +
                  mat_A[22][3] * mat_B[3][4] +
                  mat_A[22][4] * mat_B[4][4] +
                  mat_A[22][5] * mat_B[5][4] +
                  mat_A[22][6] * mat_B[6][4] +
                  mat_A[22][7] * mat_B[7][4] +
                  mat_A[22][8] * mat_B[8][4] +
                  mat_A[22][9] * mat_B[9][4] +
                  mat_A[22][10] * mat_B[10][4] +
                  mat_A[22][11] * mat_B[11][4] +
                  mat_A[22][12] * mat_B[12][4] +
                  mat_A[22][13] * mat_B[13][4] +
                  mat_A[22][14] * mat_B[14][4] +
                  mat_A[22][15] * mat_B[15][4] +
                  mat_A[22][16] * mat_B[16][4] +
                  mat_A[22][17] * mat_B[17][4] +
                  mat_A[22][18] * mat_B[18][4] +
                  mat_A[22][19] * mat_B[19][4] +
                  mat_A[22][20] * mat_B[20][4] +
                  mat_A[22][21] * mat_B[21][4] +
                  mat_A[22][22] * mat_B[22][4] +
                  mat_A[22][23] * mat_B[23][4] +
                  mat_A[22][24] * mat_B[24][4] +
                  mat_A[22][25] * mat_B[25][4] +
                  mat_A[22][26] * mat_B[26][4] +
                  mat_A[22][27] * mat_B[27][4] +
                  mat_A[22][28] * mat_B[28][4] +
                  mat_A[22][29] * mat_B[29][4] +
                  mat_A[22][30] * mat_B[30][4] +
                  mat_A[22][31] * mat_B[31][4];
    mat_C[22][5] <= 
                  mat_A[22][0] * mat_B[0][5] +
                  mat_A[22][1] * mat_B[1][5] +
                  mat_A[22][2] * mat_B[2][5] +
                  mat_A[22][3] * mat_B[3][5] +
                  mat_A[22][4] * mat_B[4][5] +
                  mat_A[22][5] * mat_B[5][5] +
                  mat_A[22][6] * mat_B[6][5] +
                  mat_A[22][7] * mat_B[7][5] +
                  mat_A[22][8] * mat_B[8][5] +
                  mat_A[22][9] * mat_B[9][5] +
                  mat_A[22][10] * mat_B[10][5] +
                  mat_A[22][11] * mat_B[11][5] +
                  mat_A[22][12] * mat_B[12][5] +
                  mat_A[22][13] * mat_B[13][5] +
                  mat_A[22][14] * mat_B[14][5] +
                  mat_A[22][15] * mat_B[15][5] +
                  mat_A[22][16] * mat_B[16][5] +
                  mat_A[22][17] * mat_B[17][5] +
                  mat_A[22][18] * mat_B[18][5] +
                  mat_A[22][19] * mat_B[19][5] +
                  mat_A[22][20] * mat_B[20][5] +
                  mat_A[22][21] * mat_B[21][5] +
                  mat_A[22][22] * mat_B[22][5] +
                  mat_A[22][23] * mat_B[23][5] +
                  mat_A[22][24] * mat_B[24][5] +
                  mat_A[22][25] * mat_B[25][5] +
                  mat_A[22][26] * mat_B[26][5] +
                  mat_A[22][27] * mat_B[27][5] +
                  mat_A[22][28] * mat_B[28][5] +
                  mat_A[22][29] * mat_B[29][5] +
                  mat_A[22][30] * mat_B[30][5] +
                  mat_A[22][31] * mat_B[31][5];
    mat_C[22][6] <= 
                  mat_A[22][0] * mat_B[0][6] +
                  mat_A[22][1] * mat_B[1][6] +
                  mat_A[22][2] * mat_B[2][6] +
                  mat_A[22][3] * mat_B[3][6] +
                  mat_A[22][4] * mat_B[4][6] +
                  mat_A[22][5] * mat_B[5][6] +
                  mat_A[22][6] * mat_B[6][6] +
                  mat_A[22][7] * mat_B[7][6] +
                  mat_A[22][8] * mat_B[8][6] +
                  mat_A[22][9] * mat_B[9][6] +
                  mat_A[22][10] * mat_B[10][6] +
                  mat_A[22][11] * mat_B[11][6] +
                  mat_A[22][12] * mat_B[12][6] +
                  mat_A[22][13] * mat_B[13][6] +
                  mat_A[22][14] * mat_B[14][6] +
                  mat_A[22][15] * mat_B[15][6] +
                  mat_A[22][16] * mat_B[16][6] +
                  mat_A[22][17] * mat_B[17][6] +
                  mat_A[22][18] * mat_B[18][6] +
                  mat_A[22][19] * mat_B[19][6] +
                  mat_A[22][20] * mat_B[20][6] +
                  mat_A[22][21] * mat_B[21][6] +
                  mat_A[22][22] * mat_B[22][6] +
                  mat_A[22][23] * mat_B[23][6] +
                  mat_A[22][24] * mat_B[24][6] +
                  mat_A[22][25] * mat_B[25][6] +
                  mat_A[22][26] * mat_B[26][6] +
                  mat_A[22][27] * mat_B[27][6] +
                  mat_A[22][28] * mat_B[28][6] +
                  mat_A[22][29] * mat_B[29][6] +
                  mat_A[22][30] * mat_B[30][6] +
                  mat_A[22][31] * mat_B[31][6];
    mat_C[22][7] <= 
                  mat_A[22][0] * mat_B[0][7] +
                  mat_A[22][1] * mat_B[1][7] +
                  mat_A[22][2] * mat_B[2][7] +
                  mat_A[22][3] * mat_B[3][7] +
                  mat_A[22][4] * mat_B[4][7] +
                  mat_A[22][5] * mat_B[5][7] +
                  mat_A[22][6] * mat_B[6][7] +
                  mat_A[22][7] * mat_B[7][7] +
                  mat_A[22][8] * mat_B[8][7] +
                  mat_A[22][9] * mat_B[9][7] +
                  mat_A[22][10] * mat_B[10][7] +
                  mat_A[22][11] * mat_B[11][7] +
                  mat_A[22][12] * mat_B[12][7] +
                  mat_A[22][13] * mat_B[13][7] +
                  mat_A[22][14] * mat_B[14][7] +
                  mat_A[22][15] * mat_B[15][7] +
                  mat_A[22][16] * mat_B[16][7] +
                  mat_A[22][17] * mat_B[17][7] +
                  mat_A[22][18] * mat_B[18][7] +
                  mat_A[22][19] * mat_B[19][7] +
                  mat_A[22][20] * mat_B[20][7] +
                  mat_A[22][21] * mat_B[21][7] +
                  mat_A[22][22] * mat_B[22][7] +
                  mat_A[22][23] * mat_B[23][7] +
                  mat_A[22][24] * mat_B[24][7] +
                  mat_A[22][25] * mat_B[25][7] +
                  mat_A[22][26] * mat_B[26][7] +
                  mat_A[22][27] * mat_B[27][7] +
                  mat_A[22][28] * mat_B[28][7] +
                  mat_A[22][29] * mat_B[29][7] +
                  mat_A[22][30] * mat_B[30][7] +
                  mat_A[22][31] * mat_B[31][7];
    mat_C[22][8] <= 
                  mat_A[22][0] * mat_B[0][8] +
                  mat_A[22][1] * mat_B[1][8] +
                  mat_A[22][2] * mat_B[2][8] +
                  mat_A[22][3] * mat_B[3][8] +
                  mat_A[22][4] * mat_B[4][8] +
                  mat_A[22][5] * mat_B[5][8] +
                  mat_A[22][6] * mat_B[6][8] +
                  mat_A[22][7] * mat_B[7][8] +
                  mat_A[22][8] * mat_B[8][8] +
                  mat_A[22][9] * mat_B[9][8] +
                  mat_A[22][10] * mat_B[10][8] +
                  mat_A[22][11] * mat_B[11][8] +
                  mat_A[22][12] * mat_B[12][8] +
                  mat_A[22][13] * mat_B[13][8] +
                  mat_A[22][14] * mat_B[14][8] +
                  mat_A[22][15] * mat_B[15][8] +
                  mat_A[22][16] * mat_B[16][8] +
                  mat_A[22][17] * mat_B[17][8] +
                  mat_A[22][18] * mat_B[18][8] +
                  mat_A[22][19] * mat_B[19][8] +
                  mat_A[22][20] * mat_B[20][8] +
                  mat_A[22][21] * mat_B[21][8] +
                  mat_A[22][22] * mat_B[22][8] +
                  mat_A[22][23] * mat_B[23][8] +
                  mat_A[22][24] * mat_B[24][8] +
                  mat_A[22][25] * mat_B[25][8] +
                  mat_A[22][26] * mat_B[26][8] +
                  mat_A[22][27] * mat_B[27][8] +
                  mat_A[22][28] * mat_B[28][8] +
                  mat_A[22][29] * mat_B[29][8] +
                  mat_A[22][30] * mat_B[30][8] +
                  mat_A[22][31] * mat_B[31][8];
    mat_C[22][9] <= 
                  mat_A[22][0] * mat_B[0][9] +
                  mat_A[22][1] * mat_B[1][9] +
                  mat_A[22][2] * mat_B[2][9] +
                  mat_A[22][3] * mat_B[3][9] +
                  mat_A[22][4] * mat_B[4][9] +
                  mat_A[22][5] * mat_B[5][9] +
                  mat_A[22][6] * mat_B[6][9] +
                  mat_A[22][7] * mat_B[7][9] +
                  mat_A[22][8] * mat_B[8][9] +
                  mat_A[22][9] * mat_B[9][9] +
                  mat_A[22][10] * mat_B[10][9] +
                  mat_A[22][11] * mat_B[11][9] +
                  mat_A[22][12] * mat_B[12][9] +
                  mat_A[22][13] * mat_B[13][9] +
                  mat_A[22][14] * mat_B[14][9] +
                  mat_A[22][15] * mat_B[15][9] +
                  mat_A[22][16] * mat_B[16][9] +
                  mat_A[22][17] * mat_B[17][9] +
                  mat_A[22][18] * mat_B[18][9] +
                  mat_A[22][19] * mat_B[19][9] +
                  mat_A[22][20] * mat_B[20][9] +
                  mat_A[22][21] * mat_B[21][9] +
                  mat_A[22][22] * mat_B[22][9] +
                  mat_A[22][23] * mat_B[23][9] +
                  mat_A[22][24] * mat_B[24][9] +
                  mat_A[22][25] * mat_B[25][9] +
                  mat_A[22][26] * mat_B[26][9] +
                  mat_A[22][27] * mat_B[27][9] +
                  mat_A[22][28] * mat_B[28][9] +
                  mat_A[22][29] * mat_B[29][9] +
                  mat_A[22][30] * mat_B[30][9] +
                  mat_A[22][31] * mat_B[31][9];
    mat_C[22][10] <= 
                  mat_A[22][0] * mat_B[0][10] +
                  mat_A[22][1] * mat_B[1][10] +
                  mat_A[22][2] * mat_B[2][10] +
                  mat_A[22][3] * mat_B[3][10] +
                  mat_A[22][4] * mat_B[4][10] +
                  mat_A[22][5] * mat_B[5][10] +
                  mat_A[22][6] * mat_B[6][10] +
                  mat_A[22][7] * mat_B[7][10] +
                  mat_A[22][8] * mat_B[8][10] +
                  mat_A[22][9] * mat_B[9][10] +
                  mat_A[22][10] * mat_B[10][10] +
                  mat_A[22][11] * mat_B[11][10] +
                  mat_A[22][12] * mat_B[12][10] +
                  mat_A[22][13] * mat_B[13][10] +
                  mat_A[22][14] * mat_B[14][10] +
                  mat_A[22][15] * mat_B[15][10] +
                  mat_A[22][16] * mat_B[16][10] +
                  mat_A[22][17] * mat_B[17][10] +
                  mat_A[22][18] * mat_B[18][10] +
                  mat_A[22][19] * mat_B[19][10] +
                  mat_A[22][20] * mat_B[20][10] +
                  mat_A[22][21] * mat_B[21][10] +
                  mat_A[22][22] * mat_B[22][10] +
                  mat_A[22][23] * mat_B[23][10] +
                  mat_A[22][24] * mat_B[24][10] +
                  mat_A[22][25] * mat_B[25][10] +
                  mat_A[22][26] * mat_B[26][10] +
                  mat_A[22][27] * mat_B[27][10] +
                  mat_A[22][28] * mat_B[28][10] +
                  mat_A[22][29] * mat_B[29][10] +
                  mat_A[22][30] * mat_B[30][10] +
                  mat_A[22][31] * mat_B[31][10];
    mat_C[22][11] <= 
                  mat_A[22][0] * mat_B[0][11] +
                  mat_A[22][1] * mat_B[1][11] +
                  mat_A[22][2] * mat_B[2][11] +
                  mat_A[22][3] * mat_B[3][11] +
                  mat_A[22][4] * mat_B[4][11] +
                  mat_A[22][5] * mat_B[5][11] +
                  mat_A[22][6] * mat_B[6][11] +
                  mat_A[22][7] * mat_B[7][11] +
                  mat_A[22][8] * mat_B[8][11] +
                  mat_A[22][9] * mat_B[9][11] +
                  mat_A[22][10] * mat_B[10][11] +
                  mat_A[22][11] * mat_B[11][11] +
                  mat_A[22][12] * mat_B[12][11] +
                  mat_A[22][13] * mat_B[13][11] +
                  mat_A[22][14] * mat_B[14][11] +
                  mat_A[22][15] * mat_B[15][11] +
                  mat_A[22][16] * mat_B[16][11] +
                  mat_A[22][17] * mat_B[17][11] +
                  mat_A[22][18] * mat_B[18][11] +
                  mat_A[22][19] * mat_B[19][11] +
                  mat_A[22][20] * mat_B[20][11] +
                  mat_A[22][21] * mat_B[21][11] +
                  mat_A[22][22] * mat_B[22][11] +
                  mat_A[22][23] * mat_B[23][11] +
                  mat_A[22][24] * mat_B[24][11] +
                  mat_A[22][25] * mat_B[25][11] +
                  mat_A[22][26] * mat_B[26][11] +
                  mat_A[22][27] * mat_B[27][11] +
                  mat_A[22][28] * mat_B[28][11] +
                  mat_A[22][29] * mat_B[29][11] +
                  mat_A[22][30] * mat_B[30][11] +
                  mat_A[22][31] * mat_B[31][11];
    mat_C[22][12] <= 
                  mat_A[22][0] * mat_B[0][12] +
                  mat_A[22][1] * mat_B[1][12] +
                  mat_A[22][2] * mat_B[2][12] +
                  mat_A[22][3] * mat_B[3][12] +
                  mat_A[22][4] * mat_B[4][12] +
                  mat_A[22][5] * mat_B[5][12] +
                  mat_A[22][6] * mat_B[6][12] +
                  mat_A[22][7] * mat_B[7][12] +
                  mat_A[22][8] * mat_B[8][12] +
                  mat_A[22][9] * mat_B[9][12] +
                  mat_A[22][10] * mat_B[10][12] +
                  mat_A[22][11] * mat_B[11][12] +
                  mat_A[22][12] * mat_B[12][12] +
                  mat_A[22][13] * mat_B[13][12] +
                  mat_A[22][14] * mat_B[14][12] +
                  mat_A[22][15] * mat_B[15][12] +
                  mat_A[22][16] * mat_B[16][12] +
                  mat_A[22][17] * mat_B[17][12] +
                  mat_A[22][18] * mat_B[18][12] +
                  mat_A[22][19] * mat_B[19][12] +
                  mat_A[22][20] * mat_B[20][12] +
                  mat_A[22][21] * mat_B[21][12] +
                  mat_A[22][22] * mat_B[22][12] +
                  mat_A[22][23] * mat_B[23][12] +
                  mat_A[22][24] * mat_B[24][12] +
                  mat_A[22][25] * mat_B[25][12] +
                  mat_A[22][26] * mat_B[26][12] +
                  mat_A[22][27] * mat_B[27][12] +
                  mat_A[22][28] * mat_B[28][12] +
                  mat_A[22][29] * mat_B[29][12] +
                  mat_A[22][30] * mat_B[30][12] +
                  mat_A[22][31] * mat_B[31][12];
    mat_C[22][13] <= 
                  mat_A[22][0] * mat_B[0][13] +
                  mat_A[22][1] * mat_B[1][13] +
                  mat_A[22][2] * mat_B[2][13] +
                  mat_A[22][3] * mat_B[3][13] +
                  mat_A[22][4] * mat_B[4][13] +
                  mat_A[22][5] * mat_B[5][13] +
                  mat_A[22][6] * mat_B[6][13] +
                  mat_A[22][7] * mat_B[7][13] +
                  mat_A[22][8] * mat_B[8][13] +
                  mat_A[22][9] * mat_B[9][13] +
                  mat_A[22][10] * mat_B[10][13] +
                  mat_A[22][11] * mat_B[11][13] +
                  mat_A[22][12] * mat_B[12][13] +
                  mat_A[22][13] * mat_B[13][13] +
                  mat_A[22][14] * mat_B[14][13] +
                  mat_A[22][15] * mat_B[15][13] +
                  mat_A[22][16] * mat_B[16][13] +
                  mat_A[22][17] * mat_B[17][13] +
                  mat_A[22][18] * mat_B[18][13] +
                  mat_A[22][19] * mat_B[19][13] +
                  mat_A[22][20] * mat_B[20][13] +
                  mat_A[22][21] * mat_B[21][13] +
                  mat_A[22][22] * mat_B[22][13] +
                  mat_A[22][23] * mat_B[23][13] +
                  mat_A[22][24] * mat_B[24][13] +
                  mat_A[22][25] * mat_B[25][13] +
                  mat_A[22][26] * mat_B[26][13] +
                  mat_A[22][27] * mat_B[27][13] +
                  mat_A[22][28] * mat_B[28][13] +
                  mat_A[22][29] * mat_B[29][13] +
                  mat_A[22][30] * mat_B[30][13] +
                  mat_A[22][31] * mat_B[31][13];
    mat_C[22][14] <= 
                  mat_A[22][0] * mat_B[0][14] +
                  mat_A[22][1] * mat_B[1][14] +
                  mat_A[22][2] * mat_B[2][14] +
                  mat_A[22][3] * mat_B[3][14] +
                  mat_A[22][4] * mat_B[4][14] +
                  mat_A[22][5] * mat_B[5][14] +
                  mat_A[22][6] * mat_B[6][14] +
                  mat_A[22][7] * mat_B[7][14] +
                  mat_A[22][8] * mat_B[8][14] +
                  mat_A[22][9] * mat_B[9][14] +
                  mat_A[22][10] * mat_B[10][14] +
                  mat_A[22][11] * mat_B[11][14] +
                  mat_A[22][12] * mat_B[12][14] +
                  mat_A[22][13] * mat_B[13][14] +
                  mat_A[22][14] * mat_B[14][14] +
                  mat_A[22][15] * mat_B[15][14] +
                  mat_A[22][16] * mat_B[16][14] +
                  mat_A[22][17] * mat_B[17][14] +
                  mat_A[22][18] * mat_B[18][14] +
                  mat_A[22][19] * mat_B[19][14] +
                  mat_A[22][20] * mat_B[20][14] +
                  mat_A[22][21] * mat_B[21][14] +
                  mat_A[22][22] * mat_B[22][14] +
                  mat_A[22][23] * mat_B[23][14] +
                  mat_A[22][24] * mat_B[24][14] +
                  mat_A[22][25] * mat_B[25][14] +
                  mat_A[22][26] * mat_B[26][14] +
                  mat_A[22][27] * mat_B[27][14] +
                  mat_A[22][28] * mat_B[28][14] +
                  mat_A[22][29] * mat_B[29][14] +
                  mat_A[22][30] * mat_B[30][14] +
                  mat_A[22][31] * mat_B[31][14];
    mat_C[22][15] <= 
                  mat_A[22][0] * mat_B[0][15] +
                  mat_A[22][1] * mat_B[1][15] +
                  mat_A[22][2] * mat_B[2][15] +
                  mat_A[22][3] * mat_B[3][15] +
                  mat_A[22][4] * mat_B[4][15] +
                  mat_A[22][5] * mat_B[5][15] +
                  mat_A[22][6] * mat_B[6][15] +
                  mat_A[22][7] * mat_B[7][15] +
                  mat_A[22][8] * mat_B[8][15] +
                  mat_A[22][9] * mat_B[9][15] +
                  mat_A[22][10] * mat_B[10][15] +
                  mat_A[22][11] * mat_B[11][15] +
                  mat_A[22][12] * mat_B[12][15] +
                  mat_A[22][13] * mat_B[13][15] +
                  mat_A[22][14] * mat_B[14][15] +
                  mat_A[22][15] * mat_B[15][15] +
                  mat_A[22][16] * mat_B[16][15] +
                  mat_A[22][17] * mat_B[17][15] +
                  mat_A[22][18] * mat_B[18][15] +
                  mat_A[22][19] * mat_B[19][15] +
                  mat_A[22][20] * mat_B[20][15] +
                  mat_A[22][21] * mat_B[21][15] +
                  mat_A[22][22] * mat_B[22][15] +
                  mat_A[22][23] * mat_B[23][15] +
                  mat_A[22][24] * mat_B[24][15] +
                  mat_A[22][25] * mat_B[25][15] +
                  mat_A[22][26] * mat_B[26][15] +
                  mat_A[22][27] * mat_B[27][15] +
                  mat_A[22][28] * mat_B[28][15] +
                  mat_A[22][29] * mat_B[29][15] +
                  mat_A[22][30] * mat_B[30][15] +
                  mat_A[22][31] * mat_B[31][15];
    mat_C[22][16] <= 
                  mat_A[22][0] * mat_B[0][16] +
                  mat_A[22][1] * mat_B[1][16] +
                  mat_A[22][2] * mat_B[2][16] +
                  mat_A[22][3] * mat_B[3][16] +
                  mat_A[22][4] * mat_B[4][16] +
                  mat_A[22][5] * mat_B[5][16] +
                  mat_A[22][6] * mat_B[6][16] +
                  mat_A[22][7] * mat_B[7][16] +
                  mat_A[22][8] * mat_B[8][16] +
                  mat_A[22][9] * mat_B[9][16] +
                  mat_A[22][10] * mat_B[10][16] +
                  mat_A[22][11] * mat_B[11][16] +
                  mat_A[22][12] * mat_B[12][16] +
                  mat_A[22][13] * mat_B[13][16] +
                  mat_A[22][14] * mat_B[14][16] +
                  mat_A[22][15] * mat_B[15][16] +
                  mat_A[22][16] * mat_B[16][16] +
                  mat_A[22][17] * mat_B[17][16] +
                  mat_A[22][18] * mat_B[18][16] +
                  mat_A[22][19] * mat_B[19][16] +
                  mat_A[22][20] * mat_B[20][16] +
                  mat_A[22][21] * mat_B[21][16] +
                  mat_A[22][22] * mat_B[22][16] +
                  mat_A[22][23] * mat_B[23][16] +
                  mat_A[22][24] * mat_B[24][16] +
                  mat_A[22][25] * mat_B[25][16] +
                  mat_A[22][26] * mat_B[26][16] +
                  mat_A[22][27] * mat_B[27][16] +
                  mat_A[22][28] * mat_B[28][16] +
                  mat_A[22][29] * mat_B[29][16] +
                  mat_A[22][30] * mat_B[30][16] +
                  mat_A[22][31] * mat_B[31][16];
    mat_C[22][17] <= 
                  mat_A[22][0] * mat_B[0][17] +
                  mat_A[22][1] * mat_B[1][17] +
                  mat_A[22][2] * mat_B[2][17] +
                  mat_A[22][3] * mat_B[3][17] +
                  mat_A[22][4] * mat_B[4][17] +
                  mat_A[22][5] * mat_B[5][17] +
                  mat_A[22][6] * mat_B[6][17] +
                  mat_A[22][7] * mat_B[7][17] +
                  mat_A[22][8] * mat_B[8][17] +
                  mat_A[22][9] * mat_B[9][17] +
                  mat_A[22][10] * mat_B[10][17] +
                  mat_A[22][11] * mat_B[11][17] +
                  mat_A[22][12] * mat_B[12][17] +
                  mat_A[22][13] * mat_B[13][17] +
                  mat_A[22][14] * mat_B[14][17] +
                  mat_A[22][15] * mat_B[15][17] +
                  mat_A[22][16] * mat_B[16][17] +
                  mat_A[22][17] * mat_B[17][17] +
                  mat_A[22][18] * mat_B[18][17] +
                  mat_A[22][19] * mat_B[19][17] +
                  mat_A[22][20] * mat_B[20][17] +
                  mat_A[22][21] * mat_B[21][17] +
                  mat_A[22][22] * mat_B[22][17] +
                  mat_A[22][23] * mat_B[23][17] +
                  mat_A[22][24] * mat_B[24][17] +
                  mat_A[22][25] * mat_B[25][17] +
                  mat_A[22][26] * mat_B[26][17] +
                  mat_A[22][27] * mat_B[27][17] +
                  mat_A[22][28] * mat_B[28][17] +
                  mat_A[22][29] * mat_B[29][17] +
                  mat_A[22][30] * mat_B[30][17] +
                  mat_A[22][31] * mat_B[31][17];
    mat_C[22][18] <= 
                  mat_A[22][0] * mat_B[0][18] +
                  mat_A[22][1] * mat_B[1][18] +
                  mat_A[22][2] * mat_B[2][18] +
                  mat_A[22][3] * mat_B[3][18] +
                  mat_A[22][4] * mat_B[4][18] +
                  mat_A[22][5] * mat_B[5][18] +
                  mat_A[22][6] * mat_B[6][18] +
                  mat_A[22][7] * mat_B[7][18] +
                  mat_A[22][8] * mat_B[8][18] +
                  mat_A[22][9] * mat_B[9][18] +
                  mat_A[22][10] * mat_B[10][18] +
                  mat_A[22][11] * mat_B[11][18] +
                  mat_A[22][12] * mat_B[12][18] +
                  mat_A[22][13] * mat_B[13][18] +
                  mat_A[22][14] * mat_B[14][18] +
                  mat_A[22][15] * mat_B[15][18] +
                  mat_A[22][16] * mat_B[16][18] +
                  mat_A[22][17] * mat_B[17][18] +
                  mat_A[22][18] * mat_B[18][18] +
                  mat_A[22][19] * mat_B[19][18] +
                  mat_A[22][20] * mat_B[20][18] +
                  mat_A[22][21] * mat_B[21][18] +
                  mat_A[22][22] * mat_B[22][18] +
                  mat_A[22][23] * mat_B[23][18] +
                  mat_A[22][24] * mat_B[24][18] +
                  mat_A[22][25] * mat_B[25][18] +
                  mat_A[22][26] * mat_B[26][18] +
                  mat_A[22][27] * mat_B[27][18] +
                  mat_A[22][28] * mat_B[28][18] +
                  mat_A[22][29] * mat_B[29][18] +
                  mat_A[22][30] * mat_B[30][18] +
                  mat_A[22][31] * mat_B[31][18];
    mat_C[22][19] <= 
                  mat_A[22][0] * mat_B[0][19] +
                  mat_A[22][1] * mat_B[1][19] +
                  mat_A[22][2] * mat_B[2][19] +
                  mat_A[22][3] * mat_B[3][19] +
                  mat_A[22][4] * mat_B[4][19] +
                  mat_A[22][5] * mat_B[5][19] +
                  mat_A[22][6] * mat_B[6][19] +
                  mat_A[22][7] * mat_B[7][19] +
                  mat_A[22][8] * mat_B[8][19] +
                  mat_A[22][9] * mat_B[9][19] +
                  mat_A[22][10] * mat_B[10][19] +
                  mat_A[22][11] * mat_B[11][19] +
                  mat_A[22][12] * mat_B[12][19] +
                  mat_A[22][13] * mat_B[13][19] +
                  mat_A[22][14] * mat_B[14][19] +
                  mat_A[22][15] * mat_B[15][19] +
                  mat_A[22][16] * mat_B[16][19] +
                  mat_A[22][17] * mat_B[17][19] +
                  mat_A[22][18] * mat_B[18][19] +
                  mat_A[22][19] * mat_B[19][19] +
                  mat_A[22][20] * mat_B[20][19] +
                  mat_A[22][21] * mat_B[21][19] +
                  mat_A[22][22] * mat_B[22][19] +
                  mat_A[22][23] * mat_B[23][19] +
                  mat_A[22][24] * mat_B[24][19] +
                  mat_A[22][25] * mat_B[25][19] +
                  mat_A[22][26] * mat_B[26][19] +
                  mat_A[22][27] * mat_B[27][19] +
                  mat_A[22][28] * mat_B[28][19] +
                  mat_A[22][29] * mat_B[29][19] +
                  mat_A[22][30] * mat_B[30][19] +
                  mat_A[22][31] * mat_B[31][19];
    mat_C[22][20] <= 
                  mat_A[22][0] * mat_B[0][20] +
                  mat_A[22][1] * mat_B[1][20] +
                  mat_A[22][2] * mat_B[2][20] +
                  mat_A[22][3] * mat_B[3][20] +
                  mat_A[22][4] * mat_B[4][20] +
                  mat_A[22][5] * mat_B[5][20] +
                  mat_A[22][6] * mat_B[6][20] +
                  mat_A[22][7] * mat_B[7][20] +
                  mat_A[22][8] * mat_B[8][20] +
                  mat_A[22][9] * mat_B[9][20] +
                  mat_A[22][10] * mat_B[10][20] +
                  mat_A[22][11] * mat_B[11][20] +
                  mat_A[22][12] * mat_B[12][20] +
                  mat_A[22][13] * mat_B[13][20] +
                  mat_A[22][14] * mat_B[14][20] +
                  mat_A[22][15] * mat_B[15][20] +
                  mat_A[22][16] * mat_B[16][20] +
                  mat_A[22][17] * mat_B[17][20] +
                  mat_A[22][18] * mat_B[18][20] +
                  mat_A[22][19] * mat_B[19][20] +
                  mat_A[22][20] * mat_B[20][20] +
                  mat_A[22][21] * mat_B[21][20] +
                  mat_A[22][22] * mat_B[22][20] +
                  mat_A[22][23] * mat_B[23][20] +
                  mat_A[22][24] * mat_B[24][20] +
                  mat_A[22][25] * mat_B[25][20] +
                  mat_A[22][26] * mat_B[26][20] +
                  mat_A[22][27] * mat_B[27][20] +
                  mat_A[22][28] * mat_B[28][20] +
                  mat_A[22][29] * mat_B[29][20] +
                  mat_A[22][30] * mat_B[30][20] +
                  mat_A[22][31] * mat_B[31][20];
    mat_C[22][21] <= 
                  mat_A[22][0] * mat_B[0][21] +
                  mat_A[22][1] * mat_B[1][21] +
                  mat_A[22][2] * mat_B[2][21] +
                  mat_A[22][3] * mat_B[3][21] +
                  mat_A[22][4] * mat_B[4][21] +
                  mat_A[22][5] * mat_B[5][21] +
                  mat_A[22][6] * mat_B[6][21] +
                  mat_A[22][7] * mat_B[7][21] +
                  mat_A[22][8] * mat_B[8][21] +
                  mat_A[22][9] * mat_B[9][21] +
                  mat_A[22][10] * mat_B[10][21] +
                  mat_A[22][11] * mat_B[11][21] +
                  mat_A[22][12] * mat_B[12][21] +
                  mat_A[22][13] * mat_B[13][21] +
                  mat_A[22][14] * mat_B[14][21] +
                  mat_A[22][15] * mat_B[15][21] +
                  mat_A[22][16] * mat_B[16][21] +
                  mat_A[22][17] * mat_B[17][21] +
                  mat_A[22][18] * mat_B[18][21] +
                  mat_A[22][19] * mat_B[19][21] +
                  mat_A[22][20] * mat_B[20][21] +
                  mat_A[22][21] * mat_B[21][21] +
                  mat_A[22][22] * mat_B[22][21] +
                  mat_A[22][23] * mat_B[23][21] +
                  mat_A[22][24] * mat_B[24][21] +
                  mat_A[22][25] * mat_B[25][21] +
                  mat_A[22][26] * mat_B[26][21] +
                  mat_A[22][27] * mat_B[27][21] +
                  mat_A[22][28] * mat_B[28][21] +
                  mat_A[22][29] * mat_B[29][21] +
                  mat_A[22][30] * mat_B[30][21] +
                  mat_A[22][31] * mat_B[31][21];
    mat_C[22][22] <= 
                  mat_A[22][0] * mat_B[0][22] +
                  mat_A[22][1] * mat_B[1][22] +
                  mat_A[22][2] * mat_B[2][22] +
                  mat_A[22][3] * mat_B[3][22] +
                  mat_A[22][4] * mat_B[4][22] +
                  mat_A[22][5] * mat_B[5][22] +
                  mat_A[22][6] * mat_B[6][22] +
                  mat_A[22][7] * mat_B[7][22] +
                  mat_A[22][8] * mat_B[8][22] +
                  mat_A[22][9] * mat_B[9][22] +
                  mat_A[22][10] * mat_B[10][22] +
                  mat_A[22][11] * mat_B[11][22] +
                  mat_A[22][12] * mat_B[12][22] +
                  mat_A[22][13] * mat_B[13][22] +
                  mat_A[22][14] * mat_B[14][22] +
                  mat_A[22][15] * mat_B[15][22] +
                  mat_A[22][16] * mat_B[16][22] +
                  mat_A[22][17] * mat_B[17][22] +
                  mat_A[22][18] * mat_B[18][22] +
                  mat_A[22][19] * mat_B[19][22] +
                  mat_A[22][20] * mat_B[20][22] +
                  mat_A[22][21] * mat_B[21][22] +
                  mat_A[22][22] * mat_B[22][22] +
                  mat_A[22][23] * mat_B[23][22] +
                  mat_A[22][24] * mat_B[24][22] +
                  mat_A[22][25] * mat_B[25][22] +
                  mat_A[22][26] * mat_B[26][22] +
                  mat_A[22][27] * mat_B[27][22] +
                  mat_A[22][28] * mat_B[28][22] +
                  mat_A[22][29] * mat_B[29][22] +
                  mat_A[22][30] * mat_B[30][22] +
                  mat_A[22][31] * mat_B[31][22];
    mat_C[22][23] <= 
                  mat_A[22][0] * mat_B[0][23] +
                  mat_A[22][1] * mat_B[1][23] +
                  mat_A[22][2] * mat_B[2][23] +
                  mat_A[22][3] * mat_B[3][23] +
                  mat_A[22][4] * mat_B[4][23] +
                  mat_A[22][5] * mat_B[5][23] +
                  mat_A[22][6] * mat_B[6][23] +
                  mat_A[22][7] * mat_B[7][23] +
                  mat_A[22][8] * mat_B[8][23] +
                  mat_A[22][9] * mat_B[9][23] +
                  mat_A[22][10] * mat_B[10][23] +
                  mat_A[22][11] * mat_B[11][23] +
                  mat_A[22][12] * mat_B[12][23] +
                  mat_A[22][13] * mat_B[13][23] +
                  mat_A[22][14] * mat_B[14][23] +
                  mat_A[22][15] * mat_B[15][23] +
                  mat_A[22][16] * mat_B[16][23] +
                  mat_A[22][17] * mat_B[17][23] +
                  mat_A[22][18] * mat_B[18][23] +
                  mat_A[22][19] * mat_B[19][23] +
                  mat_A[22][20] * mat_B[20][23] +
                  mat_A[22][21] * mat_B[21][23] +
                  mat_A[22][22] * mat_B[22][23] +
                  mat_A[22][23] * mat_B[23][23] +
                  mat_A[22][24] * mat_B[24][23] +
                  mat_A[22][25] * mat_B[25][23] +
                  mat_A[22][26] * mat_B[26][23] +
                  mat_A[22][27] * mat_B[27][23] +
                  mat_A[22][28] * mat_B[28][23] +
                  mat_A[22][29] * mat_B[29][23] +
                  mat_A[22][30] * mat_B[30][23] +
                  mat_A[22][31] * mat_B[31][23];
    mat_C[22][24] <= 
                  mat_A[22][0] * mat_B[0][24] +
                  mat_A[22][1] * mat_B[1][24] +
                  mat_A[22][2] * mat_B[2][24] +
                  mat_A[22][3] * mat_B[3][24] +
                  mat_A[22][4] * mat_B[4][24] +
                  mat_A[22][5] * mat_B[5][24] +
                  mat_A[22][6] * mat_B[6][24] +
                  mat_A[22][7] * mat_B[7][24] +
                  mat_A[22][8] * mat_B[8][24] +
                  mat_A[22][9] * mat_B[9][24] +
                  mat_A[22][10] * mat_B[10][24] +
                  mat_A[22][11] * mat_B[11][24] +
                  mat_A[22][12] * mat_B[12][24] +
                  mat_A[22][13] * mat_B[13][24] +
                  mat_A[22][14] * mat_B[14][24] +
                  mat_A[22][15] * mat_B[15][24] +
                  mat_A[22][16] * mat_B[16][24] +
                  mat_A[22][17] * mat_B[17][24] +
                  mat_A[22][18] * mat_B[18][24] +
                  mat_A[22][19] * mat_B[19][24] +
                  mat_A[22][20] * mat_B[20][24] +
                  mat_A[22][21] * mat_B[21][24] +
                  mat_A[22][22] * mat_B[22][24] +
                  mat_A[22][23] * mat_B[23][24] +
                  mat_A[22][24] * mat_B[24][24] +
                  mat_A[22][25] * mat_B[25][24] +
                  mat_A[22][26] * mat_B[26][24] +
                  mat_A[22][27] * mat_B[27][24] +
                  mat_A[22][28] * mat_B[28][24] +
                  mat_A[22][29] * mat_B[29][24] +
                  mat_A[22][30] * mat_B[30][24] +
                  mat_A[22][31] * mat_B[31][24];
    mat_C[22][25] <= 
                  mat_A[22][0] * mat_B[0][25] +
                  mat_A[22][1] * mat_B[1][25] +
                  mat_A[22][2] * mat_B[2][25] +
                  mat_A[22][3] * mat_B[3][25] +
                  mat_A[22][4] * mat_B[4][25] +
                  mat_A[22][5] * mat_B[5][25] +
                  mat_A[22][6] * mat_B[6][25] +
                  mat_A[22][7] * mat_B[7][25] +
                  mat_A[22][8] * mat_B[8][25] +
                  mat_A[22][9] * mat_B[9][25] +
                  mat_A[22][10] * mat_B[10][25] +
                  mat_A[22][11] * mat_B[11][25] +
                  mat_A[22][12] * mat_B[12][25] +
                  mat_A[22][13] * mat_B[13][25] +
                  mat_A[22][14] * mat_B[14][25] +
                  mat_A[22][15] * mat_B[15][25] +
                  mat_A[22][16] * mat_B[16][25] +
                  mat_A[22][17] * mat_B[17][25] +
                  mat_A[22][18] * mat_B[18][25] +
                  mat_A[22][19] * mat_B[19][25] +
                  mat_A[22][20] * mat_B[20][25] +
                  mat_A[22][21] * mat_B[21][25] +
                  mat_A[22][22] * mat_B[22][25] +
                  mat_A[22][23] * mat_B[23][25] +
                  mat_A[22][24] * mat_B[24][25] +
                  mat_A[22][25] * mat_B[25][25] +
                  mat_A[22][26] * mat_B[26][25] +
                  mat_A[22][27] * mat_B[27][25] +
                  mat_A[22][28] * mat_B[28][25] +
                  mat_A[22][29] * mat_B[29][25] +
                  mat_A[22][30] * mat_B[30][25] +
                  mat_A[22][31] * mat_B[31][25];
    mat_C[22][26] <= 
                  mat_A[22][0] * mat_B[0][26] +
                  mat_A[22][1] * mat_B[1][26] +
                  mat_A[22][2] * mat_B[2][26] +
                  mat_A[22][3] * mat_B[3][26] +
                  mat_A[22][4] * mat_B[4][26] +
                  mat_A[22][5] * mat_B[5][26] +
                  mat_A[22][6] * mat_B[6][26] +
                  mat_A[22][7] * mat_B[7][26] +
                  mat_A[22][8] * mat_B[8][26] +
                  mat_A[22][9] * mat_B[9][26] +
                  mat_A[22][10] * mat_B[10][26] +
                  mat_A[22][11] * mat_B[11][26] +
                  mat_A[22][12] * mat_B[12][26] +
                  mat_A[22][13] * mat_B[13][26] +
                  mat_A[22][14] * mat_B[14][26] +
                  mat_A[22][15] * mat_B[15][26] +
                  mat_A[22][16] * mat_B[16][26] +
                  mat_A[22][17] * mat_B[17][26] +
                  mat_A[22][18] * mat_B[18][26] +
                  mat_A[22][19] * mat_B[19][26] +
                  mat_A[22][20] * mat_B[20][26] +
                  mat_A[22][21] * mat_B[21][26] +
                  mat_A[22][22] * mat_B[22][26] +
                  mat_A[22][23] * mat_B[23][26] +
                  mat_A[22][24] * mat_B[24][26] +
                  mat_A[22][25] * mat_B[25][26] +
                  mat_A[22][26] * mat_B[26][26] +
                  mat_A[22][27] * mat_B[27][26] +
                  mat_A[22][28] * mat_B[28][26] +
                  mat_A[22][29] * mat_B[29][26] +
                  mat_A[22][30] * mat_B[30][26] +
                  mat_A[22][31] * mat_B[31][26];
    mat_C[22][27] <= 
                  mat_A[22][0] * mat_B[0][27] +
                  mat_A[22][1] * mat_B[1][27] +
                  mat_A[22][2] * mat_B[2][27] +
                  mat_A[22][3] * mat_B[3][27] +
                  mat_A[22][4] * mat_B[4][27] +
                  mat_A[22][5] * mat_B[5][27] +
                  mat_A[22][6] * mat_B[6][27] +
                  mat_A[22][7] * mat_B[7][27] +
                  mat_A[22][8] * mat_B[8][27] +
                  mat_A[22][9] * mat_B[9][27] +
                  mat_A[22][10] * mat_B[10][27] +
                  mat_A[22][11] * mat_B[11][27] +
                  mat_A[22][12] * mat_B[12][27] +
                  mat_A[22][13] * mat_B[13][27] +
                  mat_A[22][14] * mat_B[14][27] +
                  mat_A[22][15] * mat_B[15][27] +
                  mat_A[22][16] * mat_B[16][27] +
                  mat_A[22][17] * mat_B[17][27] +
                  mat_A[22][18] * mat_B[18][27] +
                  mat_A[22][19] * mat_B[19][27] +
                  mat_A[22][20] * mat_B[20][27] +
                  mat_A[22][21] * mat_B[21][27] +
                  mat_A[22][22] * mat_B[22][27] +
                  mat_A[22][23] * mat_B[23][27] +
                  mat_A[22][24] * mat_B[24][27] +
                  mat_A[22][25] * mat_B[25][27] +
                  mat_A[22][26] * mat_B[26][27] +
                  mat_A[22][27] * mat_B[27][27] +
                  mat_A[22][28] * mat_B[28][27] +
                  mat_A[22][29] * mat_B[29][27] +
                  mat_A[22][30] * mat_B[30][27] +
                  mat_A[22][31] * mat_B[31][27];
    mat_C[22][28] <= 
                  mat_A[22][0] * mat_B[0][28] +
                  mat_A[22][1] * mat_B[1][28] +
                  mat_A[22][2] * mat_B[2][28] +
                  mat_A[22][3] * mat_B[3][28] +
                  mat_A[22][4] * mat_B[4][28] +
                  mat_A[22][5] * mat_B[5][28] +
                  mat_A[22][6] * mat_B[6][28] +
                  mat_A[22][7] * mat_B[7][28] +
                  mat_A[22][8] * mat_B[8][28] +
                  mat_A[22][9] * mat_B[9][28] +
                  mat_A[22][10] * mat_B[10][28] +
                  mat_A[22][11] * mat_B[11][28] +
                  mat_A[22][12] * mat_B[12][28] +
                  mat_A[22][13] * mat_B[13][28] +
                  mat_A[22][14] * mat_B[14][28] +
                  mat_A[22][15] * mat_B[15][28] +
                  mat_A[22][16] * mat_B[16][28] +
                  mat_A[22][17] * mat_B[17][28] +
                  mat_A[22][18] * mat_B[18][28] +
                  mat_A[22][19] * mat_B[19][28] +
                  mat_A[22][20] * mat_B[20][28] +
                  mat_A[22][21] * mat_B[21][28] +
                  mat_A[22][22] * mat_B[22][28] +
                  mat_A[22][23] * mat_B[23][28] +
                  mat_A[22][24] * mat_B[24][28] +
                  mat_A[22][25] * mat_B[25][28] +
                  mat_A[22][26] * mat_B[26][28] +
                  mat_A[22][27] * mat_B[27][28] +
                  mat_A[22][28] * mat_B[28][28] +
                  mat_A[22][29] * mat_B[29][28] +
                  mat_A[22][30] * mat_B[30][28] +
                  mat_A[22][31] * mat_B[31][28];
    mat_C[22][29] <= 
                  mat_A[22][0] * mat_B[0][29] +
                  mat_A[22][1] * mat_B[1][29] +
                  mat_A[22][2] * mat_B[2][29] +
                  mat_A[22][3] * mat_B[3][29] +
                  mat_A[22][4] * mat_B[4][29] +
                  mat_A[22][5] * mat_B[5][29] +
                  mat_A[22][6] * mat_B[6][29] +
                  mat_A[22][7] * mat_B[7][29] +
                  mat_A[22][8] * mat_B[8][29] +
                  mat_A[22][9] * mat_B[9][29] +
                  mat_A[22][10] * mat_B[10][29] +
                  mat_A[22][11] * mat_B[11][29] +
                  mat_A[22][12] * mat_B[12][29] +
                  mat_A[22][13] * mat_B[13][29] +
                  mat_A[22][14] * mat_B[14][29] +
                  mat_A[22][15] * mat_B[15][29] +
                  mat_A[22][16] * mat_B[16][29] +
                  mat_A[22][17] * mat_B[17][29] +
                  mat_A[22][18] * mat_B[18][29] +
                  mat_A[22][19] * mat_B[19][29] +
                  mat_A[22][20] * mat_B[20][29] +
                  mat_A[22][21] * mat_B[21][29] +
                  mat_A[22][22] * mat_B[22][29] +
                  mat_A[22][23] * mat_B[23][29] +
                  mat_A[22][24] * mat_B[24][29] +
                  mat_A[22][25] * mat_B[25][29] +
                  mat_A[22][26] * mat_B[26][29] +
                  mat_A[22][27] * mat_B[27][29] +
                  mat_A[22][28] * mat_B[28][29] +
                  mat_A[22][29] * mat_B[29][29] +
                  mat_A[22][30] * mat_B[30][29] +
                  mat_A[22][31] * mat_B[31][29];
    mat_C[22][30] <= 
                  mat_A[22][0] * mat_B[0][30] +
                  mat_A[22][1] * mat_B[1][30] +
                  mat_A[22][2] * mat_B[2][30] +
                  mat_A[22][3] * mat_B[3][30] +
                  mat_A[22][4] * mat_B[4][30] +
                  mat_A[22][5] * mat_B[5][30] +
                  mat_A[22][6] * mat_B[6][30] +
                  mat_A[22][7] * mat_B[7][30] +
                  mat_A[22][8] * mat_B[8][30] +
                  mat_A[22][9] * mat_B[9][30] +
                  mat_A[22][10] * mat_B[10][30] +
                  mat_A[22][11] * mat_B[11][30] +
                  mat_A[22][12] * mat_B[12][30] +
                  mat_A[22][13] * mat_B[13][30] +
                  mat_A[22][14] * mat_B[14][30] +
                  mat_A[22][15] * mat_B[15][30] +
                  mat_A[22][16] * mat_B[16][30] +
                  mat_A[22][17] * mat_B[17][30] +
                  mat_A[22][18] * mat_B[18][30] +
                  mat_A[22][19] * mat_B[19][30] +
                  mat_A[22][20] * mat_B[20][30] +
                  mat_A[22][21] * mat_B[21][30] +
                  mat_A[22][22] * mat_B[22][30] +
                  mat_A[22][23] * mat_B[23][30] +
                  mat_A[22][24] * mat_B[24][30] +
                  mat_A[22][25] * mat_B[25][30] +
                  mat_A[22][26] * mat_B[26][30] +
                  mat_A[22][27] * mat_B[27][30] +
                  mat_A[22][28] * mat_B[28][30] +
                  mat_A[22][29] * mat_B[29][30] +
                  mat_A[22][30] * mat_B[30][30] +
                  mat_A[22][31] * mat_B[31][30];
    mat_C[22][31] <= 
                  mat_A[22][0] * mat_B[0][31] +
                  mat_A[22][1] * mat_B[1][31] +
                  mat_A[22][2] * mat_B[2][31] +
                  mat_A[22][3] * mat_B[3][31] +
                  mat_A[22][4] * mat_B[4][31] +
                  mat_A[22][5] * mat_B[5][31] +
                  mat_A[22][6] * mat_B[6][31] +
                  mat_A[22][7] * mat_B[7][31] +
                  mat_A[22][8] * mat_B[8][31] +
                  mat_A[22][9] * mat_B[9][31] +
                  mat_A[22][10] * mat_B[10][31] +
                  mat_A[22][11] * mat_B[11][31] +
                  mat_A[22][12] * mat_B[12][31] +
                  mat_A[22][13] * mat_B[13][31] +
                  mat_A[22][14] * mat_B[14][31] +
                  mat_A[22][15] * mat_B[15][31] +
                  mat_A[22][16] * mat_B[16][31] +
                  mat_A[22][17] * mat_B[17][31] +
                  mat_A[22][18] * mat_B[18][31] +
                  mat_A[22][19] * mat_B[19][31] +
                  mat_A[22][20] * mat_B[20][31] +
                  mat_A[22][21] * mat_B[21][31] +
                  mat_A[22][22] * mat_B[22][31] +
                  mat_A[22][23] * mat_B[23][31] +
                  mat_A[22][24] * mat_B[24][31] +
                  mat_A[22][25] * mat_B[25][31] +
                  mat_A[22][26] * mat_B[26][31] +
                  mat_A[22][27] * mat_B[27][31] +
                  mat_A[22][28] * mat_B[28][31] +
                  mat_A[22][29] * mat_B[29][31] +
                  mat_A[22][30] * mat_B[30][31] +
                  mat_A[22][31] * mat_B[31][31];
    mat_C[23][0] <= 
                  mat_A[23][0] * mat_B[0][0] +
                  mat_A[23][1] * mat_B[1][0] +
                  mat_A[23][2] * mat_B[2][0] +
                  mat_A[23][3] * mat_B[3][0] +
                  mat_A[23][4] * mat_B[4][0] +
                  mat_A[23][5] * mat_B[5][0] +
                  mat_A[23][6] * mat_B[6][0] +
                  mat_A[23][7] * mat_B[7][0] +
                  mat_A[23][8] * mat_B[8][0] +
                  mat_A[23][9] * mat_B[9][0] +
                  mat_A[23][10] * mat_B[10][0] +
                  mat_A[23][11] * mat_B[11][0] +
                  mat_A[23][12] * mat_B[12][0] +
                  mat_A[23][13] * mat_B[13][0] +
                  mat_A[23][14] * mat_B[14][0] +
                  mat_A[23][15] * mat_B[15][0] +
                  mat_A[23][16] * mat_B[16][0] +
                  mat_A[23][17] * mat_B[17][0] +
                  mat_A[23][18] * mat_B[18][0] +
                  mat_A[23][19] * mat_B[19][0] +
                  mat_A[23][20] * mat_B[20][0] +
                  mat_A[23][21] * mat_B[21][0] +
                  mat_A[23][22] * mat_B[22][0] +
                  mat_A[23][23] * mat_B[23][0] +
                  mat_A[23][24] * mat_B[24][0] +
                  mat_A[23][25] * mat_B[25][0] +
                  mat_A[23][26] * mat_B[26][0] +
                  mat_A[23][27] * mat_B[27][0] +
                  mat_A[23][28] * mat_B[28][0] +
                  mat_A[23][29] * mat_B[29][0] +
                  mat_A[23][30] * mat_B[30][0] +
                  mat_A[23][31] * mat_B[31][0];
    mat_C[23][1] <= 
                  mat_A[23][0] * mat_B[0][1] +
                  mat_A[23][1] * mat_B[1][1] +
                  mat_A[23][2] * mat_B[2][1] +
                  mat_A[23][3] * mat_B[3][1] +
                  mat_A[23][4] * mat_B[4][1] +
                  mat_A[23][5] * mat_B[5][1] +
                  mat_A[23][6] * mat_B[6][1] +
                  mat_A[23][7] * mat_B[7][1] +
                  mat_A[23][8] * mat_B[8][1] +
                  mat_A[23][9] * mat_B[9][1] +
                  mat_A[23][10] * mat_B[10][1] +
                  mat_A[23][11] * mat_B[11][1] +
                  mat_A[23][12] * mat_B[12][1] +
                  mat_A[23][13] * mat_B[13][1] +
                  mat_A[23][14] * mat_B[14][1] +
                  mat_A[23][15] * mat_B[15][1] +
                  mat_A[23][16] * mat_B[16][1] +
                  mat_A[23][17] * mat_B[17][1] +
                  mat_A[23][18] * mat_B[18][1] +
                  mat_A[23][19] * mat_B[19][1] +
                  mat_A[23][20] * mat_B[20][1] +
                  mat_A[23][21] * mat_B[21][1] +
                  mat_A[23][22] * mat_B[22][1] +
                  mat_A[23][23] * mat_B[23][1] +
                  mat_A[23][24] * mat_B[24][1] +
                  mat_A[23][25] * mat_B[25][1] +
                  mat_A[23][26] * mat_B[26][1] +
                  mat_A[23][27] * mat_B[27][1] +
                  mat_A[23][28] * mat_B[28][1] +
                  mat_A[23][29] * mat_B[29][1] +
                  mat_A[23][30] * mat_B[30][1] +
                  mat_A[23][31] * mat_B[31][1];
    mat_C[23][2] <= 
                  mat_A[23][0] * mat_B[0][2] +
                  mat_A[23][1] * mat_B[1][2] +
                  mat_A[23][2] * mat_B[2][2] +
                  mat_A[23][3] * mat_B[3][2] +
                  mat_A[23][4] * mat_B[4][2] +
                  mat_A[23][5] * mat_B[5][2] +
                  mat_A[23][6] * mat_B[6][2] +
                  mat_A[23][7] * mat_B[7][2] +
                  mat_A[23][8] * mat_B[8][2] +
                  mat_A[23][9] * mat_B[9][2] +
                  mat_A[23][10] * mat_B[10][2] +
                  mat_A[23][11] * mat_B[11][2] +
                  mat_A[23][12] * mat_B[12][2] +
                  mat_A[23][13] * mat_B[13][2] +
                  mat_A[23][14] * mat_B[14][2] +
                  mat_A[23][15] * mat_B[15][2] +
                  mat_A[23][16] * mat_B[16][2] +
                  mat_A[23][17] * mat_B[17][2] +
                  mat_A[23][18] * mat_B[18][2] +
                  mat_A[23][19] * mat_B[19][2] +
                  mat_A[23][20] * mat_B[20][2] +
                  mat_A[23][21] * mat_B[21][2] +
                  mat_A[23][22] * mat_B[22][2] +
                  mat_A[23][23] * mat_B[23][2] +
                  mat_A[23][24] * mat_B[24][2] +
                  mat_A[23][25] * mat_B[25][2] +
                  mat_A[23][26] * mat_B[26][2] +
                  mat_A[23][27] * mat_B[27][2] +
                  mat_A[23][28] * mat_B[28][2] +
                  mat_A[23][29] * mat_B[29][2] +
                  mat_A[23][30] * mat_B[30][2] +
                  mat_A[23][31] * mat_B[31][2];
    mat_C[23][3] <= 
                  mat_A[23][0] * mat_B[0][3] +
                  mat_A[23][1] * mat_B[1][3] +
                  mat_A[23][2] * mat_B[2][3] +
                  mat_A[23][3] * mat_B[3][3] +
                  mat_A[23][4] * mat_B[4][3] +
                  mat_A[23][5] * mat_B[5][3] +
                  mat_A[23][6] * mat_B[6][3] +
                  mat_A[23][7] * mat_B[7][3] +
                  mat_A[23][8] * mat_B[8][3] +
                  mat_A[23][9] * mat_B[9][3] +
                  mat_A[23][10] * mat_B[10][3] +
                  mat_A[23][11] * mat_B[11][3] +
                  mat_A[23][12] * mat_B[12][3] +
                  mat_A[23][13] * mat_B[13][3] +
                  mat_A[23][14] * mat_B[14][3] +
                  mat_A[23][15] * mat_B[15][3] +
                  mat_A[23][16] * mat_B[16][3] +
                  mat_A[23][17] * mat_B[17][3] +
                  mat_A[23][18] * mat_B[18][3] +
                  mat_A[23][19] * mat_B[19][3] +
                  mat_A[23][20] * mat_B[20][3] +
                  mat_A[23][21] * mat_B[21][3] +
                  mat_A[23][22] * mat_B[22][3] +
                  mat_A[23][23] * mat_B[23][3] +
                  mat_A[23][24] * mat_B[24][3] +
                  mat_A[23][25] * mat_B[25][3] +
                  mat_A[23][26] * mat_B[26][3] +
                  mat_A[23][27] * mat_B[27][3] +
                  mat_A[23][28] * mat_B[28][3] +
                  mat_A[23][29] * mat_B[29][3] +
                  mat_A[23][30] * mat_B[30][3] +
                  mat_A[23][31] * mat_B[31][3];
    mat_C[23][4] <= 
                  mat_A[23][0] * mat_B[0][4] +
                  mat_A[23][1] * mat_B[1][4] +
                  mat_A[23][2] * mat_B[2][4] +
                  mat_A[23][3] * mat_B[3][4] +
                  mat_A[23][4] * mat_B[4][4] +
                  mat_A[23][5] * mat_B[5][4] +
                  mat_A[23][6] * mat_B[6][4] +
                  mat_A[23][7] * mat_B[7][4] +
                  mat_A[23][8] * mat_B[8][4] +
                  mat_A[23][9] * mat_B[9][4] +
                  mat_A[23][10] * mat_B[10][4] +
                  mat_A[23][11] * mat_B[11][4] +
                  mat_A[23][12] * mat_B[12][4] +
                  mat_A[23][13] * mat_B[13][4] +
                  mat_A[23][14] * mat_B[14][4] +
                  mat_A[23][15] * mat_B[15][4] +
                  mat_A[23][16] * mat_B[16][4] +
                  mat_A[23][17] * mat_B[17][4] +
                  mat_A[23][18] * mat_B[18][4] +
                  mat_A[23][19] * mat_B[19][4] +
                  mat_A[23][20] * mat_B[20][4] +
                  mat_A[23][21] * mat_B[21][4] +
                  mat_A[23][22] * mat_B[22][4] +
                  mat_A[23][23] * mat_B[23][4] +
                  mat_A[23][24] * mat_B[24][4] +
                  mat_A[23][25] * mat_B[25][4] +
                  mat_A[23][26] * mat_B[26][4] +
                  mat_A[23][27] * mat_B[27][4] +
                  mat_A[23][28] * mat_B[28][4] +
                  mat_A[23][29] * mat_B[29][4] +
                  mat_A[23][30] * mat_B[30][4] +
                  mat_A[23][31] * mat_B[31][4];
    mat_C[23][5] <= 
                  mat_A[23][0] * mat_B[0][5] +
                  mat_A[23][1] * mat_B[1][5] +
                  mat_A[23][2] * mat_B[2][5] +
                  mat_A[23][3] * mat_B[3][5] +
                  mat_A[23][4] * mat_B[4][5] +
                  mat_A[23][5] * mat_B[5][5] +
                  mat_A[23][6] * mat_B[6][5] +
                  mat_A[23][7] * mat_B[7][5] +
                  mat_A[23][8] * mat_B[8][5] +
                  mat_A[23][9] * mat_B[9][5] +
                  mat_A[23][10] * mat_B[10][5] +
                  mat_A[23][11] * mat_B[11][5] +
                  mat_A[23][12] * mat_B[12][5] +
                  mat_A[23][13] * mat_B[13][5] +
                  mat_A[23][14] * mat_B[14][5] +
                  mat_A[23][15] * mat_B[15][5] +
                  mat_A[23][16] * mat_B[16][5] +
                  mat_A[23][17] * mat_B[17][5] +
                  mat_A[23][18] * mat_B[18][5] +
                  mat_A[23][19] * mat_B[19][5] +
                  mat_A[23][20] * mat_B[20][5] +
                  mat_A[23][21] * mat_B[21][5] +
                  mat_A[23][22] * mat_B[22][5] +
                  mat_A[23][23] * mat_B[23][5] +
                  mat_A[23][24] * mat_B[24][5] +
                  mat_A[23][25] * mat_B[25][5] +
                  mat_A[23][26] * mat_B[26][5] +
                  mat_A[23][27] * mat_B[27][5] +
                  mat_A[23][28] * mat_B[28][5] +
                  mat_A[23][29] * mat_B[29][5] +
                  mat_A[23][30] * mat_B[30][5] +
                  mat_A[23][31] * mat_B[31][5];
    mat_C[23][6] <= 
                  mat_A[23][0] * mat_B[0][6] +
                  mat_A[23][1] * mat_B[1][6] +
                  mat_A[23][2] * mat_B[2][6] +
                  mat_A[23][3] * mat_B[3][6] +
                  mat_A[23][4] * mat_B[4][6] +
                  mat_A[23][5] * mat_B[5][6] +
                  mat_A[23][6] * mat_B[6][6] +
                  mat_A[23][7] * mat_B[7][6] +
                  mat_A[23][8] * mat_B[8][6] +
                  mat_A[23][9] * mat_B[9][6] +
                  mat_A[23][10] * mat_B[10][6] +
                  mat_A[23][11] * mat_B[11][6] +
                  mat_A[23][12] * mat_B[12][6] +
                  mat_A[23][13] * mat_B[13][6] +
                  mat_A[23][14] * mat_B[14][6] +
                  mat_A[23][15] * mat_B[15][6] +
                  mat_A[23][16] * mat_B[16][6] +
                  mat_A[23][17] * mat_B[17][6] +
                  mat_A[23][18] * mat_B[18][6] +
                  mat_A[23][19] * mat_B[19][6] +
                  mat_A[23][20] * mat_B[20][6] +
                  mat_A[23][21] * mat_B[21][6] +
                  mat_A[23][22] * mat_B[22][6] +
                  mat_A[23][23] * mat_B[23][6] +
                  mat_A[23][24] * mat_B[24][6] +
                  mat_A[23][25] * mat_B[25][6] +
                  mat_A[23][26] * mat_B[26][6] +
                  mat_A[23][27] * mat_B[27][6] +
                  mat_A[23][28] * mat_B[28][6] +
                  mat_A[23][29] * mat_B[29][6] +
                  mat_A[23][30] * mat_B[30][6] +
                  mat_A[23][31] * mat_B[31][6];
    mat_C[23][7] <= 
                  mat_A[23][0] * mat_B[0][7] +
                  mat_A[23][1] * mat_B[1][7] +
                  mat_A[23][2] * mat_B[2][7] +
                  mat_A[23][3] * mat_B[3][7] +
                  mat_A[23][4] * mat_B[4][7] +
                  mat_A[23][5] * mat_B[5][7] +
                  mat_A[23][6] * mat_B[6][7] +
                  mat_A[23][7] * mat_B[7][7] +
                  mat_A[23][8] * mat_B[8][7] +
                  mat_A[23][9] * mat_B[9][7] +
                  mat_A[23][10] * mat_B[10][7] +
                  mat_A[23][11] * mat_B[11][7] +
                  mat_A[23][12] * mat_B[12][7] +
                  mat_A[23][13] * mat_B[13][7] +
                  mat_A[23][14] * mat_B[14][7] +
                  mat_A[23][15] * mat_B[15][7] +
                  mat_A[23][16] * mat_B[16][7] +
                  mat_A[23][17] * mat_B[17][7] +
                  mat_A[23][18] * mat_B[18][7] +
                  mat_A[23][19] * mat_B[19][7] +
                  mat_A[23][20] * mat_B[20][7] +
                  mat_A[23][21] * mat_B[21][7] +
                  mat_A[23][22] * mat_B[22][7] +
                  mat_A[23][23] * mat_B[23][7] +
                  mat_A[23][24] * mat_B[24][7] +
                  mat_A[23][25] * mat_B[25][7] +
                  mat_A[23][26] * mat_B[26][7] +
                  mat_A[23][27] * mat_B[27][7] +
                  mat_A[23][28] * mat_B[28][7] +
                  mat_A[23][29] * mat_B[29][7] +
                  mat_A[23][30] * mat_B[30][7] +
                  mat_A[23][31] * mat_B[31][7];
    mat_C[23][8] <= 
                  mat_A[23][0] * mat_B[0][8] +
                  mat_A[23][1] * mat_B[1][8] +
                  mat_A[23][2] * mat_B[2][8] +
                  mat_A[23][3] * mat_B[3][8] +
                  mat_A[23][4] * mat_B[4][8] +
                  mat_A[23][5] * mat_B[5][8] +
                  mat_A[23][6] * mat_B[6][8] +
                  mat_A[23][7] * mat_B[7][8] +
                  mat_A[23][8] * mat_B[8][8] +
                  mat_A[23][9] * mat_B[9][8] +
                  mat_A[23][10] * mat_B[10][8] +
                  mat_A[23][11] * mat_B[11][8] +
                  mat_A[23][12] * mat_B[12][8] +
                  mat_A[23][13] * mat_B[13][8] +
                  mat_A[23][14] * mat_B[14][8] +
                  mat_A[23][15] * mat_B[15][8] +
                  mat_A[23][16] * mat_B[16][8] +
                  mat_A[23][17] * mat_B[17][8] +
                  mat_A[23][18] * mat_B[18][8] +
                  mat_A[23][19] * mat_B[19][8] +
                  mat_A[23][20] * mat_B[20][8] +
                  mat_A[23][21] * mat_B[21][8] +
                  mat_A[23][22] * mat_B[22][8] +
                  mat_A[23][23] * mat_B[23][8] +
                  mat_A[23][24] * mat_B[24][8] +
                  mat_A[23][25] * mat_B[25][8] +
                  mat_A[23][26] * mat_B[26][8] +
                  mat_A[23][27] * mat_B[27][8] +
                  mat_A[23][28] * mat_B[28][8] +
                  mat_A[23][29] * mat_B[29][8] +
                  mat_A[23][30] * mat_B[30][8] +
                  mat_A[23][31] * mat_B[31][8];
    mat_C[23][9] <= 
                  mat_A[23][0] * mat_B[0][9] +
                  mat_A[23][1] * mat_B[1][9] +
                  mat_A[23][2] * mat_B[2][9] +
                  mat_A[23][3] * mat_B[3][9] +
                  mat_A[23][4] * mat_B[4][9] +
                  mat_A[23][5] * mat_B[5][9] +
                  mat_A[23][6] * mat_B[6][9] +
                  mat_A[23][7] * mat_B[7][9] +
                  mat_A[23][8] * mat_B[8][9] +
                  mat_A[23][9] * mat_B[9][9] +
                  mat_A[23][10] * mat_B[10][9] +
                  mat_A[23][11] * mat_B[11][9] +
                  mat_A[23][12] * mat_B[12][9] +
                  mat_A[23][13] * mat_B[13][9] +
                  mat_A[23][14] * mat_B[14][9] +
                  mat_A[23][15] * mat_B[15][9] +
                  mat_A[23][16] * mat_B[16][9] +
                  mat_A[23][17] * mat_B[17][9] +
                  mat_A[23][18] * mat_B[18][9] +
                  mat_A[23][19] * mat_B[19][9] +
                  mat_A[23][20] * mat_B[20][9] +
                  mat_A[23][21] * mat_B[21][9] +
                  mat_A[23][22] * mat_B[22][9] +
                  mat_A[23][23] * mat_B[23][9] +
                  mat_A[23][24] * mat_B[24][9] +
                  mat_A[23][25] * mat_B[25][9] +
                  mat_A[23][26] * mat_B[26][9] +
                  mat_A[23][27] * mat_B[27][9] +
                  mat_A[23][28] * mat_B[28][9] +
                  mat_A[23][29] * mat_B[29][9] +
                  mat_A[23][30] * mat_B[30][9] +
                  mat_A[23][31] * mat_B[31][9];
    mat_C[23][10] <= 
                  mat_A[23][0] * mat_B[0][10] +
                  mat_A[23][1] * mat_B[1][10] +
                  mat_A[23][2] * mat_B[2][10] +
                  mat_A[23][3] * mat_B[3][10] +
                  mat_A[23][4] * mat_B[4][10] +
                  mat_A[23][5] * mat_B[5][10] +
                  mat_A[23][6] * mat_B[6][10] +
                  mat_A[23][7] * mat_B[7][10] +
                  mat_A[23][8] * mat_B[8][10] +
                  mat_A[23][9] * mat_B[9][10] +
                  mat_A[23][10] * mat_B[10][10] +
                  mat_A[23][11] * mat_B[11][10] +
                  mat_A[23][12] * mat_B[12][10] +
                  mat_A[23][13] * mat_B[13][10] +
                  mat_A[23][14] * mat_B[14][10] +
                  mat_A[23][15] * mat_B[15][10] +
                  mat_A[23][16] * mat_B[16][10] +
                  mat_A[23][17] * mat_B[17][10] +
                  mat_A[23][18] * mat_B[18][10] +
                  mat_A[23][19] * mat_B[19][10] +
                  mat_A[23][20] * mat_B[20][10] +
                  mat_A[23][21] * mat_B[21][10] +
                  mat_A[23][22] * mat_B[22][10] +
                  mat_A[23][23] * mat_B[23][10] +
                  mat_A[23][24] * mat_B[24][10] +
                  mat_A[23][25] * mat_B[25][10] +
                  mat_A[23][26] * mat_B[26][10] +
                  mat_A[23][27] * mat_B[27][10] +
                  mat_A[23][28] * mat_B[28][10] +
                  mat_A[23][29] * mat_B[29][10] +
                  mat_A[23][30] * mat_B[30][10] +
                  mat_A[23][31] * mat_B[31][10];
    mat_C[23][11] <= 
                  mat_A[23][0] * mat_B[0][11] +
                  mat_A[23][1] * mat_B[1][11] +
                  mat_A[23][2] * mat_B[2][11] +
                  mat_A[23][3] * mat_B[3][11] +
                  mat_A[23][4] * mat_B[4][11] +
                  mat_A[23][5] * mat_B[5][11] +
                  mat_A[23][6] * mat_B[6][11] +
                  mat_A[23][7] * mat_B[7][11] +
                  mat_A[23][8] * mat_B[8][11] +
                  mat_A[23][9] * mat_B[9][11] +
                  mat_A[23][10] * mat_B[10][11] +
                  mat_A[23][11] * mat_B[11][11] +
                  mat_A[23][12] * mat_B[12][11] +
                  mat_A[23][13] * mat_B[13][11] +
                  mat_A[23][14] * mat_B[14][11] +
                  mat_A[23][15] * mat_B[15][11] +
                  mat_A[23][16] * mat_B[16][11] +
                  mat_A[23][17] * mat_B[17][11] +
                  mat_A[23][18] * mat_B[18][11] +
                  mat_A[23][19] * mat_B[19][11] +
                  mat_A[23][20] * mat_B[20][11] +
                  mat_A[23][21] * mat_B[21][11] +
                  mat_A[23][22] * mat_B[22][11] +
                  mat_A[23][23] * mat_B[23][11] +
                  mat_A[23][24] * mat_B[24][11] +
                  mat_A[23][25] * mat_B[25][11] +
                  mat_A[23][26] * mat_B[26][11] +
                  mat_A[23][27] * mat_B[27][11] +
                  mat_A[23][28] * mat_B[28][11] +
                  mat_A[23][29] * mat_B[29][11] +
                  mat_A[23][30] * mat_B[30][11] +
                  mat_A[23][31] * mat_B[31][11];
    mat_C[23][12] <= 
                  mat_A[23][0] * mat_B[0][12] +
                  mat_A[23][1] * mat_B[1][12] +
                  mat_A[23][2] * mat_B[2][12] +
                  mat_A[23][3] * mat_B[3][12] +
                  mat_A[23][4] * mat_B[4][12] +
                  mat_A[23][5] * mat_B[5][12] +
                  mat_A[23][6] * mat_B[6][12] +
                  mat_A[23][7] * mat_B[7][12] +
                  mat_A[23][8] * mat_B[8][12] +
                  mat_A[23][9] * mat_B[9][12] +
                  mat_A[23][10] * mat_B[10][12] +
                  mat_A[23][11] * mat_B[11][12] +
                  mat_A[23][12] * mat_B[12][12] +
                  mat_A[23][13] * mat_B[13][12] +
                  mat_A[23][14] * mat_B[14][12] +
                  mat_A[23][15] * mat_B[15][12] +
                  mat_A[23][16] * mat_B[16][12] +
                  mat_A[23][17] * mat_B[17][12] +
                  mat_A[23][18] * mat_B[18][12] +
                  mat_A[23][19] * mat_B[19][12] +
                  mat_A[23][20] * mat_B[20][12] +
                  mat_A[23][21] * mat_B[21][12] +
                  mat_A[23][22] * mat_B[22][12] +
                  mat_A[23][23] * mat_B[23][12] +
                  mat_A[23][24] * mat_B[24][12] +
                  mat_A[23][25] * mat_B[25][12] +
                  mat_A[23][26] * mat_B[26][12] +
                  mat_A[23][27] * mat_B[27][12] +
                  mat_A[23][28] * mat_B[28][12] +
                  mat_A[23][29] * mat_B[29][12] +
                  mat_A[23][30] * mat_B[30][12] +
                  mat_A[23][31] * mat_B[31][12];
    mat_C[23][13] <= 
                  mat_A[23][0] * mat_B[0][13] +
                  mat_A[23][1] * mat_B[1][13] +
                  mat_A[23][2] * mat_B[2][13] +
                  mat_A[23][3] * mat_B[3][13] +
                  mat_A[23][4] * mat_B[4][13] +
                  mat_A[23][5] * mat_B[5][13] +
                  mat_A[23][6] * mat_B[6][13] +
                  mat_A[23][7] * mat_B[7][13] +
                  mat_A[23][8] * mat_B[8][13] +
                  mat_A[23][9] * mat_B[9][13] +
                  mat_A[23][10] * mat_B[10][13] +
                  mat_A[23][11] * mat_B[11][13] +
                  mat_A[23][12] * mat_B[12][13] +
                  mat_A[23][13] * mat_B[13][13] +
                  mat_A[23][14] * mat_B[14][13] +
                  mat_A[23][15] * mat_B[15][13] +
                  mat_A[23][16] * mat_B[16][13] +
                  mat_A[23][17] * mat_B[17][13] +
                  mat_A[23][18] * mat_B[18][13] +
                  mat_A[23][19] * mat_B[19][13] +
                  mat_A[23][20] * mat_B[20][13] +
                  mat_A[23][21] * mat_B[21][13] +
                  mat_A[23][22] * mat_B[22][13] +
                  mat_A[23][23] * mat_B[23][13] +
                  mat_A[23][24] * mat_B[24][13] +
                  mat_A[23][25] * mat_B[25][13] +
                  mat_A[23][26] * mat_B[26][13] +
                  mat_A[23][27] * mat_B[27][13] +
                  mat_A[23][28] * mat_B[28][13] +
                  mat_A[23][29] * mat_B[29][13] +
                  mat_A[23][30] * mat_B[30][13] +
                  mat_A[23][31] * mat_B[31][13];
    mat_C[23][14] <= 
                  mat_A[23][0] * mat_B[0][14] +
                  mat_A[23][1] * mat_B[1][14] +
                  mat_A[23][2] * mat_B[2][14] +
                  mat_A[23][3] * mat_B[3][14] +
                  mat_A[23][4] * mat_B[4][14] +
                  mat_A[23][5] * mat_B[5][14] +
                  mat_A[23][6] * mat_B[6][14] +
                  mat_A[23][7] * mat_B[7][14] +
                  mat_A[23][8] * mat_B[8][14] +
                  mat_A[23][9] * mat_B[9][14] +
                  mat_A[23][10] * mat_B[10][14] +
                  mat_A[23][11] * mat_B[11][14] +
                  mat_A[23][12] * mat_B[12][14] +
                  mat_A[23][13] * mat_B[13][14] +
                  mat_A[23][14] * mat_B[14][14] +
                  mat_A[23][15] * mat_B[15][14] +
                  mat_A[23][16] * mat_B[16][14] +
                  mat_A[23][17] * mat_B[17][14] +
                  mat_A[23][18] * mat_B[18][14] +
                  mat_A[23][19] * mat_B[19][14] +
                  mat_A[23][20] * mat_B[20][14] +
                  mat_A[23][21] * mat_B[21][14] +
                  mat_A[23][22] * mat_B[22][14] +
                  mat_A[23][23] * mat_B[23][14] +
                  mat_A[23][24] * mat_B[24][14] +
                  mat_A[23][25] * mat_B[25][14] +
                  mat_A[23][26] * mat_B[26][14] +
                  mat_A[23][27] * mat_B[27][14] +
                  mat_A[23][28] * mat_B[28][14] +
                  mat_A[23][29] * mat_B[29][14] +
                  mat_A[23][30] * mat_B[30][14] +
                  mat_A[23][31] * mat_B[31][14];
    mat_C[23][15] <= 
                  mat_A[23][0] * mat_B[0][15] +
                  mat_A[23][1] * mat_B[1][15] +
                  mat_A[23][2] * mat_B[2][15] +
                  mat_A[23][3] * mat_B[3][15] +
                  mat_A[23][4] * mat_B[4][15] +
                  mat_A[23][5] * mat_B[5][15] +
                  mat_A[23][6] * mat_B[6][15] +
                  mat_A[23][7] * mat_B[7][15] +
                  mat_A[23][8] * mat_B[8][15] +
                  mat_A[23][9] * mat_B[9][15] +
                  mat_A[23][10] * mat_B[10][15] +
                  mat_A[23][11] * mat_B[11][15] +
                  mat_A[23][12] * mat_B[12][15] +
                  mat_A[23][13] * mat_B[13][15] +
                  mat_A[23][14] * mat_B[14][15] +
                  mat_A[23][15] * mat_B[15][15] +
                  mat_A[23][16] * mat_B[16][15] +
                  mat_A[23][17] * mat_B[17][15] +
                  mat_A[23][18] * mat_B[18][15] +
                  mat_A[23][19] * mat_B[19][15] +
                  mat_A[23][20] * mat_B[20][15] +
                  mat_A[23][21] * mat_B[21][15] +
                  mat_A[23][22] * mat_B[22][15] +
                  mat_A[23][23] * mat_B[23][15] +
                  mat_A[23][24] * mat_B[24][15] +
                  mat_A[23][25] * mat_B[25][15] +
                  mat_A[23][26] * mat_B[26][15] +
                  mat_A[23][27] * mat_B[27][15] +
                  mat_A[23][28] * mat_B[28][15] +
                  mat_A[23][29] * mat_B[29][15] +
                  mat_A[23][30] * mat_B[30][15] +
                  mat_A[23][31] * mat_B[31][15];
    mat_C[23][16] <= 
                  mat_A[23][0] * mat_B[0][16] +
                  mat_A[23][1] * mat_B[1][16] +
                  mat_A[23][2] * mat_B[2][16] +
                  mat_A[23][3] * mat_B[3][16] +
                  mat_A[23][4] * mat_B[4][16] +
                  mat_A[23][5] * mat_B[5][16] +
                  mat_A[23][6] * mat_B[6][16] +
                  mat_A[23][7] * mat_B[7][16] +
                  mat_A[23][8] * mat_B[8][16] +
                  mat_A[23][9] * mat_B[9][16] +
                  mat_A[23][10] * mat_B[10][16] +
                  mat_A[23][11] * mat_B[11][16] +
                  mat_A[23][12] * mat_B[12][16] +
                  mat_A[23][13] * mat_B[13][16] +
                  mat_A[23][14] * mat_B[14][16] +
                  mat_A[23][15] * mat_B[15][16] +
                  mat_A[23][16] * mat_B[16][16] +
                  mat_A[23][17] * mat_B[17][16] +
                  mat_A[23][18] * mat_B[18][16] +
                  mat_A[23][19] * mat_B[19][16] +
                  mat_A[23][20] * mat_B[20][16] +
                  mat_A[23][21] * mat_B[21][16] +
                  mat_A[23][22] * mat_B[22][16] +
                  mat_A[23][23] * mat_B[23][16] +
                  mat_A[23][24] * mat_B[24][16] +
                  mat_A[23][25] * mat_B[25][16] +
                  mat_A[23][26] * mat_B[26][16] +
                  mat_A[23][27] * mat_B[27][16] +
                  mat_A[23][28] * mat_B[28][16] +
                  mat_A[23][29] * mat_B[29][16] +
                  mat_A[23][30] * mat_B[30][16] +
                  mat_A[23][31] * mat_B[31][16];
    mat_C[23][17] <= 
                  mat_A[23][0] * mat_B[0][17] +
                  mat_A[23][1] * mat_B[1][17] +
                  mat_A[23][2] * mat_B[2][17] +
                  mat_A[23][3] * mat_B[3][17] +
                  mat_A[23][4] * mat_B[4][17] +
                  mat_A[23][5] * mat_B[5][17] +
                  mat_A[23][6] * mat_B[6][17] +
                  mat_A[23][7] * mat_B[7][17] +
                  mat_A[23][8] * mat_B[8][17] +
                  mat_A[23][9] * mat_B[9][17] +
                  mat_A[23][10] * mat_B[10][17] +
                  mat_A[23][11] * mat_B[11][17] +
                  mat_A[23][12] * mat_B[12][17] +
                  mat_A[23][13] * mat_B[13][17] +
                  mat_A[23][14] * mat_B[14][17] +
                  mat_A[23][15] * mat_B[15][17] +
                  mat_A[23][16] * mat_B[16][17] +
                  mat_A[23][17] * mat_B[17][17] +
                  mat_A[23][18] * mat_B[18][17] +
                  mat_A[23][19] * mat_B[19][17] +
                  mat_A[23][20] * mat_B[20][17] +
                  mat_A[23][21] * mat_B[21][17] +
                  mat_A[23][22] * mat_B[22][17] +
                  mat_A[23][23] * mat_B[23][17] +
                  mat_A[23][24] * mat_B[24][17] +
                  mat_A[23][25] * mat_B[25][17] +
                  mat_A[23][26] * mat_B[26][17] +
                  mat_A[23][27] * mat_B[27][17] +
                  mat_A[23][28] * mat_B[28][17] +
                  mat_A[23][29] * mat_B[29][17] +
                  mat_A[23][30] * mat_B[30][17] +
                  mat_A[23][31] * mat_B[31][17];
    mat_C[23][18] <= 
                  mat_A[23][0] * mat_B[0][18] +
                  mat_A[23][1] * mat_B[1][18] +
                  mat_A[23][2] * mat_B[2][18] +
                  mat_A[23][3] * mat_B[3][18] +
                  mat_A[23][4] * mat_B[4][18] +
                  mat_A[23][5] * mat_B[5][18] +
                  mat_A[23][6] * mat_B[6][18] +
                  mat_A[23][7] * mat_B[7][18] +
                  mat_A[23][8] * mat_B[8][18] +
                  mat_A[23][9] * mat_B[9][18] +
                  mat_A[23][10] * mat_B[10][18] +
                  mat_A[23][11] * mat_B[11][18] +
                  mat_A[23][12] * mat_B[12][18] +
                  mat_A[23][13] * mat_B[13][18] +
                  mat_A[23][14] * mat_B[14][18] +
                  mat_A[23][15] * mat_B[15][18] +
                  mat_A[23][16] * mat_B[16][18] +
                  mat_A[23][17] * mat_B[17][18] +
                  mat_A[23][18] * mat_B[18][18] +
                  mat_A[23][19] * mat_B[19][18] +
                  mat_A[23][20] * mat_B[20][18] +
                  mat_A[23][21] * mat_B[21][18] +
                  mat_A[23][22] * mat_B[22][18] +
                  mat_A[23][23] * mat_B[23][18] +
                  mat_A[23][24] * mat_B[24][18] +
                  mat_A[23][25] * mat_B[25][18] +
                  mat_A[23][26] * mat_B[26][18] +
                  mat_A[23][27] * mat_B[27][18] +
                  mat_A[23][28] * mat_B[28][18] +
                  mat_A[23][29] * mat_B[29][18] +
                  mat_A[23][30] * mat_B[30][18] +
                  mat_A[23][31] * mat_B[31][18];
    mat_C[23][19] <= 
                  mat_A[23][0] * mat_B[0][19] +
                  mat_A[23][1] * mat_B[1][19] +
                  mat_A[23][2] * mat_B[2][19] +
                  mat_A[23][3] * mat_B[3][19] +
                  mat_A[23][4] * mat_B[4][19] +
                  mat_A[23][5] * mat_B[5][19] +
                  mat_A[23][6] * mat_B[6][19] +
                  mat_A[23][7] * mat_B[7][19] +
                  mat_A[23][8] * mat_B[8][19] +
                  mat_A[23][9] * mat_B[9][19] +
                  mat_A[23][10] * mat_B[10][19] +
                  mat_A[23][11] * mat_B[11][19] +
                  mat_A[23][12] * mat_B[12][19] +
                  mat_A[23][13] * mat_B[13][19] +
                  mat_A[23][14] * mat_B[14][19] +
                  mat_A[23][15] * mat_B[15][19] +
                  mat_A[23][16] * mat_B[16][19] +
                  mat_A[23][17] * mat_B[17][19] +
                  mat_A[23][18] * mat_B[18][19] +
                  mat_A[23][19] * mat_B[19][19] +
                  mat_A[23][20] * mat_B[20][19] +
                  mat_A[23][21] * mat_B[21][19] +
                  mat_A[23][22] * mat_B[22][19] +
                  mat_A[23][23] * mat_B[23][19] +
                  mat_A[23][24] * mat_B[24][19] +
                  mat_A[23][25] * mat_B[25][19] +
                  mat_A[23][26] * mat_B[26][19] +
                  mat_A[23][27] * mat_B[27][19] +
                  mat_A[23][28] * mat_B[28][19] +
                  mat_A[23][29] * mat_B[29][19] +
                  mat_A[23][30] * mat_B[30][19] +
                  mat_A[23][31] * mat_B[31][19];
    mat_C[23][20] <= 
                  mat_A[23][0] * mat_B[0][20] +
                  mat_A[23][1] * mat_B[1][20] +
                  mat_A[23][2] * mat_B[2][20] +
                  mat_A[23][3] * mat_B[3][20] +
                  mat_A[23][4] * mat_B[4][20] +
                  mat_A[23][5] * mat_B[5][20] +
                  mat_A[23][6] * mat_B[6][20] +
                  mat_A[23][7] * mat_B[7][20] +
                  mat_A[23][8] * mat_B[8][20] +
                  mat_A[23][9] * mat_B[9][20] +
                  mat_A[23][10] * mat_B[10][20] +
                  mat_A[23][11] * mat_B[11][20] +
                  mat_A[23][12] * mat_B[12][20] +
                  mat_A[23][13] * mat_B[13][20] +
                  mat_A[23][14] * mat_B[14][20] +
                  mat_A[23][15] * mat_B[15][20] +
                  mat_A[23][16] * mat_B[16][20] +
                  mat_A[23][17] * mat_B[17][20] +
                  mat_A[23][18] * mat_B[18][20] +
                  mat_A[23][19] * mat_B[19][20] +
                  mat_A[23][20] * mat_B[20][20] +
                  mat_A[23][21] * mat_B[21][20] +
                  mat_A[23][22] * mat_B[22][20] +
                  mat_A[23][23] * mat_B[23][20] +
                  mat_A[23][24] * mat_B[24][20] +
                  mat_A[23][25] * mat_B[25][20] +
                  mat_A[23][26] * mat_B[26][20] +
                  mat_A[23][27] * mat_B[27][20] +
                  mat_A[23][28] * mat_B[28][20] +
                  mat_A[23][29] * mat_B[29][20] +
                  mat_A[23][30] * mat_B[30][20] +
                  mat_A[23][31] * mat_B[31][20];
    mat_C[23][21] <= 
                  mat_A[23][0] * mat_B[0][21] +
                  mat_A[23][1] * mat_B[1][21] +
                  mat_A[23][2] * mat_B[2][21] +
                  mat_A[23][3] * mat_B[3][21] +
                  mat_A[23][4] * mat_B[4][21] +
                  mat_A[23][5] * mat_B[5][21] +
                  mat_A[23][6] * mat_B[6][21] +
                  mat_A[23][7] * mat_B[7][21] +
                  mat_A[23][8] * mat_B[8][21] +
                  mat_A[23][9] * mat_B[9][21] +
                  mat_A[23][10] * mat_B[10][21] +
                  mat_A[23][11] * mat_B[11][21] +
                  mat_A[23][12] * mat_B[12][21] +
                  mat_A[23][13] * mat_B[13][21] +
                  mat_A[23][14] * mat_B[14][21] +
                  mat_A[23][15] * mat_B[15][21] +
                  mat_A[23][16] * mat_B[16][21] +
                  mat_A[23][17] * mat_B[17][21] +
                  mat_A[23][18] * mat_B[18][21] +
                  mat_A[23][19] * mat_B[19][21] +
                  mat_A[23][20] * mat_B[20][21] +
                  mat_A[23][21] * mat_B[21][21] +
                  mat_A[23][22] * mat_B[22][21] +
                  mat_A[23][23] * mat_B[23][21] +
                  mat_A[23][24] * mat_B[24][21] +
                  mat_A[23][25] * mat_B[25][21] +
                  mat_A[23][26] * mat_B[26][21] +
                  mat_A[23][27] * mat_B[27][21] +
                  mat_A[23][28] * mat_B[28][21] +
                  mat_A[23][29] * mat_B[29][21] +
                  mat_A[23][30] * mat_B[30][21] +
                  mat_A[23][31] * mat_B[31][21];
    mat_C[23][22] <= 
                  mat_A[23][0] * mat_B[0][22] +
                  mat_A[23][1] * mat_B[1][22] +
                  mat_A[23][2] * mat_B[2][22] +
                  mat_A[23][3] * mat_B[3][22] +
                  mat_A[23][4] * mat_B[4][22] +
                  mat_A[23][5] * mat_B[5][22] +
                  mat_A[23][6] * mat_B[6][22] +
                  mat_A[23][7] * mat_B[7][22] +
                  mat_A[23][8] * mat_B[8][22] +
                  mat_A[23][9] * mat_B[9][22] +
                  mat_A[23][10] * mat_B[10][22] +
                  mat_A[23][11] * mat_B[11][22] +
                  mat_A[23][12] * mat_B[12][22] +
                  mat_A[23][13] * mat_B[13][22] +
                  mat_A[23][14] * mat_B[14][22] +
                  mat_A[23][15] * mat_B[15][22] +
                  mat_A[23][16] * mat_B[16][22] +
                  mat_A[23][17] * mat_B[17][22] +
                  mat_A[23][18] * mat_B[18][22] +
                  mat_A[23][19] * mat_B[19][22] +
                  mat_A[23][20] * mat_B[20][22] +
                  mat_A[23][21] * mat_B[21][22] +
                  mat_A[23][22] * mat_B[22][22] +
                  mat_A[23][23] * mat_B[23][22] +
                  mat_A[23][24] * mat_B[24][22] +
                  mat_A[23][25] * mat_B[25][22] +
                  mat_A[23][26] * mat_B[26][22] +
                  mat_A[23][27] * mat_B[27][22] +
                  mat_A[23][28] * mat_B[28][22] +
                  mat_A[23][29] * mat_B[29][22] +
                  mat_A[23][30] * mat_B[30][22] +
                  mat_A[23][31] * mat_B[31][22];
    mat_C[23][23] <= 
                  mat_A[23][0] * mat_B[0][23] +
                  mat_A[23][1] * mat_B[1][23] +
                  mat_A[23][2] * mat_B[2][23] +
                  mat_A[23][3] * mat_B[3][23] +
                  mat_A[23][4] * mat_B[4][23] +
                  mat_A[23][5] * mat_B[5][23] +
                  mat_A[23][6] * mat_B[6][23] +
                  mat_A[23][7] * mat_B[7][23] +
                  mat_A[23][8] * mat_B[8][23] +
                  mat_A[23][9] * mat_B[9][23] +
                  mat_A[23][10] * mat_B[10][23] +
                  mat_A[23][11] * mat_B[11][23] +
                  mat_A[23][12] * mat_B[12][23] +
                  mat_A[23][13] * mat_B[13][23] +
                  mat_A[23][14] * mat_B[14][23] +
                  mat_A[23][15] * mat_B[15][23] +
                  mat_A[23][16] * mat_B[16][23] +
                  mat_A[23][17] * mat_B[17][23] +
                  mat_A[23][18] * mat_B[18][23] +
                  mat_A[23][19] * mat_B[19][23] +
                  mat_A[23][20] * mat_B[20][23] +
                  mat_A[23][21] * mat_B[21][23] +
                  mat_A[23][22] * mat_B[22][23] +
                  mat_A[23][23] * mat_B[23][23] +
                  mat_A[23][24] * mat_B[24][23] +
                  mat_A[23][25] * mat_B[25][23] +
                  mat_A[23][26] * mat_B[26][23] +
                  mat_A[23][27] * mat_B[27][23] +
                  mat_A[23][28] * mat_B[28][23] +
                  mat_A[23][29] * mat_B[29][23] +
                  mat_A[23][30] * mat_B[30][23] +
                  mat_A[23][31] * mat_B[31][23];
    mat_C[23][24] <= 
                  mat_A[23][0] * mat_B[0][24] +
                  mat_A[23][1] * mat_B[1][24] +
                  mat_A[23][2] * mat_B[2][24] +
                  mat_A[23][3] * mat_B[3][24] +
                  mat_A[23][4] * mat_B[4][24] +
                  mat_A[23][5] * mat_B[5][24] +
                  mat_A[23][6] * mat_B[6][24] +
                  mat_A[23][7] * mat_B[7][24] +
                  mat_A[23][8] * mat_B[8][24] +
                  mat_A[23][9] * mat_B[9][24] +
                  mat_A[23][10] * mat_B[10][24] +
                  mat_A[23][11] * mat_B[11][24] +
                  mat_A[23][12] * mat_B[12][24] +
                  mat_A[23][13] * mat_B[13][24] +
                  mat_A[23][14] * mat_B[14][24] +
                  mat_A[23][15] * mat_B[15][24] +
                  mat_A[23][16] * mat_B[16][24] +
                  mat_A[23][17] * mat_B[17][24] +
                  mat_A[23][18] * mat_B[18][24] +
                  mat_A[23][19] * mat_B[19][24] +
                  mat_A[23][20] * mat_B[20][24] +
                  mat_A[23][21] * mat_B[21][24] +
                  mat_A[23][22] * mat_B[22][24] +
                  mat_A[23][23] * mat_B[23][24] +
                  mat_A[23][24] * mat_B[24][24] +
                  mat_A[23][25] * mat_B[25][24] +
                  mat_A[23][26] * mat_B[26][24] +
                  mat_A[23][27] * mat_B[27][24] +
                  mat_A[23][28] * mat_B[28][24] +
                  mat_A[23][29] * mat_B[29][24] +
                  mat_A[23][30] * mat_B[30][24] +
                  mat_A[23][31] * mat_B[31][24];
    mat_C[23][25] <= 
                  mat_A[23][0] * mat_B[0][25] +
                  mat_A[23][1] * mat_B[1][25] +
                  mat_A[23][2] * mat_B[2][25] +
                  mat_A[23][3] * mat_B[3][25] +
                  mat_A[23][4] * mat_B[4][25] +
                  mat_A[23][5] * mat_B[5][25] +
                  mat_A[23][6] * mat_B[6][25] +
                  mat_A[23][7] * mat_B[7][25] +
                  mat_A[23][8] * mat_B[8][25] +
                  mat_A[23][9] * mat_B[9][25] +
                  mat_A[23][10] * mat_B[10][25] +
                  mat_A[23][11] * mat_B[11][25] +
                  mat_A[23][12] * mat_B[12][25] +
                  mat_A[23][13] * mat_B[13][25] +
                  mat_A[23][14] * mat_B[14][25] +
                  mat_A[23][15] * mat_B[15][25] +
                  mat_A[23][16] * mat_B[16][25] +
                  mat_A[23][17] * mat_B[17][25] +
                  mat_A[23][18] * mat_B[18][25] +
                  mat_A[23][19] * mat_B[19][25] +
                  mat_A[23][20] * mat_B[20][25] +
                  mat_A[23][21] * mat_B[21][25] +
                  mat_A[23][22] * mat_B[22][25] +
                  mat_A[23][23] * mat_B[23][25] +
                  mat_A[23][24] * mat_B[24][25] +
                  mat_A[23][25] * mat_B[25][25] +
                  mat_A[23][26] * mat_B[26][25] +
                  mat_A[23][27] * mat_B[27][25] +
                  mat_A[23][28] * mat_B[28][25] +
                  mat_A[23][29] * mat_B[29][25] +
                  mat_A[23][30] * mat_B[30][25] +
                  mat_A[23][31] * mat_B[31][25];
    mat_C[23][26] <= 
                  mat_A[23][0] * mat_B[0][26] +
                  mat_A[23][1] * mat_B[1][26] +
                  mat_A[23][2] * mat_B[2][26] +
                  mat_A[23][3] * mat_B[3][26] +
                  mat_A[23][4] * mat_B[4][26] +
                  mat_A[23][5] * mat_B[5][26] +
                  mat_A[23][6] * mat_B[6][26] +
                  mat_A[23][7] * mat_B[7][26] +
                  mat_A[23][8] * mat_B[8][26] +
                  mat_A[23][9] * mat_B[9][26] +
                  mat_A[23][10] * mat_B[10][26] +
                  mat_A[23][11] * mat_B[11][26] +
                  mat_A[23][12] * mat_B[12][26] +
                  mat_A[23][13] * mat_B[13][26] +
                  mat_A[23][14] * mat_B[14][26] +
                  mat_A[23][15] * mat_B[15][26] +
                  mat_A[23][16] * mat_B[16][26] +
                  mat_A[23][17] * mat_B[17][26] +
                  mat_A[23][18] * mat_B[18][26] +
                  mat_A[23][19] * mat_B[19][26] +
                  mat_A[23][20] * mat_B[20][26] +
                  mat_A[23][21] * mat_B[21][26] +
                  mat_A[23][22] * mat_B[22][26] +
                  mat_A[23][23] * mat_B[23][26] +
                  mat_A[23][24] * mat_B[24][26] +
                  mat_A[23][25] * mat_B[25][26] +
                  mat_A[23][26] * mat_B[26][26] +
                  mat_A[23][27] * mat_B[27][26] +
                  mat_A[23][28] * mat_B[28][26] +
                  mat_A[23][29] * mat_B[29][26] +
                  mat_A[23][30] * mat_B[30][26] +
                  mat_A[23][31] * mat_B[31][26];
    mat_C[23][27] <= 
                  mat_A[23][0] * mat_B[0][27] +
                  mat_A[23][1] * mat_B[1][27] +
                  mat_A[23][2] * mat_B[2][27] +
                  mat_A[23][3] * mat_B[3][27] +
                  mat_A[23][4] * mat_B[4][27] +
                  mat_A[23][5] * mat_B[5][27] +
                  mat_A[23][6] * mat_B[6][27] +
                  mat_A[23][7] * mat_B[7][27] +
                  mat_A[23][8] * mat_B[8][27] +
                  mat_A[23][9] * mat_B[9][27] +
                  mat_A[23][10] * mat_B[10][27] +
                  mat_A[23][11] * mat_B[11][27] +
                  mat_A[23][12] * mat_B[12][27] +
                  mat_A[23][13] * mat_B[13][27] +
                  mat_A[23][14] * mat_B[14][27] +
                  mat_A[23][15] * mat_B[15][27] +
                  mat_A[23][16] * mat_B[16][27] +
                  mat_A[23][17] * mat_B[17][27] +
                  mat_A[23][18] * mat_B[18][27] +
                  mat_A[23][19] * mat_B[19][27] +
                  mat_A[23][20] * mat_B[20][27] +
                  mat_A[23][21] * mat_B[21][27] +
                  mat_A[23][22] * mat_B[22][27] +
                  mat_A[23][23] * mat_B[23][27] +
                  mat_A[23][24] * mat_B[24][27] +
                  mat_A[23][25] * mat_B[25][27] +
                  mat_A[23][26] * mat_B[26][27] +
                  mat_A[23][27] * mat_B[27][27] +
                  mat_A[23][28] * mat_B[28][27] +
                  mat_A[23][29] * mat_B[29][27] +
                  mat_A[23][30] * mat_B[30][27] +
                  mat_A[23][31] * mat_B[31][27];
    mat_C[23][28] <= 
                  mat_A[23][0] * mat_B[0][28] +
                  mat_A[23][1] * mat_B[1][28] +
                  mat_A[23][2] * mat_B[2][28] +
                  mat_A[23][3] * mat_B[3][28] +
                  mat_A[23][4] * mat_B[4][28] +
                  mat_A[23][5] * mat_B[5][28] +
                  mat_A[23][6] * mat_B[6][28] +
                  mat_A[23][7] * mat_B[7][28] +
                  mat_A[23][8] * mat_B[8][28] +
                  mat_A[23][9] * mat_B[9][28] +
                  mat_A[23][10] * mat_B[10][28] +
                  mat_A[23][11] * mat_B[11][28] +
                  mat_A[23][12] * mat_B[12][28] +
                  mat_A[23][13] * mat_B[13][28] +
                  mat_A[23][14] * mat_B[14][28] +
                  mat_A[23][15] * mat_B[15][28] +
                  mat_A[23][16] * mat_B[16][28] +
                  mat_A[23][17] * mat_B[17][28] +
                  mat_A[23][18] * mat_B[18][28] +
                  mat_A[23][19] * mat_B[19][28] +
                  mat_A[23][20] * mat_B[20][28] +
                  mat_A[23][21] * mat_B[21][28] +
                  mat_A[23][22] * mat_B[22][28] +
                  mat_A[23][23] * mat_B[23][28] +
                  mat_A[23][24] * mat_B[24][28] +
                  mat_A[23][25] * mat_B[25][28] +
                  mat_A[23][26] * mat_B[26][28] +
                  mat_A[23][27] * mat_B[27][28] +
                  mat_A[23][28] * mat_B[28][28] +
                  mat_A[23][29] * mat_B[29][28] +
                  mat_A[23][30] * mat_B[30][28] +
                  mat_A[23][31] * mat_B[31][28];
    mat_C[23][29] <= 
                  mat_A[23][0] * mat_B[0][29] +
                  mat_A[23][1] * mat_B[1][29] +
                  mat_A[23][2] * mat_B[2][29] +
                  mat_A[23][3] * mat_B[3][29] +
                  mat_A[23][4] * mat_B[4][29] +
                  mat_A[23][5] * mat_B[5][29] +
                  mat_A[23][6] * mat_B[6][29] +
                  mat_A[23][7] * mat_B[7][29] +
                  mat_A[23][8] * mat_B[8][29] +
                  mat_A[23][9] * mat_B[9][29] +
                  mat_A[23][10] * mat_B[10][29] +
                  mat_A[23][11] * mat_B[11][29] +
                  mat_A[23][12] * mat_B[12][29] +
                  mat_A[23][13] * mat_B[13][29] +
                  mat_A[23][14] * mat_B[14][29] +
                  mat_A[23][15] * mat_B[15][29] +
                  mat_A[23][16] * mat_B[16][29] +
                  mat_A[23][17] * mat_B[17][29] +
                  mat_A[23][18] * mat_B[18][29] +
                  mat_A[23][19] * mat_B[19][29] +
                  mat_A[23][20] * mat_B[20][29] +
                  mat_A[23][21] * mat_B[21][29] +
                  mat_A[23][22] * mat_B[22][29] +
                  mat_A[23][23] * mat_B[23][29] +
                  mat_A[23][24] * mat_B[24][29] +
                  mat_A[23][25] * mat_B[25][29] +
                  mat_A[23][26] * mat_B[26][29] +
                  mat_A[23][27] * mat_B[27][29] +
                  mat_A[23][28] * mat_B[28][29] +
                  mat_A[23][29] * mat_B[29][29] +
                  mat_A[23][30] * mat_B[30][29] +
                  mat_A[23][31] * mat_B[31][29];
    mat_C[23][30] <= 
                  mat_A[23][0] * mat_B[0][30] +
                  mat_A[23][1] * mat_B[1][30] +
                  mat_A[23][2] * mat_B[2][30] +
                  mat_A[23][3] * mat_B[3][30] +
                  mat_A[23][4] * mat_B[4][30] +
                  mat_A[23][5] * mat_B[5][30] +
                  mat_A[23][6] * mat_B[6][30] +
                  mat_A[23][7] * mat_B[7][30] +
                  mat_A[23][8] * mat_B[8][30] +
                  mat_A[23][9] * mat_B[9][30] +
                  mat_A[23][10] * mat_B[10][30] +
                  mat_A[23][11] * mat_B[11][30] +
                  mat_A[23][12] * mat_B[12][30] +
                  mat_A[23][13] * mat_B[13][30] +
                  mat_A[23][14] * mat_B[14][30] +
                  mat_A[23][15] * mat_B[15][30] +
                  mat_A[23][16] * mat_B[16][30] +
                  mat_A[23][17] * mat_B[17][30] +
                  mat_A[23][18] * mat_B[18][30] +
                  mat_A[23][19] * mat_B[19][30] +
                  mat_A[23][20] * mat_B[20][30] +
                  mat_A[23][21] * mat_B[21][30] +
                  mat_A[23][22] * mat_B[22][30] +
                  mat_A[23][23] * mat_B[23][30] +
                  mat_A[23][24] * mat_B[24][30] +
                  mat_A[23][25] * mat_B[25][30] +
                  mat_A[23][26] * mat_B[26][30] +
                  mat_A[23][27] * mat_B[27][30] +
                  mat_A[23][28] * mat_B[28][30] +
                  mat_A[23][29] * mat_B[29][30] +
                  mat_A[23][30] * mat_B[30][30] +
                  mat_A[23][31] * mat_B[31][30];
    mat_C[23][31] <= 
                  mat_A[23][0] * mat_B[0][31] +
                  mat_A[23][1] * mat_B[1][31] +
                  mat_A[23][2] * mat_B[2][31] +
                  mat_A[23][3] * mat_B[3][31] +
                  mat_A[23][4] * mat_B[4][31] +
                  mat_A[23][5] * mat_B[5][31] +
                  mat_A[23][6] * mat_B[6][31] +
                  mat_A[23][7] * mat_B[7][31] +
                  mat_A[23][8] * mat_B[8][31] +
                  mat_A[23][9] * mat_B[9][31] +
                  mat_A[23][10] * mat_B[10][31] +
                  mat_A[23][11] * mat_B[11][31] +
                  mat_A[23][12] * mat_B[12][31] +
                  mat_A[23][13] * mat_B[13][31] +
                  mat_A[23][14] * mat_B[14][31] +
                  mat_A[23][15] * mat_B[15][31] +
                  mat_A[23][16] * mat_B[16][31] +
                  mat_A[23][17] * mat_B[17][31] +
                  mat_A[23][18] * mat_B[18][31] +
                  mat_A[23][19] * mat_B[19][31] +
                  mat_A[23][20] * mat_B[20][31] +
                  mat_A[23][21] * mat_B[21][31] +
                  mat_A[23][22] * mat_B[22][31] +
                  mat_A[23][23] * mat_B[23][31] +
                  mat_A[23][24] * mat_B[24][31] +
                  mat_A[23][25] * mat_B[25][31] +
                  mat_A[23][26] * mat_B[26][31] +
                  mat_A[23][27] * mat_B[27][31] +
                  mat_A[23][28] * mat_B[28][31] +
                  mat_A[23][29] * mat_B[29][31] +
                  mat_A[23][30] * mat_B[30][31] +
                  mat_A[23][31] * mat_B[31][31];
    mat_C[24][0] <= 
                  mat_A[24][0] * mat_B[0][0] +
                  mat_A[24][1] * mat_B[1][0] +
                  mat_A[24][2] * mat_B[2][0] +
                  mat_A[24][3] * mat_B[3][0] +
                  mat_A[24][4] * mat_B[4][0] +
                  mat_A[24][5] * mat_B[5][0] +
                  mat_A[24][6] * mat_B[6][0] +
                  mat_A[24][7] * mat_B[7][0] +
                  mat_A[24][8] * mat_B[8][0] +
                  mat_A[24][9] * mat_B[9][0] +
                  mat_A[24][10] * mat_B[10][0] +
                  mat_A[24][11] * mat_B[11][0] +
                  mat_A[24][12] * mat_B[12][0] +
                  mat_A[24][13] * mat_B[13][0] +
                  mat_A[24][14] * mat_B[14][0] +
                  mat_A[24][15] * mat_B[15][0] +
                  mat_A[24][16] * mat_B[16][0] +
                  mat_A[24][17] * mat_B[17][0] +
                  mat_A[24][18] * mat_B[18][0] +
                  mat_A[24][19] * mat_B[19][0] +
                  mat_A[24][20] * mat_B[20][0] +
                  mat_A[24][21] * mat_B[21][0] +
                  mat_A[24][22] * mat_B[22][0] +
                  mat_A[24][23] * mat_B[23][0] +
                  mat_A[24][24] * mat_B[24][0] +
                  mat_A[24][25] * mat_B[25][0] +
                  mat_A[24][26] * mat_B[26][0] +
                  mat_A[24][27] * mat_B[27][0] +
                  mat_A[24][28] * mat_B[28][0] +
                  mat_A[24][29] * mat_B[29][0] +
                  mat_A[24][30] * mat_B[30][0] +
                  mat_A[24][31] * mat_B[31][0];
    mat_C[24][1] <= 
                  mat_A[24][0] * mat_B[0][1] +
                  mat_A[24][1] * mat_B[1][1] +
                  mat_A[24][2] * mat_B[2][1] +
                  mat_A[24][3] * mat_B[3][1] +
                  mat_A[24][4] * mat_B[4][1] +
                  mat_A[24][5] * mat_B[5][1] +
                  mat_A[24][6] * mat_B[6][1] +
                  mat_A[24][7] * mat_B[7][1] +
                  mat_A[24][8] * mat_B[8][1] +
                  mat_A[24][9] * mat_B[9][1] +
                  mat_A[24][10] * mat_B[10][1] +
                  mat_A[24][11] * mat_B[11][1] +
                  mat_A[24][12] * mat_B[12][1] +
                  mat_A[24][13] * mat_B[13][1] +
                  mat_A[24][14] * mat_B[14][1] +
                  mat_A[24][15] * mat_B[15][1] +
                  mat_A[24][16] * mat_B[16][1] +
                  mat_A[24][17] * mat_B[17][1] +
                  mat_A[24][18] * mat_B[18][1] +
                  mat_A[24][19] * mat_B[19][1] +
                  mat_A[24][20] * mat_B[20][1] +
                  mat_A[24][21] * mat_B[21][1] +
                  mat_A[24][22] * mat_B[22][1] +
                  mat_A[24][23] * mat_B[23][1] +
                  mat_A[24][24] * mat_B[24][1] +
                  mat_A[24][25] * mat_B[25][1] +
                  mat_A[24][26] * mat_B[26][1] +
                  mat_A[24][27] * mat_B[27][1] +
                  mat_A[24][28] * mat_B[28][1] +
                  mat_A[24][29] * mat_B[29][1] +
                  mat_A[24][30] * mat_B[30][1] +
                  mat_A[24][31] * mat_B[31][1];
    mat_C[24][2] <= 
                  mat_A[24][0] * mat_B[0][2] +
                  mat_A[24][1] * mat_B[1][2] +
                  mat_A[24][2] * mat_B[2][2] +
                  mat_A[24][3] * mat_B[3][2] +
                  mat_A[24][4] * mat_B[4][2] +
                  mat_A[24][5] * mat_B[5][2] +
                  mat_A[24][6] * mat_B[6][2] +
                  mat_A[24][7] * mat_B[7][2] +
                  mat_A[24][8] * mat_B[8][2] +
                  mat_A[24][9] * mat_B[9][2] +
                  mat_A[24][10] * mat_B[10][2] +
                  mat_A[24][11] * mat_B[11][2] +
                  mat_A[24][12] * mat_B[12][2] +
                  mat_A[24][13] * mat_B[13][2] +
                  mat_A[24][14] * mat_B[14][2] +
                  mat_A[24][15] * mat_B[15][2] +
                  mat_A[24][16] * mat_B[16][2] +
                  mat_A[24][17] * mat_B[17][2] +
                  mat_A[24][18] * mat_B[18][2] +
                  mat_A[24][19] * mat_B[19][2] +
                  mat_A[24][20] * mat_B[20][2] +
                  mat_A[24][21] * mat_B[21][2] +
                  mat_A[24][22] * mat_B[22][2] +
                  mat_A[24][23] * mat_B[23][2] +
                  mat_A[24][24] * mat_B[24][2] +
                  mat_A[24][25] * mat_B[25][2] +
                  mat_A[24][26] * mat_B[26][2] +
                  mat_A[24][27] * mat_B[27][2] +
                  mat_A[24][28] * mat_B[28][2] +
                  mat_A[24][29] * mat_B[29][2] +
                  mat_A[24][30] * mat_B[30][2] +
                  mat_A[24][31] * mat_B[31][2];
    mat_C[24][3] <= 
                  mat_A[24][0] * mat_B[0][3] +
                  mat_A[24][1] * mat_B[1][3] +
                  mat_A[24][2] * mat_B[2][3] +
                  mat_A[24][3] * mat_B[3][3] +
                  mat_A[24][4] * mat_B[4][3] +
                  mat_A[24][5] * mat_B[5][3] +
                  mat_A[24][6] * mat_B[6][3] +
                  mat_A[24][7] * mat_B[7][3] +
                  mat_A[24][8] * mat_B[8][3] +
                  mat_A[24][9] * mat_B[9][3] +
                  mat_A[24][10] * mat_B[10][3] +
                  mat_A[24][11] * mat_B[11][3] +
                  mat_A[24][12] * mat_B[12][3] +
                  mat_A[24][13] * mat_B[13][3] +
                  mat_A[24][14] * mat_B[14][3] +
                  mat_A[24][15] * mat_B[15][3] +
                  mat_A[24][16] * mat_B[16][3] +
                  mat_A[24][17] * mat_B[17][3] +
                  mat_A[24][18] * mat_B[18][3] +
                  mat_A[24][19] * mat_B[19][3] +
                  mat_A[24][20] * mat_B[20][3] +
                  mat_A[24][21] * mat_B[21][3] +
                  mat_A[24][22] * mat_B[22][3] +
                  mat_A[24][23] * mat_B[23][3] +
                  mat_A[24][24] * mat_B[24][3] +
                  mat_A[24][25] * mat_B[25][3] +
                  mat_A[24][26] * mat_B[26][3] +
                  mat_A[24][27] * mat_B[27][3] +
                  mat_A[24][28] * mat_B[28][3] +
                  mat_A[24][29] * mat_B[29][3] +
                  mat_A[24][30] * mat_B[30][3] +
                  mat_A[24][31] * mat_B[31][3];
    mat_C[24][4] <= 
                  mat_A[24][0] * mat_B[0][4] +
                  mat_A[24][1] * mat_B[1][4] +
                  mat_A[24][2] * mat_B[2][4] +
                  mat_A[24][3] * mat_B[3][4] +
                  mat_A[24][4] * mat_B[4][4] +
                  mat_A[24][5] * mat_B[5][4] +
                  mat_A[24][6] * mat_B[6][4] +
                  mat_A[24][7] * mat_B[7][4] +
                  mat_A[24][8] * mat_B[8][4] +
                  mat_A[24][9] * mat_B[9][4] +
                  mat_A[24][10] * mat_B[10][4] +
                  mat_A[24][11] * mat_B[11][4] +
                  mat_A[24][12] * mat_B[12][4] +
                  mat_A[24][13] * mat_B[13][4] +
                  mat_A[24][14] * mat_B[14][4] +
                  mat_A[24][15] * mat_B[15][4] +
                  mat_A[24][16] * mat_B[16][4] +
                  mat_A[24][17] * mat_B[17][4] +
                  mat_A[24][18] * mat_B[18][4] +
                  mat_A[24][19] * mat_B[19][4] +
                  mat_A[24][20] * mat_B[20][4] +
                  mat_A[24][21] * mat_B[21][4] +
                  mat_A[24][22] * mat_B[22][4] +
                  mat_A[24][23] * mat_B[23][4] +
                  mat_A[24][24] * mat_B[24][4] +
                  mat_A[24][25] * mat_B[25][4] +
                  mat_A[24][26] * mat_B[26][4] +
                  mat_A[24][27] * mat_B[27][4] +
                  mat_A[24][28] * mat_B[28][4] +
                  mat_A[24][29] * mat_B[29][4] +
                  mat_A[24][30] * mat_B[30][4] +
                  mat_A[24][31] * mat_B[31][4];
    mat_C[24][5] <= 
                  mat_A[24][0] * mat_B[0][5] +
                  mat_A[24][1] * mat_B[1][5] +
                  mat_A[24][2] * mat_B[2][5] +
                  mat_A[24][3] * mat_B[3][5] +
                  mat_A[24][4] * mat_B[4][5] +
                  mat_A[24][5] * mat_B[5][5] +
                  mat_A[24][6] * mat_B[6][5] +
                  mat_A[24][7] * mat_B[7][5] +
                  mat_A[24][8] * mat_B[8][5] +
                  mat_A[24][9] * mat_B[9][5] +
                  mat_A[24][10] * mat_B[10][5] +
                  mat_A[24][11] * mat_B[11][5] +
                  mat_A[24][12] * mat_B[12][5] +
                  mat_A[24][13] * mat_B[13][5] +
                  mat_A[24][14] * mat_B[14][5] +
                  mat_A[24][15] * mat_B[15][5] +
                  mat_A[24][16] * mat_B[16][5] +
                  mat_A[24][17] * mat_B[17][5] +
                  mat_A[24][18] * mat_B[18][5] +
                  mat_A[24][19] * mat_B[19][5] +
                  mat_A[24][20] * mat_B[20][5] +
                  mat_A[24][21] * mat_B[21][5] +
                  mat_A[24][22] * mat_B[22][5] +
                  mat_A[24][23] * mat_B[23][5] +
                  mat_A[24][24] * mat_B[24][5] +
                  mat_A[24][25] * mat_B[25][5] +
                  mat_A[24][26] * mat_B[26][5] +
                  mat_A[24][27] * mat_B[27][5] +
                  mat_A[24][28] * mat_B[28][5] +
                  mat_A[24][29] * mat_B[29][5] +
                  mat_A[24][30] * mat_B[30][5] +
                  mat_A[24][31] * mat_B[31][5];
    mat_C[24][6] <= 
                  mat_A[24][0] * mat_B[0][6] +
                  mat_A[24][1] * mat_B[1][6] +
                  mat_A[24][2] * mat_B[2][6] +
                  mat_A[24][3] * mat_B[3][6] +
                  mat_A[24][4] * mat_B[4][6] +
                  mat_A[24][5] * mat_B[5][6] +
                  mat_A[24][6] * mat_B[6][6] +
                  mat_A[24][7] * mat_B[7][6] +
                  mat_A[24][8] * mat_B[8][6] +
                  mat_A[24][9] * mat_B[9][6] +
                  mat_A[24][10] * mat_B[10][6] +
                  mat_A[24][11] * mat_B[11][6] +
                  mat_A[24][12] * mat_B[12][6] +
                  mat_A[24][13] * mat_B[13][6] +
                  mat_A[24][14] * mat_B[14][6] +
                  mat_A[24][15] * mat_B[15][6] +
                  mat_A[24][16] * mat_B[16][6] +
                  mat_A[24][17] * mat_B[17][6] +
                  mat_A[24][18] * mat_B[18][6] +
                  mat_A[24][19] * mat_B[19][6] +
                  mat_A[24][20] * mat_B[20][6] +
                  mat_A[24][21] * mat_B[21][6] +
                  mat_A[24][22] * mat_B[22][6] +
                  mat_A[24][23] * mat_B[23][6] +
                  mat_A[24][24] * mat_B[24][6] +
                  mat_A[24][25] * mat_B[25][6] +
                  mat_A[24][26] * mat_B[26][6] +
                  mat_A[24][27] * mat_B[27][6] +
                  mat_A[24][28] * mat_B[28][6] +
                  mat_A[24][29] * mat_B[29][6] +
                  mat_A[24][30] * mat_B[30][6] +
                  mat_A[24][31] * mat_B[31][6];
    mat_C[24][7] <= 
                  mat_A[24][0] * mat_B[0][7] +
                  mat_A[24][1] * mat_B[1][7] +
                  mat_A[24][2] * mat_B[2][7] +
                  mat_A[24][3] * mat_B[3][7] +
                  mat_A[24][4] * mat_B[4][7] +
                  mat_A[24][5] * mat_B[5][7] +
                  mat_A[24][6] * mat_B[6][7] +
                  mat_A[24][7] * mat_B[7][7] +
                  mat_A[24][8] * mat_B[8][7] +
                  mat_A[24][9] * mat_B[9][7] +
                  mat_A[24][10] * mat_B[10][7] +
                  mat_A[24][11] * mat_B[11][7] +
                  mat_A[24][12] * mat_B[12][7] +
                  mat_A[24][13] * mat_B[13][7] +
                  mat_A[24][14] * mat_B[14][7] +
                  mat_A[24][15] * mat_B[15][7] +
                  mat_A[24][16] * mat_B[16][7] +
                  mat_A[24][17] * mat_B[17][7] +
                  mat_A[24][18] * mat_B[18][7] +
                  mat_A[24][19] * mat_B[19][7] +
                  mat_A[24][20] * mat_B[20][7] +
                  mat_A[24][21] * mat_B[21][7] +
                  mat_A[24][22] * mat_B[22][7] +
                  mat_A[24][23] * mat_B[23][7] +
                  mat_A[24][24] * mat_B[24][7] +
                  mat_A[24][25] * mat_B[25][7] +
                  mat_A[24][26] * mat_B[26][7] +
                  mat_A[24][27] * mat_B[27][7] +
                  mat_A[24][28] * mat_B[28][7] +
                  mat_A[24][29] * mat_B[29][7] +
                  mat_A[24][30] * mat_B[30][7] +
                  mat_A[24][31] * mat_B[31][7];
    mat_C[24][8] <= 
                  mat_A[24][0] * mat_B[0][8] +
                  mat_A[24][1] * mat_B[1][8] +
                  mat_A[24][2] * mat_B[2][8] +
                  mat_A[24][3] * mat_B[3][8] +
                  mat_A[24][4] * mat_B[4][8] +
                  mat_A[24][5] * mat_B[5][8] +
                  mat_A[24][6] * mat_B[6][8] +
                  mat_A[24][7] * mat_B[7][8] +
                  mat_A[24][8] * mat_B[8][8] +
                  mat_A[24][9] * mat_B[9][8] +
                  mat_A[24][10] * mat_B[10][8] +
                  mat_A[24][11] * mat_B[11][8] +
                  mat_A[24][12] * mat_B[12][8] +
                  mat_A[24][13] * mat_B[13][8] +
                  mat_A[24][14] * mat_B[14][8] +
                  mat_A[24][15] * mat_B[15][8] +
                  mat_A[24][16] * mat_B[16][8] +
                  mat_A[24][17] * mat_B[17][8] +
                  mat_A[24][18] * mat_B[18][8] +
                  mat_A[24][19] * mat_B[19][8] +
                  mat_A[24][20] * mat_B[20][8] +
                  mat_A[24][21] * mat_B[21][8] +
                  mat_A[24][22] * mat_B[22][8] +
                  mat_A[24][23] * mat_B[23][8] +
                  mat_A[24][24] * mat_B[24][8] +
                  mat_A[24][25] * mat_B[25][8] +
                  mat_A[24][26] * mat_B[26][8] +
                  mat_A[24][27] * mat_B[27][8] +
                  mat_A[24][28] * mat_B[28][8] +
                  mat_A[24][29] * mat_B[29][8] +
                  mat_A[24][30] * mat_B[30][8] +
                  mat_A[24][31] * mat_B[31][8];
    mat_C[24][9] <= 
                  mat_A[24][0] * mat_B[0][9] +
                  mat_A[24][1] * mat_B[1][9] +
                  mat_A[24][2] * mat_B[2][9] +
                  mat_A[24][3] * mat_B[3][9] +
                  mat_A[24][4] * mat_B[4][9] +
                  mat_A[24][5] * mat_B[5][9] +
                  mat_A[24][6] * mat_B[6][9] +
                  mat_A[24][7] * mat_B[7][9] +
                  mat_A[24][8] * mat_B[8][9] +
                  mat_A[24][9] * mat_B[9][9] +
                  mat_A[24][10] * mat_B[10][9] +
                  mat_A[24][11] * mat_B[11][9] +
                  mat_A[24][12] * mat_B[12][9] +
                  mat_A[24][13] * mat_B[13][9] +
                  mat_A[24][14] * mat_B[14][9] +
                  mat_A[24][15] * mat_B[15][9] +
                  mat_A[24][16] * mat_B[16][9] +
                  mat_A[24][17] * mat_B[17][9] +
                  mat_A[24][18] * mat_B[18][9] +
                  mat_A[24][19] * mat_B[19][9] +
                  mat_A[24][20] * mat_B[20][9] +
                  mat_A[24][21] * mat_B[21][9] +
                  mat_A[24][22] * mat_B[22][9] +
                  mat_A[24][23] * mat_B[23][9] +
                  mat_A[24][24] * mat_B[24][9] +
                  mat_A[24][25] * mat_B[25][9] +
                  mat_A[24][26] * mat_B[26][9] +
                  mat_A[24][27] * mat_B[27][9] +
                  mat_A[24][28] * mat_B[28][9] +
                  mat_A[24][29] * mat_B[29][9] +
                  mat_A[24][30] * mat_B[30][9] +
                  mat_A[24][31] * mat_B[31][9];
    mat_C[24][10] <= 
                  mat_A[24][0] * mat_B[0][10] +
                  mat_A[24][1] * mat_B[1][10] +
                  mat_A[24][2] * mat_B[2][10] +
                  mat_A[24][3] * mat_B[3][10] +
                  mat_A[24][4] * mat_B[4][10] +
                  mat_A[24][5] * mat_B[5][10] +
                  mat_A[24][6] * mat_B[6][10] +
                  mat_A[24][7] * mat_B[7][10] +
                  mat_A[24][8] * mat_B[8][10] +
                  mat_A[24][9] * mat_B[9][10] +
                  mat_A[24][10] * mat_B[10][10] +
                  mat_A[24][11] * mat_B[11][10] +
                  mat_A[24][12] * mat_B[12][10] +
                  mat_A[24][13] * mat_B[13][10] +
                  mat_A[24][14] * mat_B[14][10] +
                  mat_A[24][15] * mat_B[15][10] +
                  mat_A[24][16] * mat_B[16][10] +
                  mat_A[24][17] * mat_B[17][10] +
                  mat_A[24][18] * mat_B[18][10] +
                  mat_A[24][19] * mat_B[19][10] +
                  mat_A[24][20] * mat_B[20][10] +
                  mat_A[24][21] * mat_B[21][10] +
                  mat_A[24][22] * mat_B[22][10] +
                  mat_A[24][23] * mat_B[23][10] +
                  mat_A[24][24] * mat_B[24][10] +
                  mat_A[24][25] * mat_B[25][10] +
                  mat_A[24][26] * mat_B[26][10] +
                  mat_A[24][27] * mat_B[27][10] +
                  mat_A[24][28] * mat_B[28][10] +
                  mat_A[24][29] * mat_B[29][10] +
                  mat_A[24][30] * mat_B[30][10] +
                  mat_A[24][31] * mat_B[31][10];
    mat_C[24][11] <= 
                  mat_A[24][0] * mat_B[0][11] +
                  mat_A[24][1] * mat_B[1][11] +
                  mat_A[24][2] * mat_B[2][11] +
                  mat_A[24][3] * mat_B[3][11] +
                  mat_A[24][4] * mat_B[4][11] +
                  mat_A[24][5] * mat_B[5][11] +
                  mat_A[24][6] * mat_B[6][11] +
                  mat_A[24][7] * mat_B[7][11] +
                  mat_A[24][8] * mat_B[8][11] +
                  mat_A[24][9] * mat_B[9][11] +
                  mat_A[24][10] * mat_B[10][11] +
                  mat_A[24][11] * mat_B[11][11] +
                  mat_A[24][12] * mat_B[12][11] +
                  mat_A[24][13] * mat_B[13][11] +
                  mat_A[24][14] * mat_B[14][11] +
                  mat_A[24][15] * mat_B[15][11] +
                  mat_A[24][16] * mat_B[16][11] +
                  mat_A[24][17] * mat_B[17][11] +
                  mat_A[24][18] * mat_B[18][11] +
                  mat_A[24][19] * mat_B[19][11] +
                  mat_A[24][20] * mat_B[20][11] +
                  mat_A[24][21] * mat_B[21][11] +
                  mat_A[24][22] * mat_B[22][11] +
                  mat_A[24][23] * mat_B[23][11] +
                  mat_A[24][24] * mat_B[24][11] +
                  mat_A[24][25] * mat_B[25][11] +
                  mat_A[24][26] * mat_B[26][11] +
                  mat_A[24][27] * mat_B[27][11] +
                  mat_A[24][28] * mat_B[28][11] +
                  mat_A[24][29] * mat_B[29][11] +
                  mat_A[24][30] * mat_B[30][11] +
                  mat_A[24][31] * mat_B[31][11];
    mat_C[24][12] <= 
                  mat_A[24][0] * mat_B[0][12] +
                  mat_A[24][1] * mat_B[1][12] +
                  mat_A[24][2] * mat_B[2][12] +
                  mat_A[24][3] * mat_B[3][12] +
                  mat_A[24][4] * mat_B[4][12] +
                  mat_A[24][5] * mat_B[5][12] +
                  mat_A[24][6] * mat_B[6][12] +
                  mat_A[24][7] * mat_B[7][12] +
                  mat_A[24][8] * mat_B[8][12] +
                  mat_A[24][9] * mat_B[9][12] +
                  mat_A[24][10] * mat_B[10][12] +
                  mat_A[24][11] * mat_B[11][12] +
                  mat_A[24][12] * mat_B[12][12] +
                  mat_A[24][13] * mat_B[13][12] +
                  mat_A[24][14] * mat_B[14][12] +
                  mat_A[24][15] * mat_B[15][12] +
                  mat_A[24][16] * mat_B[16][12] +
                  mat_A[24][17] * mat_B[17][12] +
                  mat_A[24][18] * mat_B[18][12] +
                  mat_A[24][19] * mat_B[19][12] +
                  mat_A[24][20] * mat_B[20][12] +
                  mat_A[24][21] * mat_B[21][12] +
                  mat_A[24][22] * mat_B[22][12] +
                  mat_A[24][23] * mat_B[23][12] +
                  mat_A[24][24] * mat_B[24][12] +
                  mat_A[24][25] * mat_B[25][12] +
                  mat_A[24][26] * mat_B[26][12] +
                  mat_A[24][27] * mat_B[27][12] +
                  mat_A[24][28] * mat_B[28][12] +
                  mat_A[24][29] * mat_B[29][12] +
                  mat_A[24][30] * mat_B[30][12] +
                  mat_A[24][31] * mat_B[31][12];
    mat_C[24][13] <= 
                  mat_A[24][0] * mat_B[0][13] +
                  mat_A[24][1] * mat_B[1][13] +
                  mat_A[24][2] * mat_B[2][13] +
                  mat_A[24][3] * mat_B[3][13] +
                  mat_A[24][4] * mat_B[4][13] +
                  mat_A[24][5] * mat_B[5][13] +
                  mat_A[24][6] * mat_B[6][13] +
                  mat_A[24][7] * mat_B[7][13] +
                  mat_A[24][8] * mat_B[8][13] +
                  mat_A[24][9] * mat_B[9][13] +
                  mat_A[24][10] * mat_B[10][13] +
                  mat_A[24][11] * mat_B[11][13] +
                  mat_A[24][12] * mat_B[12][13] +
                  mat_A[24][13] * mat_B[13][13] +
                  mat_A[24][14] * mat_B[14][13] +
                  mat_A[24][15] * mat_B[15][13] +
                  mat_A[24][16] * mat_B[16][13] +
                  mat_A[24][17] * mat_B[17][13] +
                  mat_A[24][18] * mat_B[18][13] +
                  mat_A[24][19] * mat_B[19][13] +
                  mat_A[24][20] * mat_B[20][13] +
                  mat_A[24][21] * mat_B[21][13] +
                  mat_A[24][22] * mat_B[22][13] +
                  mat_A[24][23] * mat_B[23][13] +
                  mat_A[24][24] * mat_B[24][13] +
                  mat_A[24][25] * mat_B[25][13] +
                  mat_A[24][26] * mat_B[26][13] +
                  mat_A[24][27] * mat_B[27][13] +
                  mat_A[24][28] * mat_B[28][13] +
                  mat_A[24][29] * mat_B[29][13] +
                  mat_A[24][30] * mat_B[30][13] +
                  mat_A[24][31] * mat_B[31][13];
    mat_C[24][14] <= 
                  mat_A[24][0] * mat_B[0][14] +
                  mat_A[24][1] * mat_B[1][14] +
                  mat_A[24][2] * mat_B[2][14] +
                  mat_A[24][3] * mat_B[3][14] +
                  mat_A[24][4] * mat_B[4][14] +
                  mat_A[24][5] * mat_B[5][14] +
                  mat_A[24][6] * mat_B[6][14] +
                  mat_A[24][7] * mat_B[7][14] +
                  mat_A[24][8] * mat_B[8][14] +
                  mat_A[24][9] * mat_B[9][14] +
                  mat_A[24][10] * mat_B[10][14] +
                  mat_A[24][11] * mat_B[11][14] +
                  mat_A[24][12] * mat_B[12][14] +
                  mat_A[24][13] * mat_B[13][14] +
                  mat_A[24][14] * mat_B[14][14] +
                  mat_A[24][15] * mat_B[15][14] +
                  mat_A[24][16] * mat_B[16][14] +
                  mat_A[24][17] * mat_B[17][14] +
                  mat_A[24][18] * mat_B[18][14] +
                  mat_A[24][19] * mat_B[19][14] +
                  mat_A[24][20] * mat_B[20][14] +
                  mat_A[24][21] * mat_B[21][14] +
                  mat_A[24][22] * mat_B[22][14] +
                  mat_A[24][23] * mat_B[23][14] +
                  mat_A[24][24] * mat_B[24][14] +
                  mat_A[24][25] * mat_B[25][14] +
                  mat_A[24][26] * mat_B[26][14] +
                  mat_A[24][27] * mat_B[27][14] +
                  mat_A[24][28] * mat_B[28][14] +
                  mat_A[24][29] * mat_B[29][14] +
                  mat_A[24][30] * mat_B[30][14] +
                  mat_A[24][31] * mat_B[31][14];
    mat_C[24][15] <= 
                  mat_A[24][0] * mat_B[0][15] +
                  mat_A[24][1] * mat_B[1][15] +
                  mat_A[24][2] * mat_B[2][15] +
                  mat_A[24][3] * mat_B[3][15] +
                  mat_A[24][4] * mat_B[4][15] +
                  mat_A[24][5] * mat_B[5][15] +
                  mat_A[24][6] * mat_B[6][15] +
                  mat_A[24][7] * mat_B[7][15] +
                  mat_A[24][8] * mat_B[8][15] +
                  mat_A[24][9] * mat_B[9][15] +
                  mat_A[24][10] * mat_B[10][15] +
                  mat_A[24][11] * mat_B[11][15] +
                  mat_A[24][12] * mat_B[12][15] +
                  mat_A[24][13] * mat_B[13][15] +
                  mat_A[24][14] * mat_B[14][15] +
                  mat_A[24][15] * mat_B[15][15] +
                  mat_A[24][16] * mat_B[16][15] +
                  mat_A[24][17] * mat_B[17][15] +
                  mat_A[24][18] * mat_B[18][15] +
                  mat_A[24][19] * mat_B[19][15] +
                  mat_A[24][20] * mat_B[20][15] +
                  mat_A[24][21] * mat_B[21][15] +
                  mat_A[24][22] * mat_B[22][15] +
                  mat_A[24][23] * mat_B[23][15] +
                  mat_A[24][24] * mat_B[24][15] +
                  mat_A[24][25] * mat_B[25][15] +
                  mat_A[24][26] * mat_B[26][15] +
                  mat_A[24][27] * mat_B[27][15] +
                  mat_A[24][28] * mat_B[28][15] +
                  mat_A[24][29] * mat_B[29][15] +
                  mat_A[24][30] * mat_B[30][15] +
                  mat_A[24][31] * mat_B[31][15];
    mat_C[24][16] <= 
                  mat_A[24][0] * mat_B[0][16] +
                  mat_A[24][1] * mat_B[1][16] +
                  mat_A[24][2] * mat_B[2][16] +
                  mat_A[24][3] * mat_B[3][16] +
                  mat_A[24][4] * mat_B[4][16] +
                  mat_A[24][5] * mat_B[5][16] +
                  mat_A[24][6] * mat_B[6][16] +
                  mat_A[24][7] * mat_B[7][16] +
                  mat_A[24][8] * mat_B[8][16] +
                  mat_A[24][9] * mat_B[9][16] +
                  mat_A[24][10] * mat_B[10][16] +
                  mat_A[24][11] * mat_B[11][16] +
                  mat_A[24][12] * mat_B[12][16] +
                  mat_A[24][13] * mat_B[13][16] +
                  mat_A[24][14] * mat_B[14][16] +
                  mat_A[24][15] * mat_B[15][16] +
                  mat_A[24][16] * mat_B[16][16] +
                  mat_A[24][17] * mat_B[17][16] +
                  mat_A[24][18] * mat_B[18][16] +
                  mat_A[24][19] * mat_B[19][16] +
                  mat_A[24][20] * mat_B[20][16] +
                  mat_A[24][21] * mat_B[21][16] +
                  mat_A[24][22] * mat_B[22][16] +
                  mat_A[24][23] * mat_B[23][16] +
                  mat_A[24][24] * mat_B[24][16] +
                  mat_A[24][25] * mat_B[25][16] +
                  mat_A[24][26] * mat_B[26][16] +
                  mat_A[24][27] * mat_B[27][16] +
                  mat_A[24][28] * mat_B[28][16] +
                  mat_A[24][29] * mat_B[29][16] +
                  mat_A[24][30] * mat_B[30][16] +
                  mat_A[24][31] * mat_B[31][16];
    mat_C[24][17] <= 
                  mat_A[24][0] * mat_B[0][17] +
                  mat_A[24][1] * mat_B[1][17] +
                  mat_A[24][2] * mat_B[2][17] +
                  mat_A[24][3] * mat_B[3][17] +
                  mat_A[24][4] * mat_B[4][17] +
                  mat_A[24][5] * mat_B[5][17] +
                  mat_A[24][6] * mat_B[6][17] +
                  mat_A[24][7] * mat_B[7][17] +
                  mat_A[24][8] * mat_B[8][17] +
                  mat_A[24][9] * mat_B[9][17] +
                  mat_A[24][10] * mat_B[10][17] +
                  mat_A[24][11] * mat_B[11][17] +
                  mat_A[24][12] * mat_B[12][17] +
                  mat_A[24][13] * mat_B[13][17] +
                  mat_A[24][14] * mat_B[14][17] +
                  mat_A[24][15] * mat_B[15][17] +
                  mat_A[24][16] * mat_B[16][17] +
                  mat_A[24][17] * mat_B[17][17] +
                  mat_A[24][18] * mat_B[18][17] +
                  mat_A[24][19] * mat_B[19][17] +
                  mat_A[24][20] * mat_B[20][17] +
                  mat_A[24][21] * mat_B[21][17] +
                  mat_A[24][22] * mat_B[22][17] +
                  mat_A[24][23] * mat_B[23][17] +
                  mat_A[24][24] * mat_B[24][17] +
                  mat_A[24][25] * mat_B[25][17] +
                  mat_A[24][26] * mat_B[26][17] +
                  mat_A[24][27] * mat_B[27][17] +
                  mat_A[24][28] * mat_B[28][17] +
                  mat_A[24][29] * mat_B[29][17] +
                  mat_A[24][30] * mat_B[30][17] +
                  mat_A[24][31] * mat_B[31][17];
    mat_C[24][18] <= 
                  mat_A[24][0] * mat_B[0][18] +
                  mat_A[24][1] * mat_B[1][18] +
                  mat_A[24][2] * mat_B[2][18] +
                  mat_A[24][3] * mat_B[3][18] +
                  mat_A[24][4] * mat_B[4][18] +
                  mat_A[24][5] * mat_B[5][18] +
                  mat_A[24][6] * mat_B[6][18] +
                  mat_A[24][7] * mat_B[7][18] +
                  mat_A[24][8] * mat_B[8][18] +
                  mat_A[24][9] * mat_B[9][18] +
                  mat_A[24][10] * mat_B[10][18] +
                  mat_A[24][11] * mat_B[11][18] +
                  mat_A[24][12] * mat_B[12][18] +
                  mat_A[24][13] * mat_B[13][18] +
                  mat_A[24][14] * mat_B[14][18] +
                  mat_A[24][15] * mat_B[15][18] +
                  mat_A[24][16] * mat_B[16][18] +
                  mat_A[24][17] * mat_B[17][18] +
                  mat_A[24][18] * mat_B[18][18] +
                  mat_A[24][19] * mat_B[19][18] +
                  mat_A[24][20] * mat_B[20][18] +
                  mat_A[24][21] * mat_B[21][18] +
                  mat_A[24][22] * mat_B[22][18] +
                  mat_A[24][23] * mat_B[23][18] +
                  mat_A[24][24] * mat_B[24][18] +
                  mat_A[24][25] * mat_B[25][18] +
                  mat_A[24][26] * mat_B[26][18] +
                  mat_A[24][27] * mat_B[27][18] +
                  mat_A[24][28] * mat_B[28][18] +
                  mat_A[24][29] * mat_B[29][18] +
                  mat_A[24][30] * mat_B[30][18] +
                  mat_A[24][31] * mat_B[31][18];
    mat_C[24][19] <= 
                  mat_A[24][0] * mat_B[0][19] +
                  mat_A[24][1] * mat_B[1][19] +
                  mat_A[24][2] * mat_B[2][19] +
                  mat_A[24][3] * mat_B[3][19] +
                  mat_A[24][4] * mat_B[4][19] +
                  mat_A[24][5] * mat_B[5][19] +
                  mat_A[24][6] * mat_B[6][19] +
                  mat_A[24][7] * mat_B[7][19] +
                  mat_A[24][8] * mat_B[8][19] +
                  mat_A[24][9] * mat_B[9][19] +
                  mat_A[24][10] * mat_B[10][19] +
                  mat_A[24][11] * mat_B[11][19] +
                  mat_A[24][12] * mat_B[12][19] +
                  mat_A[24][13] * mat_B[13][19] +
                  mat_A[24][14] * mat_B[14][19] +
                  mat_A[24][15] * mat_B[15][19] +
                  mat_A[24][16] * mat_B[16][19] +
                  mat_A[24][17] * mat_B[17][19] +
                  mat_A[24][18] * mat_B[18][19] +
                  mat_A[24][19] * mat_B[19][19] +
                  mat_A[24][20] * mat_B[20][19] +
                  mat_A[24][21] * mat_B[21][19] +
                  mat_A[24][22] * mat_B[22][19] +
                  mat_A[24][23] * mat_B[23][19] +
                  mat_A[24][24] * mat_B[24][19] +
                  mat_A[24][25] * mat_B[25][19] +
                  mat_A[24][26] * mat_B[26][19] +
                  mat_A[24][27] * mat_B[27][19] +
                  mat_A[24][28] * mat_B[28][19] +
                  mat_A[24][29] * mat_B[29][19] +
                  mat_A[24][30] * mat_B[30][19] +
                  mat_A[24][31] * mat_B[31][19];
    mat_C[24][20] <= 
                  mat_A[24][0] * mat_B[0][20] +
                  mat_A[24][1] * mat_B[1][20] +
                  mat_A[24][2] * mat_B[2][20] +
                  mat_A[24][3] * mat_B[3][20] +
                  mat_A[24][4] * mat_B[4][20] +
                  mat_A[24][5] * mat_B[5][20] +
                  mat_A[24][6] * mat_B[6][20] +
                  mat_A[24][7] * mat_B[7][20] +
                  mat_A[24][8] * mat_B[8][20] +
                  mat_A[24][9] * mat_B[9][20] +
                  mat_A[24][10] * mat_B[10][20] +
                  mat_A[24][11] * mat_B[11][20] +
                  mat_A[24][12] * mat_B[12][20] +
                  mat_A[24][13] * mat_B[13][20] +
                  mat_A[24][14] * mat_B[14][20] +
                  mat_A[24][15] * mat_B[15][20] +
                  mat_A[24][16] * mat_B[16][20] +
                  mat_A[24][17] * mat_B[17][20] +
                  mat_A[24][18] * mat_B[18][20] +
                  mat_A[24][19] * mat_B[19][20] +
                  mat_A[24][20] * mat_B[20][20] +
                  mat_A[24][21] * mat_B[21][20] +
                  mat_A[24][22] * mat_B[22][20] +
                  mat_A[24][23] * mat_B[23][20] +
                  mat_A[24][24] * mat_B[24][20] +
                  mat_A[24][25] * mat_B[25][20] +
                  mat_A[24][26] * mat_B[26][20] +
                  mat_A[24][27] * mat_B[27][20] +
                  mat_A[24][28] * mat_B[28][20] +
                  mat_A[24][29] * mat_B[29][20] +
                  mat_A[24][30] * mat_B[30][20] +
                  mat_A[24][31] * mat_B[31][20];
    mat_C[24][21] <= 
                  mat_A[24][0] * mat_B[0][21] +
                  mat_A[24][1] * mat_B[1][21] +
                  mat_A[24][2] * mat_B[2][21] +
                  mat_A[24][3] * mat_B[3][21] +
                  mat_A[24][4] * mat_B[4][21] +
                  mat_A[24][5] * mat_B[5][21] +
                  mat_A[24][6] * mat_B[6][21] +
                  mat_A[24][7] * mat_B[7][21] +
                  mat_A[24][8] * mat_B[8][21] +
                  mat_A[24][9] * mat_B[9][21] +
                  mat_A[24][10] * mat_B[10][21] +
                  mat_A[24][11] * mat_B[11][21] +
                  mat_A[24][12] * mat_B[12][21] +
                  mat_A[24][13] * mat_B[13][21] +
                  mat_A[24][14] * mat_B[14][21] +
                  mat_A[24][15] * mat_B[15][21] +
                  mat_A[24][16] * mat_B[16][21] +
                  mat_A[24][17] * mat_B[17][21] +
                  mat_A[24][18] * mat_B[18][21] +
                  mat_A[24][19] * mat_B[19][21] +
                  mat_A[24][20] * mat_B[20][21] +
                  mat_A[24][21] * mat_B[21][21] +
                  mat_A[24][22] * mat_B[22][21] +
                  mat_A[24][23] * mat_B[23][21] +
                  mat_A[24][24] * mat_B[24][21] +
                  mat_A[24][25] * mat_B[25][21] +
                  mat_A[24][26] * mat_B[26][21] +
                  mat_A[24][27] * mat_B[27][21] +
                  mat_A[24][28] * mat_B[28][21] +
                  mat_A[24][29] * mat_B[29][21] +
                  mat_A[24][30] * mat_B[30][21] +
                  mat_A[24][31] * mat_B[31][21];
    mat_C[24][22] <= 
                  mat_A[24][0] * mat_B[0][22] +
                  mat_A[24][1] * mat_B[1][22] +
                  mat_A[24][2] * mat_B[2][22] +
                  mat_A[24][3] * mat_B[3][22] +
                  mat_A[24][4] * mat_B[4][22] +
                  mat_A[24][5] * mat_B[5][22] +
                  mat_A[24][6] * mat_B[6][22] +
                  mat_A[24][7] * mat_B[7][22] +
                  mat_A[24][8] * mat_B[8][22] +
                  mat_A[24][9] * mat_B[9][22] +
                  mat_A[24][10] * mat_B[10][22] +
                  mat_A[24][11] * mat_B[11][22] +
                  mat_A[24][12] * mat_B[12][22] +
                  mat_A[24][13] * mat_B[13][22] +
                  mat_A[24][14] * mat_B[14][22] +
                  mat_A[24][15] * mat_B[15][22] +
                  mat_A[24][16] * mat_B[16][22] +
                  mat_A[24][17] * mat_B[17][22] +
                  mat_A[24][18] * mat_B[18][22] +
                  mat_A[24][19] * mat_B[19][22] +
                  mat_A[24][20] * mat_B[20][22] +
                  mat_A[24][21] * mat_B[21][22] +
                  mat_A[24][22] * mat_B[22][22] +
                  mat_A[24][23] * mat_B[23][22] +
                  mat_A[24][24] * mat_B[24][22] +
                  mat_A[24][25] * mat_B[25][22] +
                  mat_A[24][26] * mat_B[26][22] +
                  mat_A[24][27] * mat_B[27][22] +
                  mat_A[24][28] * mat_B[28][22] +
                  mat_A[24][29] * mat_B[29][22] +
                  mat_A[24][30] * mat_B[30][22] +
                  mat_A[24][31] * mat_B[31][22];
    mat_C[24][23] <= 
                  mat_A[24][0] * mat_B[0][23] +
                  mat_A[24][1] * mat_B[1][23] +
                  mat_A[24][2] * mat_B[2][23] +
                  mat_A[24][3] * mat_B[3][23] +
                  mat_A[24][4] * mat_B[4][23] +
                  mat_A[24][5] * mat_B[5][23] +
                  mat_A[24][6] * mat_B[6][23] +
                  mat_A[24][7] * mat_B[7][23] +
                  mat_A[24][8] * mat_B[8][23] +
                  mat_A[24][9] * mat_B[9][23] +
                  mat_A[24][10] * mat_B[10][23] +
                  mat_A[24][11] * mat_B[11][23] +
                  mat_A[24][12] * mat_B[12][23] +
                  mat_A[24][13] * mat_B[13][23] +
                  mat_A[24][14] * mat_B[14][23] +
                  mat_A[24][15] * mat_B[15][23] +
                  mat_A[24][16] * mat_B[16][23] +
                  mat_A[24][17] * mat_B[17][23] +
                  mat_A[24][18] * mat_B[18][23] +
                  mat_A[24][19] * mat_B[19][23] +
                  mat_A[24][20] * mat_B[20][23] +
                  mat_A[24][21] * mat_B[21][23] +
                  mat_A[24][22] * mat_B[22][23] +
                  mat_A[24][23] * mat_B[23][23] +
                  mat_A[24][24] * mat_B[24][23] +
                  mat_A[24][25] * mat_B[25][23] +
                  mat_A[24][26] * mat_B[26][23] +
                  mat_A[24][27] * mat_B[27][23] +
                  mat_A[24][28] * mat_B[28][23] +
                  mat_A[24][29] * mat_B[29][23] +
                  mat_A[24][30] * mat_B[30][23] +
                  mat_A[24][31] * mat_B[31][23];
    mat_C[24][24] <= 
                  mat_A[24][0] * mat_B[0][24] +
                  mat_A[24][1] * mat_B[1][24] +
                  mat_A[24][2] * mat_B[2][24] +
                  mat_A[24][3] * mat_B[3][24] +
                  mat_A[24][4] * mat_B[4][24] +
                  mat_A[24][5] * mat_B[5][24] +
                  mat_A[24][6] * mat_B[6][24] +
                  mat_A[24][7] * mat_B[7][24] +
                  mat_A[24][8] * mat_B[8][24] +
                  mat_A[24][9] * mat_B[9][24] +
                  mat_A[24][10] * mat_B[10][24] +
                  mat_A[24][11] * mat_B[11][24] +
                  mat_A[24][12] * mat_B[12][24] +
                  mat_A[24][13] * mat_B[13][24] +
                  mat_A[24][14] * mat_B[14][24] +
                  mat_A[24][15] * mat_B[15][24] +
                  mat_A[24][16] * mat_B[16][24] +
                  mat_A[24][17] * mat_B[17][24] +
                  mat_A[24][18] * mat_B[18][24] +
                  mat_A[24][19] * mat_B[19][24] +
                  mat_A[24][20] * mat_B[20][24] +
                  mat_A[24][21] * mat_B[21][24] +
                  mat_A[24][22] * mat_B[22][24] +
                  mat_A[24][23] * mat_B[23][24] +
                  mat_A[24][24] * mat_B[24][24] +
                  mat_A[24][25] * mat_B[25][24] +
                  mat_A[24][26] * mat_B[26][24] +
                  mat_A[24][27] * mat_B[27][24] +
                  mat_A[24][28] * mat_B[28][24] +
                  mat_A[24][29] * mat_B[29][24] +
                  mat_A[24][30] * mat_B[30][24] +
                  mat_A[24][31] * mat_B[31][24];
    mat_C[24][25] <= 
                  mat_A[24][0] * mat_B[0][25] +
                  mat_A[24][1] * mat_B[1][25] +
                  mat_A[24][2] * mat_B[2][25] +
                  mat_A[24][3] * mat_B[3][25] +
                  mat_A[24][4] * mat_B[4][25] +
                  mat_A[24][5] * mat_B[5][25] +
                  mat_A[24][6] * mat_B[6][25] +
                  mat_A[24][7] * mat_B[7][25] +
                  mat_A[24][8] * mat_B[8][25] +
                  mat_A[24][9] * mat_B[9][25] +
                  mat_A[24][10] * mat_B[10][25] +
                  mat_A[24][11] * mat_B[11][25] +
                  mat_A[24][12] * mat_B[12][25] +
                  mat_A[24][13] * mat_B[13][25] +
                  mat_A[24][14] * mat_B[14][25] +
                  mat_A[24][15] * mat_B[15][25] +
                  mat_A[24][16] * mat_B[16][25] +
                  mat_A[24][17] * mat_B[17][25] +
                  mat_A[24][18] * mat_B[18][25] +
                  mat_A[24][19] * mat_B[19][25] +
                  mat_A[24][20] * mat_B[20][25] +
                  mat_A[24][21] * mat_B[21][25] +
                  mat_A[24][22] * mat_B[22][25] +
                  mat_A[24][23] * mat_B[23][25] +
                  mat_A[24][24] * mat_B[24][25] +
                  mat_A[24][25] * mat_B[25][25] +
                  mat_A[24][26] * mat_B[26][25] +
                  mat_A[24][27] * mat_B[27][25] +
                  mat_A[24][28] * mat_B[28][25] +
                  mat_A[24][29] * mat_B[29][25] +
                  mat_A[24][30] * mat_B[30][25] +
                  mat_A[24][31] * mat_B[31][25];
    mat_C[24][26] <= 
                  mat_A[24][0] * mat_B[0][26] +
                  mat_A[24][1] * mat_B[1][26] +
                  mat_A[24][2] * mat_B[2][26] +
                  mat_A[24][3] * mat_B[3][26] +
                  mat_A[24][4] * mat_B[4][26] +
                  mat_A[24][5] * mat_B[5][26] +
                  mat_A[24][6] * mat_B[6][26] +
                  mat_A[24][7] * mat_B[7][26] +
                  mat_A[24][8] * mat_B[8][26] +
                  mat_A[24][9] * mat_B[9][26] +
                  mat_A[24][10] * mat_B[10][26] +
                  mat_A[24][11] * mat_B[11][26] +
                  mat_A[24][12] * mat_B[12][26] +
                  mat_A[24][13] * mat_B[13][26] +
                  mat_A[24][14] * mat_B[14][26] +
                  mat_A[24][15] * mat_B[15][26] +
                  mat_A[24][16] * mat_B[16][26] +
                  mat_A[24][17] * mat_B[17][26] +
                  mat_A[24][18] * mat_B[18][26] +
                  mat_A[24][19] * mat_B[19][26] +
                  mat_A[24][20] * mat_B[20][26] +
                  mat_A[24][21] * mat_B[21][26] +
                  mat_A[24][22] * mat_B[22][26] +
                  mat_A[24][23] * mat_B[23][26] +
                  mat_A[24][24] * mat_B[24][26] +
                  mat_A[24][25] * mat_B[25][26] +
                  mat_A[24][26] * mat_B[26][26] +
                  mat_A[24][27] * mat_B[27][26] +
                  mat_A[24][28] * mat_B[28][26] +
                  mat_A[24][29] * mat_B[29][26] +
                  mat_A[24][30] * mat_B[30][26] +
                  mat_A[24][31] * mat_B[31][26];
    mat_C[24][27] <= 
                  mat_A[24][0] * mat_B[0][27] +
                  mat_A[24][1] * mat_B[1][27] +
                  mat_A[24][2] * mat_B[2][27] +
                  mat_A[24][3] * mat_B[3][27] +
                  mat_A[24][4] * mat_B[4][27] +
                  mat_A[24][5] * mat_B[5][27] +
                  mat_A[24][6] * mat_B[6][27] +
                  mat_A[24][7] * mat_B[7][27] +
                  mat_A[24][8] * mat_B[8][27] +
                  mat_A[24][9] * mat_B[9][27] +
                  mat_A[24][10] * mat_B[10][27] +
                  mat_A[24][11] * mat_B[11][27] +
                  mat_A[24][12] * mat_B[12][27] +
                  mat_A[24][13] * mat_B[13][27] +
                  mat_A[24][14] * mat_B[14][27] +
                  mat_A[24][15] * mat_B[15][27] +
                  mat_A[24][16] * mat_B[16][27] +
                  mat_A[24][17] * mat_B[17][27] +
                  mat_A[24][18] * mat_B[18][27] +
                  mat_A[24][19] * mat_B[19][27] +
                  mat_A[24][20] * mat_B[20][27] +
                  mat_A[24][21] * mat_B[21][27] +
                  mat_A[24][22] * mat_B[22][27] +
                  mat_A[24][23] * mat_B[23][27] +
                  mat_A[24][24] * mat_B[24][27] +
                  mat_A[24][25] * mat_B[25][27] +
                  mat_A[24][26] * mat_B[26][27] +
                  mat_A[24][27] * mat_B[27][27] +
                  mat_A[24][28] * mat_B[28][27] +
                  mat_A[24][29] * mat_B[29][27] +
                  mat_A[24][30] * mat_B[30][27] +
                  mat_A[24][31] * mat_B[31][27];
    mat_C[24][28] <= 
                  mat_A[24][0] * mat_B[0][28] +
                  mat_A[24][1] * mat_B[1][28] +
                  mat_A[24][2] * mat_B[2][28] +
                  mat_A[24][3] * mat_B[3][28] +
                  mat_A[24][4] * mat_B[4][28] +
                  mat_A[24][5] * mat_B[5][28] +
                  mat_A[24][6] * mat_B[6][28] +
                  mat_A[24][7] * mat_B[7][28] +
                  mat_A[24][8] * mat_B[8][28] +
                  mat_A[24][9] * mat_B[9][28] +
                  mat_A[24][10] * mat_B[10][28] +
                  mat_A[24][11] * mat_B[11][28] +
                  mat_A[24][12] * mat_B[12][28] +
                  mat_A[24][13] * mat_B[13][28] +
                  mat_A[24][14] * mat_B[14][28] +
                  mat_A[24][15] * mat_B[15][28] +
                  mat_A[24][16] * mat_B[16][28] +
                  mat_A[24][17] * mat_B[17][28] +
                  mat_A[24][18] * mat_B[18][28] +
                  mat_A[24][19] * mat_B[19][28] +
                  mat_A[24][20] * mat_B[20][28] +
                  mat_A[24][21] * mat_B[21][28] +
                  mat_A[24][22] * mat_B[22][28] +
                  mat_A[24][23] * mat_B[23][28] +
                  mat_A[24][24] * mat_B[24][28] +
                  mat_A[24][25] * mat_B[25][28] +
                  mat_A[24][26] * mat_B[26][28] +
                  mat_A[24][27] * mat_B[27][28] +
                  mat_A[24][28] * mat_B[28][28] +
                  mat_A[24][29] * mat_B[29][28] +
                  mat_A[24][30] * mat_B[30][28] +
                  mat_A[24][31] * mat_B[31][28];
    mat_C[24][29] <= 
                  mat_A[24][0] * mat_B[0][29] +
                  mat_A[24][1] * mat_B[1][29] +
                  mat_A[24][2] * mat_B[2][29] +
                  mat_A[24][3] * mat_B[3][29] +
                  mat_A[24][4] * mat_B[4][29] +
                  mat_A[24][5] * mat_B[5][29] +
                  mat_A[24][6] * mat_B[6][29] +
                  mat_A[24][7] * mat_B[7][29] +
                  mat_A[24][8] * mat_B[8][29] +
                  mat_A[24][9] * mat_B[9][29] +
                  mat_A[24][10] * mat_B[10][29] +
                  mat_A[24][11] * mat_B[11][29] +
                  mat_A[24][12] * mat_B[12][29] +
                  mat_A[24][13] * mat_B[13][29] +
                  mat_A[24][14] * mat_B[14][29] +
                  mat_A[24][15] * mat_B[15][29] +
                  mat_A[24][16] * mat_B[16][29] +
                  mat_A[24][17] * mat_B[17][29] +
                  mat_A[24][18] * mat_B[18][29] +
                  mat_A[24][19] * mat_B[19][29] +
                  mat_A[24][20] * mat_B[20][29] +
                  mat_A[24][21] * mat_B[21][29] +
                  mat_A[24][22] * mat_B[22][29] +
                  mat_A[24][23] * mat_B[23][29] +
                  mat_A[24][24] * mat_B[24][29] +
                  mat_A[24][25] * mat_B[25][29] +
                  mat_A[24][26] * mat_B[26][29] +
                  mat_A[24][27] * mat_B[27][29] +
                  mat_A[24][28] * mat_B[28][29] +
                  mat_A[24][29] * mat_B[29][29] +
                  mat_A[24][30] * mat_B[30][29] +
                  mat_A[24][31] * mat_B[31][29];
    mat_C[24][30] <= 
                  mat_A[24][0] * mat_B[0][30] +
                  mat_A[24][1] * mat_B[1][30] +
                  mat_A[24][2] * mat_B[2][30] +
                  mat_A[24][3] * mat_B[3][30] +
                  mat_A[24][4] * mat_B[4][30] +
                  mat_A[24][5] * mat_B[5][30] +
                  mat_A[24][6] * mat_B[6][30] +
                  mat_A[24][7] * mat_B[7][30] +
                  mat_A[24][8] * mat_B[8][30] +
                  mat_A[24][9] * mat_B[9][30] +
                  mat_A[24][10] * mat_B[10][30] +
                  mat_A[24][11] * mat_B[11][30] +
                  mat_A[24][12] * mat_B[12][30] +
                  mat_A[24][13] * mat_B[13][30] +
                  mat_A[24][14] * mat_B[14][30] +
                  mat_A[24][15] * mat_B[15][30] +
                  mat_A[24][16] * mat_B[16][30] +
                  mat_A[24][17] * mat_B[17][30] +
                  mat_A[24][18] * mat_B[18][30] +
                  mat_A[24][19] * mat_B[19][30] +
                  mat_A[24][20] * mat_B[20][30] +
                  mat_A[24][21] * mat_B[21][30] +
                  mat_A[24][22] * mat_B[22][30] +
                  mat_A[24][23] * mat_B[23][30] +
                  mat_A[24][24] * mat_B[24][30] +
                  mat_A[24][25] * mat_B[25][30] +
                  mat_A[24][26] * mat_B[26][30] +
                  mat_A[24][27] * mat_B[27][30] +
                  mat_A[24][28] * mat_B[28][30] +
                  mat_A[24][29] * mat_B[29][30] +
                  mat_A[24][30] * mat_B[30][30] +
                  mat_A[24][31] * mat_B[31][30];
    mat_C[24][31] <= 
                  mat_A[24][0] * mat_B[0][31] +
                  mat_A[24][1] * mat_B[1][31] +
                  mat_A[24][2] * mat_B[2][31] +
                  mat_A[24][3] * mat_B[3][31] +
                  mat_A[24][4] * mat_B[4][31] +
                  mat_A[24][5] * mat_B[5][31] +
                  mat_A[24][6] * mat_B[6][31] +
                  mat_A[24][7] * mat_B[7][31] +
                  mat_A[24][8] * mat_B[8][31] +
                  mat_A[24][9] * mat_B[9][31] +
                  mat_A[24][10] * mat_B[10][31] +
                  mat_A[24][11] * mat_B[11][31] +
                  mat_A[24][12] * mat_B[12][31] +
                  mat_A[24][13] * mat_B[13][31] +
                  mat_A[24][14] * mat_B[14][31] +
                  mat_A[24][15] * mat_B[15][31] +
                  mat_A[24][16] * mat_B[16][31] +
                  mat_A[24][17] * mat_B[17][31] +
                  mat_A[24][18] * mat_B[18][31] +
                  mat_A[24][19] * mat_B[19][31] +
                  mat_A[24][20] * mat_B[20][31] +
                  mat_A[24][21] * mat_B[21][31] +
                  mat_A[24][22] * mat_B[22][31] +
                  mat_A[24][23] * mat_B[23][31] +
                  mat_A[24][24] * mat_B[24][31] +
                  mat_A[24][25] * mat_B[25][31] +
                  mat_A[24][26] * mat_B[26][31] +
                  mat_A[24][27] * mat_B[27][31] +
                  mat_A[24][28] * mat_B[28][31] +
                  mat_A[24][29] * mat_B[29][31] +
                  mat_A[24][30] * mat_B[30][31] +
                  mat_A[24][31] * mat_B[31][31];
    mat_C[25][0] <= 
                  mat_A[25][0] * mat_B[0][0] +
                  mat_A[25][1] * mat_B[1][0] +
                  mat_A[25][2] * mat_B[2][0] +
                  mat_A[25][3] * mat_B[3][0] +
                  mat_A[25][4] * mat_B[4][0] +
                  mat_A[25][5] * mat_B[5][0] +
                  mat_A[25][6] * mat_B[6][0] +
                  mat_A[25][7] * mat_B[7][0] +
                  mat_A[25][8] * mat_B[8][0] +
                  mat_A[25][9] * mat_B[9][0] +
                  mat_A[25][10] * mat_B[10][0] +
                  mat_A[25][11] * mat_B[11][0] +
                  mat_A[25][12] * mat_B[12][0] +
                  mat_A[25][13] * mat_B[13][0] +
                  mat_A[25][14] * mat_B[14][0] +
                  mat_A[25][15] * mat_B[15][0] +
                  mat_A[25][16] * mat_B[16][0] +
                  mat_A[25][17] * mat_B[17][0] +
                  mat_A[25][18] * mat_B[18][0] +
                  mat_A[25][19] * mat_B[19][0] +
                  mat_A[25][20] * mat_B[20][0] +
                  mat_A[25][21] * mat_B[21][0] +
                  mat_A[25][22] * mat_B[22][0] +
                  mat_A[25][23] * mat_B[23][0] +
                  mat_A[25][24] * mat_B[24][0] +
                  mat_A[25][25] * mat_B[25][0] +
                  mat_A[25][26] * mat_B[26][0] +
                  mat_A[25][27] * mat_B[27][0] +
                  mat_A[25][28] * mat_B[28][0] +
                  mat_A[25][29] * mat_B[29][0] +
                  mat_A[25][30] * mat_B[30][0] +
                  mat_A[25][31] * mat_B[31][0];
    mat_C[25][1] <= 
                  mat_A[25][0] * mat_B[0][1] +
                  mat_A[25][1] * mat_B[1][1] +
                  mat_A[25][2] * mat_B[2][1] +
                  mat_A[25][3] * mat_B[3][1] +
                  mat_A[25][4] * mat_B[4][1] +
                  mat_A[25][5] * mat_B[5][1] +
                  mat_A[25][6] * mat_B[6][1] +
                  mat_A[25][7] * mat_B[7][1] +
                  mat_A[25][8] * mat_B[8][1] +
                  mat_A[25][9] * mat_B[9][1] +
                  mat_A[25][10] * mat_B[10][1] +
                  mat_A[25][11] * mat_B[11][1] +
                  mat_A[25][12] * mat_B[12][1] +
                  mat_A[25][13] * mat_B[13][1] +
                  mat_A[25][14] * mat_B[14][1] +
                  mat_A[25][15] * mat_B[15][1] +
                  mat_A[25][16] * mat_B[16][1] +
                  mat_A[25][17] * mat_B[17][1] +
                  mat_A[25][18] * mat_B[18][1] +
                  mat_A[25][19] * mat_B[19][1] +
                  mat_A[25][20] * mat_B[20][1] +
                  mat_A[25][21] * mat_B[21][1] +
                  mat_A[25][22] * mat_B[22][1] +
                  mat_A[25][23] * mat_B[23][1] +
                  mat_A[25][24] * mat_B[24][1] +
                  mat_A[25][25] * mat_B[25][1] +
                  mat_A[25][26] * mat_B[26][1] +
                  mat_A[25][27] * mat_B[27][1] +
                  mat_A[25][28] * mat_B[28][1] +
                  mat_A[25][29] * mat_B[29][1] +
                  mat_A[25][30] * mat_B[30][1] +
                  mat_A[25][31] * mat_B[31][1];
    mat_C[25][2] <= 
                  mat_A[25][0] * mat_B[0][2] +
                  mat_A[25][1] * mat_B[1][2] +
                  mat_A[25][2] * mat_B[2][2] +
                  mat_A[25][3] * mat_B[3][2] +
                  mat_A[25][4] * mat_B[4][2] +
                  mat_A[25][5] * mat_B[5][2] +
                  mat_A[25][6] * mat_B[6][2] +
                  mat_A[25][7] * mat_B[7][2] +
                  mat_A[25][8] * mat_B[8][2] +
                  mat_A[25][9] * mat_B[9][2] +
                  mat_A[25][10] * mat_B[10][2] +
                  mat_A[25][11] * mat_B[11][2] +
                  mat_A[25][12] * mat_B[12][2] +
                  mat_A[25][13] * mat_B[13][2] +
                  mat_A[25][14] * mat_B[14][2] +
                  mat_A[25][15] * mat_B[15][2] +
                  mat_A[25][16] * mat_B[16][2] +
                  mat_A[25][17] * mat_B[17][2] +
                  mat_A[25][18] * mat_B[18][2] +
                  mat_A[25][19] * mat_B[19][2] +
                  mat_A[25][20] * mat_B[20][2] +
                  mat_A[25][21] * mat_B[21][2] +
                  mat_A[25][22] * mat_B[22][2] +
                  mat_A[25][23] * mat_B[23][2] +
                  mat_A[25][24] * mat_B[24][2] +
                  mat_A[25][25] * mat_B[25][2] +
                  mat_A[25][26] * mat_B[26][2] +
                  mat_A[25][27] * mat_B[27][2] +
                  mat_A[25][28] * mat_B[28][2] +
                  mat_A[25][29] * mat_B[29][2] +
                  mat_A[25][30] * mat_B[30][2] +
                  mat_A[25][31] * mat_B[31][2];
    mat_C[25][3] <= 
                  mat_A[25][0] * mat_B[0][3] +
                  mat_A[25][1] * mat_B[1][3] +
                  mat_A[25][2] * mat_B[2][3] +
                  mat_A[25][3] * mat_B[3][3] +
                  mat_A[25][4] * mat_B[4][3] +
                  mat_A[25][5] * mat_B[5][3] +
                  mat_A[25][6] * mat_B[6][3] +
                  mat_A[25][7] * mat_B[7][3] +
                  mat_A[25][8] * mat_B[8][3] +
                  mat_A[25][9] * mat_B[9][3] +
                  mat_A[25][10] * mat_B[10][3] +
                  mat_A[25][11] * mat_B[11][3] +
                  mat_A[25][12] * mat_B[12][3] +
                  mat_A[25][13] * mat_B[13][3] +
                  mat_A[25][14] * mat_B[14][3] +
                  mat_A[25][15] * mat_B[15][3] +
                  mat_A[25][16] * mat_B[16][3] +
                  mat_A[25][17] * mat_B[17][3] +
                  mat_A[25][18] * mat_B[18][3] +
                  mat_A[25][19] * mat_B[19][3] +
                  mat_A[25][20] * mat_B[20][3] +
                  mat_A[25][21] * mat_B[21][3] +
                  mat_A[25][22] * mat_B[22][3] +
                  mat_A[25][23] * mat_B[23][3] +
                  mat_A[25][24] * mat_B[24][3] +
                  mat_A[25][25] * mat_B[25][3] +
                  mat_A[25][26] * mat_B[26][3] +
                  mat_A[25][27] * mat_B[27][3] +
                  mat_A[25][28] * mat_B[28][3] +
                  mat_A[25][29] * mat_B[29][3] +
                  mat_A[25][30] * mat_B[30][3] +
                  mat_A[25][31] * mat_B[31][3];
    mat_C[25][4] <= 
                  mat_A[25][0] * mat_B[0][4] +
                  mat_A[25][1] * mat_B[1][4] +
                  mat_A[25][2] * mat_B[2][4] +
                  mat_A[25][3] * mat_B[3][4] +
                  mat_A[25][4] * mat_B[4][4] +
                  mat_A[25][5] * mat_B[5][4] +
                  mat_A[25][6] * mat_B[6][4] +
                  mat_A[25][7] * mat_B[7][4] +
                  mat_A[25][8] * mat_B[8][4] +
                  mat_A[25][9] * mat_B[9][4] +
                  mat_A[25][10] * mat_B[10][4] +
                  mat_A[25][11] * mat_B[11][4] +
                  mat_A[25][12] * mat_B[12][4] +
                  mat_A[25][13] * mat_B[13][4] +
                  mat_A[25][14] * mat_B[14][4] +
                  mat_A[25][15] * mat_B[15][4] +
                  mat_A[25][16] * mat_B[16][4] +
                  mat_A[25][17] * mat_B[17][4] +
                  mat_A[25][18] * mat_B[18][4] +
                  mat_A[25][19] * mat_B[19][4] +
                  mat_A[25][20] * mat_B[20][4] +
                  mat_A[25][21] * mat_B[21][4] +
                  mat_A[25][22] * mat_B[22][4] +
                  mat_A[25][23] * mat_B[23][4] +
                  mat_A[25][24] * mat_B[24][4] +
                  mat_A[25][25] * mat_B[25][4] +
                  mat_A[25][26] * mat_B[26][4] +
                  mat_A[25][27] * mat_B[27][4] +
                  mat_A[25][28] * mat_B[28][4] +
                  mat_A[25][29] * mat_B[29][4] +
                  mat_A[25][30] * mat_B[30][4] +
                  mat_A[25][31] * mat_B[31][4];
    mat_C[25][5] <= 
                  mat_A[25][0] * mat_B[0][5] +
                  mat_A[25][1] * mat_B[1][5] +
                  mat_A[25][2] * mat_B[2][5] +
                  mat_A[25][3] * mat_B[3][5] +
                  mat_A[25][4] * mat_B[4][5] +
                  mat_A[25][5] * mat_B[5][5] +
                  mat_A[25][6] * mat_B[6][5] +
                  mat_A[25][7] * mat_B[7][5] +
                  mat_A[25][8] * mat_B[8][5] +
                  mat_A[25][9] * mat_B[9][5] +
                  mat_A[25][10] * mat_B[10][5] +
                  mat_A[25][11] * mat_B[11][5] +
                  mat_A[25][12] * mat_B[12][5] +
                  mat_A[25][13] * mat_B[13][5] +
                  mat_A[25][14] * mat_B[14][5] +
                  mat_A[25][15] * mat_B[15][5] +
                  mat_A[25][16] * mat_B[16][5] +
                  mat_A[25][17] * mat_B[17][5] +
                  mat_A[25][18] * mat_B[18][5] +
                  mat_A[25][19] * mat_B[19][5] +
                  mat_A[25][20] * mat_B[20][5] +
                  mat_A[25][21] * mat_B[21][5] +
                  mat_A[25][22] * mat_B[22][5] +
                  mat_A[25][23] * mat_B[23][5] +
                  mat_A[25][24] * mat_B[24][5] +
                  mat_A[25][25] * mat_B[25][5] +
                  mat_A[25][26] * mat_B[26][5] +
                  mat_A[25][27] * mat_B[27][5] +
                  mat_A[25][28] * mat_B[28][5] +
                  mat_A[25][29] * mat_B[29][5] +
                  mat_A[25][30] * mat_B[30][5] +
                  mat_A[25][31] * mat_B[31][5];
    mat_C[25][6] <= 
                  mat_A[25][0] * mat_B[0][6] +
                  mat_A[25][1] * mat_B[1][6] +
                  mat_A[25][2] * mat_B[2][6] +
                  mat_A[25][3] * mat_B[3][6] +
                  mat_A[25][4] * mat_B[4][6] +
                  mat_A[25][5] * mat_B[5][6] +
                  mat_A[25][6] * mat_B[6][6] +
                  mat_A[25][7] * mat_B[7][6] +
                  mat_A[25][8] * mat_B[8][6] +
                  mat_A[25][9] * mat_B[9][6] +
                  mat_A[25][10] * mat_B[10][6] +
                  mat_A[25][11] * mat_B[11][6] +
                  mat_A[25][12] * mat_B[12][6] +
                  mat_A[25][13] * mat_B[13][6] +
                  mat_A[25][14] * mat_B[14][6] +
                  mat_A[25][15] * mat_B[15][6] +
                  mat_A[25][16] * mat_B[16][6] +
                  mat_A[25][17] * mat_B[17][6] +
                  mat_A[25][18] * mat_B[18][6] +
                  mat_A[25][19] * mat_B[19][6] +
                  mat_A[25][20] * mat_B[20][6] +
                  mat_A[25][21] * mat_B[21][6] +
                  mat_A[25][22] * mat_B[22][6] +
                  mat_A[25][23] * mat_B[23][6] +
                  mat_A[25][24] * mat_B[24][6] +
                  mat_A[25][25] * mat_B[25][6] +
                  mat_A[25][26] * mat_B[26][6] +
                  mat_A[25][27] * mat_B[27][6] +
                  mat_A[25][28] * mat_B[28][6] +
                  mat_A[25][29] * mat_B[29][6] +
                  mat_A[25][30] * mat_B[30][6] +
                  mat_A[25][31] * mat_B[31][6];
    mat_C[25][7] <= 
                  mat_A[25][0] * mat_B[0][7] +
                  mat_A[25][1] * mat_B[1][7] +
                  mat_A[25][2] * mat_B[2][7] +
                  mat_A[25][3] * mat_B[3][7] +
                  mat_A[25][4] * mat_B[4][7] +
                  mat_A[25][5] * mat_B[5][7] +
                  mat_A[25][6] * mat_B[6][7] +
                  mat_A[25][7] * mat_B[7][7] +
                  mat_A[25][8] * mat_B[8][7] +
                  mat_A[25][9] * mat_B[9][7] +
                  mat_A[25][10] * mat_B[10][7] +
                  mat_A[25][11] * mat_B[11][7] +
                  mat_A[25][12] * mat_B[12][7] +
                  mat_A[25][13] * mat_B[13][7] +
                  mat_A[25][14] * mat_B[14][7] +
                  mat_A[25][15] * mat_B[15][7] +
                  mat_A[25][16] * mat_B[16][7] +
                  mat_A[25][17] * mat_B[17][7] +
                  mat_A[25][18] * mat_B[18][7] +
                  mat_A[25][19] * mat_B[19][7] +
                  mat_A[25][20] * mat_B[20][7] +
                  mat_A[25][21] * mat_B[21][7] +
                  mat_A[25][22] * mat_B[22][7] +
                  mat_A[25][23] * mat_B[23][7] +
                  mat_A[25][24] * mat_B[24][7] +
                  mat_A[25][25] * mat_B[25][7] +
                  mat_A[25][26] * mat_B[26][7] +
                  mat_A[25][27] * mat_B[27][7] +
                  mat_A[25][28] * mat_B[28][7] +
                  mat_A[25][29] * mat_B[29][7] +
                  mat_A[25][30] * mat_B[30][7] +
                  mat_A[25][31] * mat_B[31][7];
    mat_C[25][8] <= 
                  mat_A[25][0] * mat_B[0][8] +
                  mat_A[25][1] * mat_B[1][8] +
                  mat_A[25][2] * mat_B[2][8] +
                  mat_A[25][3] * mat_B[3][8] +
                  mat_A[25][4] * mat_B[4][8] +
                  mat_A[25][5] * mat_B[5][8] +
                  mat_A[25][6] * mat_B[6][8] +
                  mat_A[25][7] * mat_B[7][8] +
                  mat_A[25][8] * mat_B[8][8] +
                  mat_A[25][9] * mat_B[9][8] +
                  mat_A[25][10] * mat_B[10][8] +
                  mat_A[25][11] * mat_B[11][8] +
                  mat_A[25][12] * mat_B[12][8] +
                  mat_A[25][13] * mat_B[13][8] +
                  mat_A[25][14] * mat_B[14][8] +
                  mat_A[25][15] * mat_B[15][8] +
                  mat_A[25][16] * mat_B[16][8] +
                  mat_A[25][17] * mat_B[17][8] +
                  mat_A[25][18] * mat_B[18][8] +
                  mat_A[25][19] * mat_B[19][8] +
                  mat_A[25][20] * mat_B[20][8] +
                  mat_A[25][21] * mat_B[21][8] +
                  mat_A[25][22] * mat_B[22][8] +
                  mat_A[25][23] * mat_B[23][8] +
                  mat_A[25][24] * mat_B[24][8] +
                  mat_A[25][25] * mat_B[25][8] +
                  mat_A[25][26] * mat_B[26][8] +
                  mat_A[25][27] * mat_B[27][8] +
                  mat_A[25][28] * mat_B[28][8] +
                  mat_A[25][29] * mat_B[29][8] +
                  mat_A[25][30] * mat_B[30][8] +
                  mat_A[25][31] * mat_B[31][8];
    mat_C[25][9] <= 
                  mat_A[25][0] * mat_B[0][9] +
                  mat_A[25][1] * mat_B[1][9] +
                  mat_A[25][2] * mat_B[2][9] +
                  mat_A[25][3] * mat_B[3][9] +
                  mat_A[25][4] * mat_B[4][9] +
                  mat_A[25][5] * mat_B[5][9] +
                  mat_A[25][6] * mat_B[6][9] +
                  mat_A[25][7] * mat_B[7][9] +
                  mat_A[25][8] * mat_B[8][9] +
                  mat_A[25][9] * mat_B[9][9] +
                  mat_A[25][10] * mat_B[10][9] +
                  mat_A[25][11] * mat_B[11][9] +
                  mat_A[25][12] * mat_B[12][9] +
                  mat_A[25][13] * mat_B[13][9] +
                  mat_A[25][14] * mat_B[14][9] +
                  mat_A[25][15] * mat_B[15][9] +
                  mat_A[25][16] * mat_B[16][9] +
                  mat_A[25][17] * mat_B[17][9] +
                  mat_A[25][18] * mat_B[18][9] +
                  mat_A[25][19] * mat_B[19][9] +
                  mat_A[25][20] * mat_B[20][9] +
                  mat_A[25][21] * mat_B[21][9] +
                  mat_A[25][22] * mat_B[22][9] +
                  mat_A[25][23] * mat_B[23][9] +
                  mat_A[25][24] * mat_B[24][9] +
                  mat_A[25][25] * mat_B[25][9] +
                  mat_A[25][26] * mat_B[26][9] +
                  mat_A[25][27] * mat_B[27][9] +
                  mat_A[25][28] * mat_B[28][9] +
                  mat_A[25][29] * mat_B[29][9] +
                  mat_A[25][30] * mat_B[30][9] +
                  mat_A[25][31] * mat_B[31][9];
    mat_C[25][10] <= 
                  mat_A[25][0] * mat_B[0][10] +
                  mat_A[25][1] * mat_B[1][10] +
                  mat_A[25][2] * mat_B[2][10] +
                  mat_A[25][3] * mat_B[3][10] +
                  mat_A[25][4] * mat_B[4][10] +
                  mat_A[25][5] * mat_B[5][10] +
                  mat_A[25][6] * mat_B[6][10] +
                  mat_A[25][7] * mat_B[7][10] +
                  mat_A[25][8] * mat_B[8][10] +
                  mat_A[25][9] * mat_B[9][10] +
                  mat_A[25][10] * mat_B[10][10] +
                  mat_A[25][11] * mat_B[11][10] +
                  mat_A[25][12] * mat_B[12][10] +
                  mat_A[25][13] * mat_B[13][10] +
                  mat_A[25][14] * mat_B[14][10] +
                  mat_A[25][15] * mat_B[15][10] +
                  mat_A[25][16] * mat_B[16][10] +
                  mat_A[25][17] * mat_B[17][10] +
                  mat_A[25][18] * mat_B[18][10] +
                  mat_A[25][19] * mat_B[19][10] +
                  mat_A[25][20] * mat_B[20][10] +
                  mat_A[25][21] * mat_B[21][10] +
                  mat_A[25][22] * mat_B[22][10] +
                  mat_A[25][23] * mat_B[23][10] +
                  mat_A[25][24] * mat_B[24][10] +
                  mat_A[25][25] * mat_B[25][10] +
                  mat_A[25][26] * mat_B[26][10] +
                  mat_A[25][27] * mat_B[27][10] +
                  mat_A[25][28] * mat_B[28][10] +
                  mat_A[25][29] * mat_B[29][10] +
                  mat_A[25][30] * mat_B[30][10] +
                  mat_A[25][31] * mat_B[31][10];
    mat_C[25][11] <= 
                  mat_A[25][0] * mat_B[0][11] +
                  mat_A[25][1] * mat_B[1][11] +
                  mat_A[25][2] * mat_B[2][11] +
                  mat_A[25][3] * mat_B[3][11] +
                  mat_A[25][4] * mat_B[4][11] +
                  mat_A[25][5] * mat_B[5][11] +
                  mat_A[25][6] * mat_B[6][11] +
                  mat_A[25][7] * mat_B[7][11] +
                  mat_A[25][8] * mat_B[8][11] +
                  mat_A[25][9] * mat_B[9][11] +
                  mat_A[25][10] * mat_B[10][11] +
                  mat_A[25][11] * mat_B[11][11] +
                  mat_A[25][12] * mat_B[12][11] +
                  mat_A[25][13] * mat_B[13][11] +
                  mat_A[25][14] * mat_B[14][11] +
                  mat_A[25][15] * mat_B[15][11] +
                  mat_A[25][16] * mat_B[16][11] +
                  mat_A[25][17] * mat_B[17][11] +
                  mat_A[25][18] * mat_B[18][11] +
                  mat_A[25][19] * mat_B[19][11] +
                  mat_A[25][20] * mat_B[20][11] +
                  mat_A[25][21] * mat_B[21][11] +
                  mat_A[25][22] * mat_B[22][11] +
                  mat_A[25][23] * mat_B[23][11] +
                  mat_A[25][24] * mat_B[24][11] +
                  mat_A[25][25] * mat_B[25][11] +
                  mat_A[25][26] * mat_B[26][11] +
                  mat_A[25][27] * mat_B[27][11] +
                  mat_A[25][28] * mat_B[28][11] +
                  mat_A[25][29] * mat_B[29][11] +
                  mat_A[25][30] * mat_B[30][11] +
                  mat_A[25][31] * mat_B[31][11];
    mat_C[25][12] <= 
                  mat_A[25][0] * mat_B[0][12] +
                  mat_A[25][1] * mat_B[1][12] +
                  mat_A[25][2] * mat_B[2][12] +
                  mat_A[25][3] * mat_B[3][12] +
                  mat_A[25][4] * mat_B[4][12] +
                  mat_A[25][5] * mat_B[5][12] +
                  mat_A[25][6] * mat_B[6][12] +
                  mat_A[25][7] * mat_B[7][12] +
                  mat_A[25][8] * mat_B[8][12] +
                  mat_A[25][9] * mat_B[9][12] +
                  mat_A[25][10] * mat_B[10][12] +
                  mat_A[25][11] * mat_B[11][12] +
                  mat_A[25][12] * mat_B[12][12] +
                  mat_A[25][13] * mat_B[13][12] +
                  mat_A[25][14] * mat_B[14][12] +
                  mat_A[25][15] * mat_B[15][12] +
                  mat_A[25][16] * mat_B[16][12] +
                  mat_A[25][17] * mat_B[17][12] +
                  mat_A[25][18] * mat_B[18][12] +
                  mat_A[25][19] * mat_B[19][12] +
                  mat_A[25][20] * mat_B[20][12] +
                  mat_A[25][21] * mat_B[21][12] +
                  mat_A[25][22] * mat_B[22][12] +
                  mat_A[25][23] * mat_B[23][12] +
                  mat_A[25][24] * mat_B[24][12] +
                  mat_A[25][25] * mat_B[25][12] +
                  mat_A[25][26] * mat_B[26][12] +
                  mat_A[25][27] * mat_B[27][12] +
                  mat_A[25][28] * mat_B[28][12] +
                  mat_A[25][29] * mat_B[29][12] +
                  mat_A[25][30] * mat_B[30][12] +
                  mat_A[25][31] * mat_B[31][12];
    mat_C[25][13] <= 
                  mat_A[25][0] * mat_B[0][13] +
                  mat_A[25][1] * mat_B[1][13] +
                  mat_A[25][2] * mat_B[2][13] +
                  mat_A[25][3] * mat_B[3][13] +
                  mat_A[25][4] * mat_B[4][13] +
                  mat_A[25][5] * mat_B[5][13] +
                  mat_A[25][6] * mat_B[6][13] +
                  mat_A[25][7] * mat_B[7][13] +
                  mat_A[25][8] * mat_B[8][13] +
                  mat_A[25][9] * mat_B[9][13] +
                  mat_A[25][10] * mat_B[10][13] +
                  mat_A[25][11] * mat_B[11][13] +
                  mat_A[25][12] * mat_B[12][13] +
                  mat_A[25][13] * mat_B[13][13] +
                  mat_A[25][14] * mat_B[14][13] +
                  mat_A[25][15] * mat_B[15][13] +
                  mat_A[25][16] * mat_B[16][13] +
                  mat_A[25][17] * mat_B[17][13] +
                  mat_A[25][18] * mat_B[18][13] +
                  mat_A[25][19] * mat_B[19][13] +
                  mat_A[25][20] * mat_B[20][13] +
                  mat_A[25][21] * mat_B[21][13] +
                  mat_A[25][22] * mat_B[22][13] +
                  mat_A[25][23] * mat_B[23][13] +
                  mat_A[25][24] * mat_B[24][13] +
                  mat_A[25][25] * mat_B[25][13] +
                  mat_A[25][26] * mat_B[26][13] +
                  mat_A[25][27] * mat_B[27][13] +
                  mat_A[25][28] * mat_B[28][13] +
                  mat_A[25][29] * mat_B[29][13] +
                  mat_A[25][30] * mat_B[30][13] +
                  mat_A[25][31] * mat_B[31][13];
    mat_C[25][14] <= 
                  mat_A[25][0] * mat_B[0][14] +
                  mat_A[25][1] * mat_B[1][14] +
                  mat_A[25][2] * mat_B[2][14] +
                  mat_A[25][3] * mat_B[3][14] +
                  mat_A[25][4] * mat_B[4][14] +
                  mat_A[25][5] * mat_B[5][14] +
                  mat_A[25][6] * mat_B[6][14] +
                  mat_A[25][7] * mat_B[7][14] +
                  mat_A[25][8] * mat_B[8][14] +
                  mat_A[25][9] * mat_B[9][14] +
                  mat_A[25][10] * mat_B[10][14] +
                  mat_A[25][11] * mat_B[11][14] +
                  mat_A[25][12] * mat_B[12][14] +
                  mat_A[25][13] * mat_B[13][14] +
                  mat_A[25][14] * mat_B[14][14] +
                  mat_A[25][15] * mat_B[15][14] +
                  mat_A[25][16] * mat_B[16][14] +
                  mat_A[25][17] * mat_B[17][14] +
                  mat_A[25][18] * mat_B[18][14] +
                  mat_A[25][19] * mat_B[19][14] +
                  mat_A[25][20] * mat_B[20][14] +
                  mat_A[25][21] * mat_B[21][14] +
                  mat_A[25][22] * mat_B[22][14] +
                  mat_A[25][23] * mat_B[23][14] +
                  mat_A[25][24] * mat_B[24][14] +
                  mat_A[25][25] * mat_B[25][14] +
                  mat_A[25][26] * mat_B[26][14] +
                  mat_A[25][27] * mat_B[27][14] +
                  mat_A[25][28] * mat_B[28][14] +
                  mat_A[25][29] * mat_B[29][14] +
                  mat_A[25][30] * mat_B[30][14] +
                  mat_A[25][31] * mat_B[31][14];
    mat_C[25][15] <= 
                  mat_A[25][0] * mat_B[0][15] +
                  mat_A[25][1] * mat_B[1][15] +
                  mat_A[25][2] * mat_B[2][15] +
                  mat_A[25][3] * mat_B[3][15] +
                  mat_A[25][4] * mat_B[4][15] +
                  mat_A[25][5] * mat_B[5][15] +
                  mat_A[25][6] * mat_B[6][15] +
                  mat_A[25][7] * mat_B[7][15] +
                  mat_A[25][8] * mat_B[8][15] +
                  mat_A[25][9] * mat_B[9][15] +
                  mat_A[25][10] * mat_B[10][15] +
                  mat_A[25][11] * mat_B[11][15] +
                  mat_A[25][12] * mat_B[12][15] +
                  mat_A[25][13] * mat_B[13][15] +
                  mat_A[25][14] * mat_B[14][15] +
                  mat_A[25][15] * mat_B[15][15] +
                  mat_A[25][16] * mat_B[16][15] +
                  mat_A[25][17] * mat_B[17][15] +
                  mat_A[25][18] * mat_B[18][15] +
                  mat_A[25][19] * mat_B[19][15] +
                  mat_A[25][20] * mat_B[20][15] +
                  mat_A[25][21] * mat_B[21][15] +
                  mat_A[25][22] * mat_B[22][15] +
                  mat_A[25][23] * mat_B[23][15] +
                  mat_A[25][24] * mat_B[24][15] +
                  mat_A[25][25] * mat_B[25][15] +
                  mat_A[25][26] * mat_B[26][15] +
                  mat_A[25][27] * mat_B[27][15] +
                  mat_A[25][28] * mat_B[28][15] +
                  mat_A[25][29] * mat_B[29][15] +
                  mat_A[25][30] * mat_B[30][15] +
                  mat_A[25][31] * mat_B[31][15];
    mat_C[25][16] <= 
                  mat_A[25][0] * mat_B[0][16] +
                  mat_A[25][1] * mat_B[1][16] +
                  mat_A[25][2] * mat_B[2][16] +
                  mat_A[25][3] * mat_B[3][16] +
                  mat_A[25][4] * mat_B[4][16] +
                  mat_A[25][5] * mat_B[5][16] +
                  mat_A[25][6] * mat_B[6][16] +
                  mat_A[25][7] * mat_B[7][16] +
                  mat_A[25][8] * mat_B[8][16] +
                  mat_A[25][9] * mat_B[9][16] +
                  mat_A[25][10] * mat_B[10][16] +
                  mat_A[25][11] * mat_B[11][16] +
                  mat_A[25][12] * mat_B[12][16] +
                  mat_A[25][13] * mat_B[13][16] +
                  mat_A[25][14] * mat_B[14][16] +
                  mat_A[25][15] * mat_B[15][16] +
                  mat_A[25][16] * mat_B[16][16] +
                  mat_A[25][17] * mat_B[17][16] +
                  mat_A[25][18] * mat_B[18][16] +
                  mat_A[25][19] * mat_B[19][16] +
                  mat_A[25][20] * mat_B[20][16] +
                  mat_A[25][21] * mat_B[21][16] +
                  mat_A[25][22] * mat_B[22][16] +
                  mat_A[25][23] * mat_B[23][16] +
                  mat_A[25][24] * mat_B[24][16] +
                  mat_A[25][25] * mat_B[25][16] +
                  mat_A[25][26] * mat_B[26][16] +
                  mat_A[25][27] * mat_B[27][16] +
                  mat_A[25][28] * mat_B[28][16] +
                  mat_A[25][29] * mat_B[29][16] +
                  mat_A[25][30] * mat_B[30][16] +
                  mat_A[25][31] * mat_B[31][16];
    mat_C[25][17] <= 
                  mat_A[25][0] * mat_B[0][17] +
                  mat_A[25][1] * mat_B[1][17] +
                  mat_A[25][2] * mat_B[2][17] +
                  mat_A[25][3] * mat_B[3][17] +
                  mat_A[25][4] * mat_B[4][17] +
                  mat_A[25][5] * mat_B[5][17] +
                  mat_A[25][6] * mat_B[6][17] +
                  mat_A[25][7] * mat_B[7][17] +
                  mat_A[25][8] * mat_B[8][17] +
                  mat_A[25][9] * mat_B[9][17] +
                  mat_A[25][10] * mat_B[10][17] +
                  mat_A[25][11] * mat_B[11][17] +
                  mat_A[25][12] * mat_B[12][17] +
                  mat_A[25][13] * mat_B[13][17] +
                  mat_A[25][14] * mat_B[14][17] +
                  mat_A[25][15] * mat_B[15][17] +
                  mat_A[25][16] * mat_B[16][17] +
                  mat_A[25][17] * mat_B[17][17] +
                  mat_A[25][18] * mat_B[18][17] +
                  mat_A[25][19] * mat_B[19][17] +
                  mat_A[25][20] * mat_B[20][17] +
                  mat_A[25][21] * mat_B[21][17] +
                  mat_A[25][22] * mat_B[22][17] +
                  mat_A[25][23] * mat_B[23][17] +
                  mat_A[25][24] * mat_B[24][17] +
                  mat_A[25][25] * mat_B[25][17] +
                  mat_A[25][26] * mat_B[26][17] +
                  mat_A[25][27] * mat_B[27][17] +
                  mat_A[25][28] * mat_B[28][17] +
                  mat_A[25][29] * mat_B[29][17] +
                  mat_A[25][30] * mat_B[30][17] +
                  mat_A[25][31] * mat_B[31][17];
    mat_C[25][18] <= 
                  mat_A[25][0] * mat_B[0][18] +
                  mat_A[25][1] * mat_B[1][18] +
                  mat_A[25][2] * mat_B[2][18] +
                  mat_A[25][3] * mat_B[3][18] +
                  mat_A[25][4] * mat_B[4][18] +
                  mat_A[25][5] * mat_B[5][18] +
                  mat_A[25][6] * mat_B[6][18] +
                  mat_A[25][7] * mat_B[7][18] +
                  mat_A[25][8] * mat_B[8][18] +
                  mat_A[25][9] * mat_B[9][18] +
                  mat_A[25][10] * mat_B[10][18] +
                  mat_A[25][11] * mat_B[11][18] +
                  mat_A[25][12] * mat_B[12][18] +
                  mat_A[25][13] * mat_B[13][18] +
                  mat_A[25][14] * mat_B[14][18] +
                  mat_A[25][15] * mat_B[15][18] +
                  mat_A[25][16] * mat_B[16][18] +
                  mat_A[25][17] * mat_B[17][18] +
                  mat_A[25][18] * mat_B[18][18] +
                  mat_A[25][19] * mat_B[19][18] +
                  mat_A[25][20] * mat_B[20][18] +
                  mat_A[25][21] * mat_B[21][18] +
                  mat_A[25][22] * mat_B[22][18] +
                  mat_A[25][23] * mat_B[23][18] +
                  mat_A[25][24] * mat_B[24][18] +
                  mat_A[25][25] * mat_B[25][18] +
                  mat_A[25][26] * mat_B[26][18] +
                  mat_A[25][27] * mat_B[27][18] +
                  mat_A[25][28] * mat_B[28][18] +
                  mat_A[25][29] * mat_B[29][18] +
                  mat_A[25][30] * mat_B[30][18] +
                  mat_A[25][31] * mat_B[31][18];
    mat_C[25][19] <= 
                  mat_A[25][0] * mat_B[0][19] +
                  mat_A[25][1] * mat_B[1][19] +
                  mat_A[25][2] * mat_B[2][19] +
                  mat_A[25][3] * mat_B[3][19] +
                  mat_A[25][4] * mat_B[4][19] +
                  mat_A[25][5] * mat_B[5][19] +
                  mat_A[25][6] * mat_B[6][19] +
                  mat_A[25][7] * mat_B[7][19] +
                  mat_A[25][8] * mat_B[8][19] +
                  mat_A[25][9] * mat_B[9][19] +
                  mat_A[25][10] * mat_B[10][19] +
                  mat_A[25][11] * mat_B[11][19] +
                  mat_A[25][12] * mat_B[12][19] +
                  mat_A[25][13] * mat_B[13][19] +
                  mat_A[25][14] * mat_B[14][19] +
                  mat_A[25][15] * mat_B[15][19] +
                  mat_A[25][16] * mat_B[16][19] +
                  mat_A[25][17] * mat_B[17][19] +
                  mat_A[25][18] * mat_B[18][19] +
                  mat_A[25][19] * mat_B[19][19] +
                  mat_A[25][20] * mat_B[20][19] +
                  mat_A[25][21] * mat_B[21][19] +
                  mat_A[25][22] * mat_B[22][19] +
                  mat_A[25][23] * mat_B[23][19] +
                  mat_A[25][24] * mat_B[24][19] +
                  mat_A[25][25] * mat_B[25][19] +
                  mat_A[25][26] * mat_B[26][19] +
                  mat_A[25][27] * mat_B[27][19] +
                  mat_A[25][28] * mat_B[28][19] +
                  mat_A[25][29] * mat_B[29][19] +
                  mat_A[25][30] * mat_B[30][19] +
                  mat_A[25][31] * mat_B[31][19];
    mat_C[25][20] <= 
                  mat_A[25][0] * mat_B[0][20] +
                  mat_A[25][1] * mat_B[1][20] +
                  mat_A[25][2] * mat_B[2][20] +
                  mat_A[25][3] * mat_B[3][20] +
                  mat_A[25][4] * mat_B[4][20] +
                  mat_A[25][5] * mat_B[5][20] +
                  mat_A[25][6] * mat_B[6][20] +
                  mat_A[25][7] * mat_B[7][20] +
                  mat_A[25][8] * mat_B[8][20] +
                  mat_A[25][9] * mat_B[9][20] +
                  mat_A[25][10] * mat_B[10][20] +
                  mat_A[25][11] * mat_B[11][20] +
                  mat_A[25][12] * mat_B[12][20] +
                  mat_A[25][13] * mat_B[13][20] +
                  mat_A[25][14] * mat_B[14][20] +
                  mat_A[25][15] * mat_B[15][20] +
                  mat_A[25][16] * mat_B[16][20] +
                  mat_A[25][17] * mat_B[17][20] +
                  mat_A[25][18] * mat_B[18][20] +
                  mat_A[25][19] * mat_B[19][20] +
                  mat_A[25][20] * mat_B[20][20] +
                  mat_A[25][21] * mat_B[21][20] +
                  mat_A[25][22] * mat_B[22][20] +
                  mat_A[25][23] * mat_B[23][20] +
                  mat_A[25][24] * mat_B[24][20] +
                  mat_A[25][25] * mat_B[25][20] +
                  mat_A[25][26] * mat_B[26][20] +
                  mat_A[25][27] * mat_B[27][20] +
                  mat_A[25][28] * mat_B[28][20] +
                  mat_A[25][29] * mat_B[29][20] +
                  mat_A[25][30] * mat_B[30][20] +
                  mat_A[25][31] * mat_B[31][20];
    mat_C[25][21] <= 
                  mat_A[25][0] * mat_B[0][21] +
                  mat_A[25][1] * mat_B[1][21] +
                  mat_A[25][2] * mat_B[2][21] +
                  mat_A[25][3] * mat_B[3][21] +
                  mat_A[25][4] * mat_B[4][21] +
                  mat_A[25][5] * mat_B[5][21] +
                  mat_A[25][6] * mat_B[6][21] +
                  mat_A[25][7] * mat_B[7][21] +
                  mat_A[25][8] * mat_B[8][21] +
                  mat_A[25][9] * mat_B[9][21] +
                  mat_A[25][10] * mat_B[10][21] +
                  mat_A[25][11] * mat_B[11][21] +
                  mat_A[25][12] * mat_B[12][21] +
                  mat_A[25][13] * mat_B[13][21] +
                  mat_A[25][14] * mat_B[14][21] +
                  mat_A[25][15] * mat_B[15][21] +
                  mat_A[25][16] * mat_B[16][21] +
                  mat_A[25][17] * mat_B[17][21] +
                  mat_A[25][18] * mat_B[18][21] +
                  mat_A[25][19] * mat_B[19][21] +
                  mat_A[25][20] * mat_B[20][21] +
                  mat_A[25][21] * mat_B[21][21] +
                  mat_A[25][22] * mat_B[22][21] +
                  mat_A[25][23] * mat_B[23][21] +
                  mat_A[25][24] * mat_B[24][21] +
                  mat_A[25][25] * mat_B[25][21] +
                  mat_A[25][26] * mat_B[26][21] +
                  mat_A[25][27] * mat_B[27][21] +
                  mat_A[25][28] * mat_B[28][21] +
                  mat_A[25][29] * mat_B[29][21] +
                  mat_A[25][30] * mat_B[30][21] +
                  mat_A[25][31] * mat_B[31][21];
    mat_C[25][22] <= 
                  mat_A[25][0] * mat_B[0][22] +
                  mat_A[25][1] * mat_B[1][22] +
                  mat_A[25][2] * mat_B[2][22] +
                  mat_A[25][3] * mat_B[3][22] +
                  mat_A[25][4] * mat_B[4][22] +
                  mat_A[25][5] * mat_B[5][22] +
                  mat_A[25][6] * mat_B[6][22] +
                  mat_A[25][7] * mat_B[7][22] +
                  mat_A[25][8] * mat_B[8][22] +
                  mat_A[25][9] * mat_B[9][22] +
                  mat_A[25][10] * mat_B[10][22] +
                  mat_A[25][11] * mat_B[11][22] +
                  mat_A[25][12] * mat_B[12][22] +
                  mat_A[25][13] * mat_B[13][22] +
                  mat_A[25][14] * mat_B[14][22] +
                  mat_A[25][15] * mat_B[15][22] +
                  mat_A[25][16] * mat_B[16][22] +
                  mat_A[25][17] * mat_B[17][22] +
                  mat_A[25][18] * mat_B[18][22] +
                  mat_A[25][19] * mat_B[19][22] +
                  mat_A[25][20] * mat_B[20][22] +
                  mat_A[25][21] * mat_B[21][22] +
                  mat_A[25][22] * mat_B[22][22] +
                  mat_A[25][23] * mat_B[23][22] +
                  mat_A[25][24] * mat_B[24][22] +
                  mat_A[25][25] * mat_B[25][22] +
                  mat_A[25][26] * mat_B[26][22] +
                  mat_A[25][27] * mat_B[27][22] +
                  mat_A[25][28] * mat_B[28][22] +
                  mat_A[25][29] * mat_B[29][22] +
                  mat_A[25][30] * mat_B[30][22] +
                  mat_A[25][31] * mat_B[31][22];
    mat_C[25][23] <= 
                  mat_A[25][0] * mat_B[0][23] +
                  mat_A[25][1] * mat_B[1][23] +
                  mat_A[25][2] * mat_B[2][23] +
                  mat_A[25][3] * mat_B[3][23] +
                  mat_A[25][4] * mat_B[4][23] +
                  mat_A[25][5] * mat_B[5][23] +
                  mat_A[25][6] * mat_B[6][23] +
                  mat_A[25][7] * mat_B[7][23] +
                  mat_A[25][8] * mat_B[8][23] +
                  mat_A[25][9] * mat_B[9][23] +
                  mat_A[25][10] * mat_B[10][23] +
                  mat_A[25][11] * mat_B[11][23] +
                  mat_A[25][12] * mat_B[12][23] +
                  mat_A[25][13] * mat_B[13][23] +
                  mat_A[25][14] * mat_B[14][23] +
                  mat_A[25][15] * mat_B[15][23] +
                  mat_A[25][16] * mat_B[16][23] +
                  mat_A[25][17] * mat_B[17][23] +
                  mat_A[25][18] * mat_B[18][23] +
                  mat_A[25][19] * mat_B[19][23] +
                  mat_A[25][20] * mat_B[20][23] +
                  mat_A[25][21] * mat_B[21][23] +
                  mat_A[25][22] * mat_B[22][23] +
                  mat_A[25][23] * mat_B[23][23] +
                  mat_A[25][24] * mat_B[24][23] +
                  mat_A[25][25] * mat_B[25][23] +
                  mat_A[25][26] * mat_B[26][23] +
                  mat_A[25][27] * mat_B[27][23] +
                  mat_A[25][28] * mat_B[28][23] +
                  mat_A[25][29] * mat_B[29][23] +
                  mat_A[25][30] * mat_B[30][23] +
                  mat_A[25][31] * mat_B[31][23];
    mat_C[25][24] <= 
                  mat_A[25][0] * mat_B[0][24] +
                  mat_A[25][1] * mat_B[1][24] +
                  mat_A[25][2] * mat_B[2][24] +
                  mat_A[25][3] * mat_B[3][24] +
                  mat_A[25][4] * mat_B[4][24] +
                  mat_A[25][5] * mat_B[5][24] +
                  mat_A[25][6] * mat_B[6][24] +
                  mat_A[25][7] * mat_B[7][24] +
                  mat_A[25][8] * mat_B[8][24] +
                  mat_A[25][9] * mat_B[9][24] +
                  mat_A[25][10] * mat_B[10][24] +
                  mat_A[25][11] * mat_B[11][24] +
                  mat_A[25][12] * mat_B[12][24] +
                  mat_A[25][13] * mat_B[13][24] +
                  mat_A[25][14] * mat_B[14][24] +
                  mat_A[25][15] * mat_B[15][24] +
                  mat_A[25][16] * mat_B[16][24] +
                  mat_A[25][17] * mat_B[17][24] +
                  mat_A[25][18] * mat_B[18][24] +
                  mat_A[25][19] * mat_B[19][24] +
                  mat_A[25][20] * mat_B[20][24] +
                  mat_A[25][21] * mat_B[21][24] +
                  mat_A[25][22] * mat_B[22][24] +
                  mat_A[25][23] * mat_B[23][24] +
                  mat_A[25][24] * mat_B[24][24] +
                  mat_A[25][25] * mat_B[25][24] +
                  mat_A[25][26] * mat_B[26][24] +
                  mat_A[25][27] * mat_B[27][24] +
                  mat_A[25][28] * mat_B[28][24] +
                  mat_A[25][29] * mat_B[29][24] +
                  mat_A[25][30] * mat_B[30][24] +
                  mat_A[25][31] * mat_B[31][24];
    mat_C[25][25] <= 
                  mat_A[25][0] * mat_B[0][25] +
                  mat_A[25][1] * mat_B[1][25] +
                  mat_A[25][2] * mat_B[2][25] +
                  mat_A[25][3] * mat_B[3][25] +
                  mat_A[25][4] * mat_B[4][25] +
                  mat_A[25][5] * mat_B[5][25] +
                  mat_A[25][6] * mat_B[6][25] +
                  mat_A[25][7] * mat_B[7][25] +
                  mat_A[25][8] * mat_B[8][25] +
                  mat_A[25][9] * mat_B[9][25] +
                  mat_A[25][10] * mat_B[10][25] +
                  mat_A[25][11] * mat_B[11][25] +
                  mat_A[25][12] * mat_B[12][25] +
                  mat_A[25][13] * mat_B[13][25] +
                  mat_A[25][14] * mat_B[14][25] +
                  mat_A[25][15] * mat_B[15][25] +
                  mat_A[25][16] * mat_B[16][25] +
                  mat_A[25][17] * mat_B[17][25] +
                  mat_A[25][18] * mat_B[18][25] +
                  mat_A[25][19] * mat_B[19][25] +
                  mat_A[25][20] * mat_B[20][25] +
                  mat_A[25][21] * mat_B[21][25] +
                  mat_A[25][22] * mat_B[22][25] +
                  mat_A[25][23] * mat_B[23][25] +
                  mat_A[25][24] * mat_B[24][25] +
                  mat_A[25][25] * mat_B[25][25] +
                  mat_A[25][26] * mat_B[26][25] +
                  mat_A[25][27] * mat_B[27][25] +
                  mat_A[25][28] * mat_B[28][25] +
                  mat_A[25][29] * mat_B[29][25] +
                  mat_A[25][30] * mat_B[30][25] +
                  mat_A[25][31] * mat_B[31][25];
    mat_C[25][26] <= 
                  mat_A[25][0] * mat_B[0][26] +
                  mat_A[25][1] * mat_B[1][26] +
                  mat_A[25][2] * mat_B[2][26] +
                  mat_A[25][3] * mat_B[3][26] +
                  mat_A[25][4] * mat_B[4][26] +
                  mat_A[25][5] * mat_B[5][26] +
                  mat_A[25][6] * mat_B[6][26] +
                  mat_A[25][7] * mat_B[7][26] +
                  mat_A[25][8] * mat_B[8][26] +
                  mat_A[25][9] * mat_B[9][26] +
                  mat_A[25][10] * mat_B[10][26] +
                  mat_A[25][11] * mat_B[11][26] +
                  mat_A[25][12] * mat_B[12][26] +
                  mat_A[25][13] * mat_B[13][26] +
                  mat_A[25][14] * mat_B[14][26] +
                  mat_A[25][15] * mat_B[15][26] +
                  mat_A[25][16] * mat_B[16][26] +
                  mat_A[25][17] * mat_B[17][26] +
                  mat_A[25][18] * mat_B[18][26] +
                  mat_A[25][19] * mat_B[19][26] +
                  mat_A[25][20] * mat_B[20][26] +
                  mat_A[25][21] * mat_B[21][26] +
                  mat_A[25][22] * mat_B[22][26] +
                  mat_A[25][23] * mat_B[23][26] +
                  mat_A[25][24] * mat_B[24][26] +
                  mat_A[25][25] * mat_B[25][26] +
                  mat_A[25][26] * mat_B[26][26] +
                  mat_A[25][27] * mat_B[27][26] +
                  mat_A[25][28] * mat_B[28][26] +
                  mat_A[25][29] * mat_B[29][26] +
                  mat_A[25][30] * mat_B[30][26] +
                  mat_A[25][31] * mat_B[31][26];
    mat_C[25][27] <= 
                  mat_A[25][0] * mat_B[0][27] +
                  mat_A[25][1] * mat_B[1][27] +
                  mat_A[25][2] * mat_B[2][27] +
                  mat_A[25][3] * mat_B[3][27] +
                  mat_A[25][4] * mat_B[4][27] +
                  mat_A[25][5] * mat_B[5][27] +
                  mat_A[25][6] * mat_B[6][27] +
                  mat_A[25][7] * mat_B[7][27] +
                  mat_A[25][8] * mat_B[8][27] +
                  mat_A[25][9] * mat_B[9][27] +
                  mat_A[25][10] * mat_B[10][27] +
                  mat_A[25][11] * mat_B[11][27] +
                  mat_A[25][12] * mat_B[12][27] +
                  mat_A[25][13] * mat_B[13][27] +
                  mat_A[25][14] * mat_B[14][27] +
                  mat_A[25][15] * mat_B[15][27] +
                  mat_A[25][16] * mat_B[16][27] +
                  mat_A[25][17] * mat_B[17][27] +
                  mat_A[25][18] * mat_B[18][27] +
                  mat_A[25][19] * mat_B[19][27] +
                  mat_A[25][20] * mat_B[20][27] +
                  mat_A[25][21] * mat_B[21][27] +
                  mat_A[25][22] * mat_B[22][27] +
                  mat_A[25][23] * mat_B[23][27] +
                  mat_A[25][24] * mat_B[24][27] +
                  mat_A[25][25] * mat_B[25][27] +
                  mat_A[25][26] * mat_B[26][27] +
                  mat_A[25][27] * mat_B[27][27] +
                  mat_A[25][28] * mat_B[28][27] +
                  mat_A[25][29] * mat_B[29][27] +
                  mat_A[25][30] * mat_B[30][27] +
                  mat_A[25][31] * mat_B[31][27];
    mat_C[25][28] <= 
                  mat_A[25][0] * mat_B[0][28] +
                  mat_A[25][1] * mat_B[1][28] +
                  mat_A[25][2] * mat_B[2][28] +
                  mat_A[25][3] * mat_B[3][28] +
                  mat_A[25][4] * mat_B[4][28] +
                  mat_A[25][5] * mat_B[5][28] +
                  mat_A[25][6] * mat_B[6][28] +
                  mat_A[25][7] * mat_B[7][28] +
                  mat_A[25][8] * mat_B[8][28] +
                  mat_A[25][9] * mat_B[9][28] +
                  mat_A[25][10] * mat_B[10][28] +
                  mat_A[25][11] * mat_B[11][28] +
                  mat_A[25][12] * mat_B[12][28] +
                  mat_A[25][13] * mat_B[13][28] +
                  mat_A[25][14] * mat_B[14][28] +
                  mat_A[25][15] * mat_B[15][28] +
                  mat_A[25][16] * mat_B[16][28] +
                  mat_A[25][17] * mat_B[17][28] +
                  mat_A[25][18] * mat_B[18][28] +
                  mat_A[25][19] * mat_B[19][28] +
                  mat_A[25][20] * mat_B[20][28] +
                  mat_A[25][21] * mat_B[21][28] +
                  mat_A[25][22] * mat_B[22][28] +
                  mat_A[25][23] * mat_B[23][28] +
                  mat_A[25][24] * mat_B[24][28] +
                  mat_A[25][25] * mat_B[25][28] +
                  mat_A[25][26] * mat_B[26][28] +
                  mat_A[25][27] * mat_B[27][28] +
                  mat_A[25][28] * mat_B[28][28] +
                  mat_A[25][29] * mat_B[29][28] +
                  mat_A[25][30] * mat_B[30][28] +
                  mat_A[25][31] * mat_B[31][28];
    mat_C[25][29] <= 
                  mat_A[25][0] * mat_B[0][29] +
                  mat_A[25][1] * mat_B[1][29] +
                  mat_A[25][2] * mat_B[2][29] +
                  mat_A[25][3] * mat_B[3][29] +
                  mat_A[25][4] * mat_B[4][29] +
                  mat_A[25][5] * mat_B[5][29] +
                  mat_A[25][6] * mat_B[6][29] +
                  mat_A[25][7] * mat_B[7][29] +
                  mat_A[25][8] * mat_B[8][29] +
                  mat_A[25][9] * mat_B[9][29] +
                  mat_A[25][10] * mat_B[10][29] +
                  mat_A[25][11] * mat_B[11][29] +
                  mat_A[25][12] * mat_B[12][29] +
                  mat_A[25][13] * mat_B[13][29] +
                  mat_A[25][14] * mat_B[14][29] +
                  mat_A[25][15] * mat_B[15][29] +
                  mat_A[25][16] * mat_B[16][29] +
                  mat_A[25][17] * mat_B[17][29] +
                  mat_A[25][18] * mat_B[18][29] +
                  mat_A[25][19] * mat_B[19][29] +
                  mat_A[25][20] * mat_B[20][29] +
                  mat_A[25][21] * mat_B[21][29] +
                  mat_A[25][22] * mat_B[22][29] +
                  mat_A[25][23] * mat_B[23][29] +
                  mat_A[25][24] * mat_B[24][29] +
                  mat_A[25][25] * mat_B[25][29] +
                  mat_A[25][26] * mat_B[26][29] +
                  mat_A[25][27] * mat_B[27][29] +
                  mat_A[25][28] * mat_B[28][29] +
                  mat_A[25][29] * mat_B[29][29] +
                  mat_A[25][30] * mat_B[30][29] +
                  mat_A[25][31] * mat_B[31][29];
    mat_C[25][30] <= 
                  mat_A[25][0] * mat_B[0][30] +
                  mat_A[25][1] * mat_B[1][30] +
                  mat_A[25][2] * mat_B[2][30] +
                  mat_A[25][3] * mat_B[3][30] +
                  mat_A[25][4] * mat_B[4][30] +
                  mat_A[25][5] * mat_B[5][30] +
                  mat_A[25][6] * mat_B[6][30] +
                  mat_A[25][7] * mat_B[7][30] +
                  mat_A[25][8] * mat_B[8][30] +
                  mat_A[25][9] * mat_B[9][30] +
                  mat_A[25][10] * mat_B[10][30] +
                  mat_A[25][11] * mat_B[11][30] +
                  mat_A[25][12] * mat_B[12][30] +
                  mat_A[25][13] * mat_B[13][30] +
                  mat_A[25][14] * mat_B[14][30] +
                  mat_A[25][15] * mat_B[15][30] +
                  mat_A[25][16] * mat_B[16][30] +
                  mat_A[25][17] * mat_B[17][30] +
                  mat_A[25][18] * mat_B[18][30] +
                  mat_A[25][19] * mat_B[19][30] +
                  mat_A[25][20] * mat_B[20][30] +
                  mat_A[25][21] * mat_B[21][30] +
                  mat_A[25][22] * mat_B[22][30] +
                  mat_A[25][23] * mat_B[23][30] +
                  mat_A[25][24] * mat_B[24][30] +
                  mat_A[25][25] * mat_B[25][30] +
                  mat_A[25][26] * mat_B[26][30] +
                  mat_A[25][27] * mat_B[27][30] +
                  mat_A[25][28] * mat_B[28][30] +
                  mat_A[25][29] * mat_B[29][30] +
                  mat_A[25][30] * mat_B[30][30] +
                  mat_A[25][31] * mat_B[31][30];
    mat_C[25][31] <= 
                  mat_A[25][0] * mat_B[0][31] +
                  mat_A[25][1] * mat_B[1][31] +
                  mat_A[25][2] * mat_B[2][31] +
                  mat_A[25][3] * mat_B[3][31] +
                  mat_A[25][4] * mat_B[4][31] +
                  mat_A[25][5] * mat_B[5][31] +
                  mat_A[25][6] * mat_B[6][31] +
                  mat_A[25][7] * mat_B[7][31] +
                  mat_A[25][8] * mat_B[8][31] +
                  mat_A[25][9] * mat_B[9][31] +
                  mat_A[25][10] * mat_B[10][31] +
                  mat_A[25][11] * mat_B[11][31] +
                  mat_A[25][12] * mat_B[12][31] +
                  mat_A[25][13] * mat_B[13][31] +
                  mat_A[25][14] * mat_B[14][31] +
                  mat_A[25][15] * mat_B[15][31] +
                  mat_A[25][16] * mat_B[16][31] +
                  mat_A[25][17] * mat_B[17][31] +
                  mat_A[25][18] * mat_B[18][31] +
                  mat_A[25][19] * mat_B[19][31] +
                  mat_A[25][20] * mat_B[20][31] +
                  mat_A[25][21] * mat_B[21][31] +
                  mat_A[25][22] * mat_B[22][31] +
                  mat_A[25][23] * mat_B[23][31] +
                  mat_A[25][24] * mat_B[24][31] +
                  mat_A[25][25] * mat_B[25][31] +
                  mat_A[25][26] * mat_B[26][31] +
                  mat_A[25][27] * mat_B[27][31] +
                  mat_A[25][28] * mat_B[28][31] +
                  mat_A[25][29] * mat_B[29][31] +
                  mat_A[25][30] * mat_B[30][31] +
                  mat_A[25][31] * mat_B[31][31];
    mat_C[26][0] <= 
                  mat_A[26][0] * mat_B[0][0] +
                  mat_A[26][1] * mat_B[1][0] +
                  mat_A[26][2] * mat_B[2][0] +
                  mat_A[26][3] * mat_B[3][0] +
                  mat_A[26][4] * mat_B[4][0] +
                  mat_A[26][5] * mat_B[5][0] +
                  mat_A[26][6] * mat_B[6][0] +
                  mat_A[26][7] * mat_B[7][0] +
                  mat_A[26][8] * mat_B[8][0] +
                  mat_A[26][9] * mat_B[9][0] +
                  mat_A[26][10] * mat_B[10][0] +
                  mat_A[26][11] * mat_B[11][0] +
                  mat_A[26][12] * mat_B[12][0] +
                  mat_A[26][13] * mat_B[13][0] +
                  mat_A[26][14] * mat_B[14][0] +
                  mat_A[26][15] * mat_B[15][0] +
                  mat_A[26][16] * mat_B[16][0] +
                  mat_A[26][17] * mat_B[17][0] +
                  mat_A[26][18] * mat_B[18][0] +
                  mat_A[26][19] * mat_B[19][0] +
                  mat_A[26][20] * mat_B[20][0] +
                  mat_A[26][21] * mat_B[21][0] +
                  mat_A[26][22] * mat_B[22][0] +
                  mat_A[26][23] * mat_B[23][0] +
                  mat_A[26][24] * mat_B[24][0] +
                  mat_A[26][25] * mat_B[25][0] +
                  mat_A[26][26] * mat_B[26][0] +
                  mat_A[26][27] * mat_B[27][0] +
                  mat_A[26][28] * mat_B[28][0] +
                  mat_A[26][29] * mat_B[29][0] +
                  mat_A[26][30] * mat_B[30][0] +
                  mat_A[26][31] * mat_B[31][0];
    mat_C[26][1] <= 
                  mat_A[26][0] * mat_B[0][1] +
                  mat_A[26][1] * mat_B[1][1] +
                  mat_A[26][2] * mat_B[2][1] +
                  mat_A[26][3] * mat_B[3][1] +
                  mat_A[26][4] * mat_B[4][1] +
                  mat_A[26][5] * mat_B[5][1] +
                  mat_A[26][6] * mat_B[6][1] +
                  mat_A[26][7] * mat_B[7][1] +
                  mat_A[26][8] * mat_B[8][1] +
                  mat_A[26][9] * mat_B[9][1] +
                  mat_A[26][10] * mat_B[10][1] +
                  mat_A[26][11] * mat_B[11][1] +
                  mat_A[26][12] * mat_B[12][1] +
                  mat_A[26][13] * mat_B[13][1] +
                  mat_A[26][14] * mat_B[14][1] +
                  mat_A[26][15] * mat_B[15][1] +
                  mat_A[26][16] * mat_B[16][1] +
                  mat_A[26][17] * mat_B[17][1] +
                  mat_A[26][18] * mat_B[18][1] +
                  mat_A[26][19] * mat_B[19][1] +
                  mat_A[26][20] * mat_B[20][1] +
                  mat_A[26][21] * mat_B[21][1] +
                  mat_A[26][22] * mat_B[22][1] +
                  mat_A[26][23] * mat_B[23][1] +
                  mat_A[26][24] * mat_B[24][1] +
                  mat_A[26][25] * mat_B[25][1] +
                  mat_A[26][26] * mat_B[26][1] +
                  mat_A[26][27] * mat_B[27][1] +
                  mat_A[26][28] * mat_B[28][1] +
                  mat_A[26][29] * mat_B[29][1] +
                  mat_A[26][30] * mat_B[30][1] +
                  mat_A[26][31] * mat_B[31][1];
    mat_C[26][2] <= 
                  mat_A[26][0] * mat_B[0][2] +
                  mat_A[26][1] * mat_B[1][2] +
                  mat_A[26][2] * mat_B[2][2] +
                  mat_A[26][3] * mat_B[3][2] +
                  mat_A[26][4] * mat_B[4][2] +
                  mat_A[26][5] * mat_B[5][2] +
                  mat_A[26][6] * mat_B[6][2] +
                  mat_A[26][7] * mat_B[7][2] +
                  mat_A[26][8] * mat_B[8][2] +
                  mat_A[26][9] * mat_B[9][2] +
                  mat_A[26][10] * mat_B[10][2] +
                  mat_A[26][11] * mat_B[11][2] +
                  mat_A[26][12] * mat_B[12][2] +
                  mat_A[26][13] * mat_B[13][2] +
                  mat_A[26][14] * mat_B[14][2] +
                  mat_A[26][15] * mat_B[15][2] +
                  mat_A[26][16] * mat_B[16][2] +
                  mat_A[26][17] * mat_B[17][2] +
                  mat_A[26][18] * mat_B[18][2] +
                  mat_A[26][19] * mat_B[19][2] +
                  mat_A[26][20] * mat_B[20][2] +
                  mat_A[26][21] * mat_B[21][2] +
                  mat_A[26][22] * mat_B[22][2] +
                  mat_A[26][23] * mat_B[23][2] +
                  mat_A[26][24] * mat_B[24][2] +
                  mat_A[26][25] * mat_B[25][2] +
                  mat_A[26][26] * mat_B[26][2] +
                  mat_A[26][27] * mat_B[27][2] +
                  mat_A[26][28] * mat_B[28][2] +
                  mat_A[26][29] * mat_B[29][2] +
                  mat_A[26][30] * mat_B[30][2] +
                  mat_A[26][31] * mat_B[31][2];
    mat_C[26][3] <= 
                  mat_A[26][0] * mat_B[0][3] +
                  mat_A[26][1] * mat_B[1][3] +
                  mat_A[26][2] * mat_B[2][3] +
                  mat_A[26][3] * mat_B[3][3] +
                  mat_A[26][4] * mat_B[4][3] +
                  mat_A[26][5] * mat_B[5][3] +
                  mat_A[26][6] * mat_B[6][3] +
                  mat_A[26][7] * mat_B[7][3] +
                  mat_A[26][8] * mat_B[8][3] +
                  mat_A[26][9] * mat_B[9][3] +
                  mat_A[26][10] * mat_B[10][3] +
                  mat_A[26][11] * mat_B[11][3] +
                  mat_A[26][12] * mat_B[12][3] +
                  mat_A[26][13] * mat_B[13][3] +
                  mat_A[26][14] * mat_B[14][3] +
                  mat_A[26][15] * mat_B[15][3] +
                  mat_A[26][16] * mat_B[16][3] +
                  mat_A[26][17] * mat_B[17][3] +
                  mat_A[26][18] * mat_B[18][3] +
                  mat_A[26][19] * mat_B[19][3] +
                  mat_A[26][20] * mat_B[20][3] +
                  mat_A[26][21] * mat_B[21][3] +
                  mat_A[26][22] * mat_B[22][3] +
                  mat_A[26][23] * mat_B[23][3] +
                  mat_A[26][24] * mat_B[24][3] +
                  mat_A[26][25] * mat_B[25][3] +
                  mat_A[26][26] * mat_B[26][3] +
                  mat_A[26][27] * mat_B[27][3] +
                  mat_A[26][28] * mat_B[28][3] +
                  mat_A[26][29] * mat_B[29][3] +
                  mat_A[26][30] * mat_B[30][3] +
                  mat_A[26][31] * mat_B[31][3];
    mat_C[26][4] <= 
                  mat_A[26][0] * mat_B[0][4] +
                  mat_A[26][1] * mat_B[1][4] +
                  mat_A[26][2] * mat_B[2][4] +
                  mat_A[26][3] * mat_B[3][4] +
                  mat_A[26][4] * mat_B[4][4] +
                  mat_A[26][5] * mat_B[5][4] +
                  mat_A[26][6] * mat_B[6][4] +
                  mat_A[26][7] * mat_B[7][4] +
                  mat_A[26][8] * mat_B[8][4] +
                  mat_A[26][9] * mat_B[9][4] +
                  mat_A[26][10] * mat_B[10][4] +
                  mat_A[26][11] * mat_B[11][4] +
                  mat_A[26][12] * mat_B[12][4] +
                  mat_A[26][13] * mat_B[13][4] +
                  mat_A[26][14] * mat_B[14][4] +
                  mat_A[26][15] * mat_B[15][4] +
                  mat_A[26][16] * mat_B[16][4] +
                  mat_A[26][17] * mat_B[17][4] +
                  mat_A[26][18] * mat_B[18][4] +
                  mat_A[26][19] * mat_B[19][4] +
                  mat_A[26][20] * mat_B[20][4] +
                  mat_A[26][21] * mat_B[21][4] +
                  mat_A[26][22] * mat_B[22][4] +
                  mat_A[26][23] * mat_B[23][4] +
                  mat_A[26][24] * mat_B[24][4] +
                  mat_A[26][25] * mat_B[25][4] +
                  mat_A[26][26] * mat_B[26][4] +
                  mat_A[26][27] * mat_B[27][4] +
                  mat_A[26][28] * mat_B[28][4] +
                  mat_A[26][29] * mat_B[29][4] +
                  mat_A[26][30] * mat_B[30][4] +
                  mat_A[26][31] * mat_B[31][4];
    mat_C[26][5] <= 
                  mat_A[26][0] * mat_B[0][5] +
                  mat_A[26][1] * mat_B[1][5] +
                  mat_A[26][2] * mat_B[2][5] +
                  mat_A[26][3] * mat_B[3][5] +
                  mat_A[26][4] * mat_B[4][5] +
                  mat_A[26][5] * mat_B[5][5] +
                  mat_A[26][6] * mat_B[6][5] +
                  mat_A[26][7] * mat_B[7][5] +
                  mat_A[26][8] * mat_B[8][5] +
                  mat_A[26][9] * mat_B[9][5] +
                  mat_A[26][10] * mat_B[10][5] +
                  mat_A[26][11] * mat_B[11][5] +
                  mat_A[26][12] * mat_B[12][5] +
                  mat_A[26][13] * mat_B[13][5] +
                  mat_A[26][14] * mat_B[14][5] +
                  mat_A[26][15] * mat_B[15][5] +
                  mat_A[26][16] * mat_B[16][5] +
                  mat_A[26][17] * mat_B[17][5] +
                  mat_A[26][18] * mat_B[18][5] +
                  mat_A[26][19] * mat_B[19][5] +
                  mat_A[26][20] * mat_B[20][5] +
                  mat_A[26][21] * mat_B[21][5] +
                  mat_A[26][22] * mat_B[22][5] +
                  mat_A[26][23] * mat_B[23][5] +
                  mat_A[26][24] * mat_B[24][5] +
                  mat_A[26][25] * mat_B[25][5] +
                  mat_A[26][26] * mat_B[26][5] +
                  mat_A[26][27] * mat_B[27][5] +
                  mat_A[26][28] * mat_B[28][5] +
                  mat_A[26][29] * mat_B[29][5] +
                  mat_A[26][30] * mat_B[30][5] +
                  mat_A[26][31] * mat_B[31][5];
    mat_C[26][6] <= 
                  mat_A[26][0] * mat_B[0][6] +
                  mat_A[26][1] * mat_B[1][6] +
                  mat_A[26][2] * mat_B[2][6] +
                  mat_A[26][3] * mat_B[3][6] +
                  mat_A[26][4] * mat_B[4][6] +
                  mat_A[26][5] * mat_B[5][6] +
                  mat_A[26][6] * mat_B[6][6] +
                  mat_A[26][7] * mat_B[7][6] +
                  mat_A[26][8] * mat_B[8][6] +
                  mat_A[26][9] * mat_B[9][6] +
                  mat_A[26][10] * mat_B[10][6] +
                  mat_A[26][11] * mat_B[11][6] +
                  mat_A[26][12] * mat_B[12][6] +
                  mat_A[26][13] * mat_B[13][6] +
                  mat_A[26][14] * mat_B[14][6] +
                  mat_A[26][15] * mat_B[15][6] +
                  mat_A[26][16] * mat_B[16][6] +
                  mat_A[26][17] * mat_B[17][6] +
                  mat_A[26][18] * mat_B[18][6] +
                  mat_A[26][19] * mat_B[19][6] +
                  mat_A[26][20] * mat_B[20][6] +
                  mat_A[26][21] * mat_B[21][6] +
                  mat_A[26][22] * mat_B[22][6] +
                  mat_A[26][23] * mat_B[23][6] +
                  mat_A[26][24] * mat_B[24][6] +
                  mat_A[26][25] * mat_B[25][6] +
                  mat_A[26][26] * mat_B[26][6] +
                  mat_A[26][27] * mat_B[27][6] +
                  mat_A[26][28] * mat_B[28][6] +
                  mat_A[26][29] * mat_B[29][6] +
                  mat_A[26][30] * mat_B[30][6] +
                  mat_A[26][31] * mat_B[31][6];
    mat_C[26][7] <= 
                  mat_A[26][0] * mat_B[0][7] +
                  mat_A[26][1] * mat_B[1][7] +
                  mat_A[26][2] * mat_B[2][7] +
                  mat_A[26][3] * mat_B[3][7] +
                  mat_A[26][4] * mat_B[4][7] +
                  mat_A[26][5] * mat_B[5][7] +
                  mat_A[26][6] * mat_B[6][7] +
                  mat_A[26][7] * mat_B[7][7] +
                  mat_A[26][8] * mat_B[8][7] +
                  mat_A[26][9] * mat_B[9][7] +
                  mat_A[26][10] * mat_B[10][7] +
                  mat_A[26][11] * mat_B[11][7] +
                  mat_A[26][12] * mat_B[12][7] +
                  mat_A[26][13] * mat_B[13][7] +
                  mat_A[26][14] * mat_B[14][7] +
                  mat_A[26][15] * mat_B[15][7] +
                  mat_A[26][16] * mat_B[16][7] +
                  mat_A[26][17] * mat_B[17][7] +
                  mat_A[26][18] * mat_B[18][7] +
                  mat_A[26][19] * mat_B[19][7] +
                  mat_A[26][20] * mat_B[20][7] +
                  mat_A[26][21] * mat_B[21][7] +
                  mat_A[26][22] * mat_B[22][7] +
                  mat_A[26][23] * mat_B[23][7] +
                  mat_A[26][24] * mat_B[24][7] +
                  mat_A[26][25] * mat_B[25][7] +
                  mat_A[26][26] * mat_B[26][7] +
                  mat_A[26][27] * mat_B[27][7] +
                  mat_A[26][28] * mat_B[28][7] +
                  mat_A[26][29] * mat_B[29][7] +
                  mat_A[26][30] * mat_B[30][7] +
                  mat_A[26][31] * mat_B[31][7];
    mat_C[26][8] <= 
                  mat_A[26][0] * mat_B[0][8] +
                  mat_A[26][1] * mat_B[1][8] +
                  mat_A[26][2] * mat_B[2][8] +
                  mat_A[26][3] * mat_B[3][8] +
                  mat_A[26][4] * mat_B[4][8] +
                  mat_A[26][5] * mat_B[5][8] +
                  mat_A[26][6] * mat_B[6][8] +
                  mat_A[26][7] * mat_B[7][8] +
                  mat_A[26][8] * mat_B[8][8] +
                  mat_A[26][9] * mat_B[9][8] +
                  mat_A[26][10] * mat_B[10][8] +
                  mat_A[26][11] * mat_B[11][8] +
                  mat_A[26][12] * mat_B[12][8] +
                  mat_A[26][13] * mat_B[13][8] +
                  mat_A[26][14] * mat_B[14][8] +
                  mat_A[26][15] * mat_B[15][8] +
                  mat_A[26][16] * mat_B[16][8] +
                  mat_A[26][17] * mat_B[17][8] +
                  mat_A[26][18] * mat_B[18][8] +
                  mat_A[26][19] * mat_B[19][8] +
                  mat_A[26][20] * mat_B[20][8] +
                  mat_A[26][21] * mat_B[21][8] +
                  mat_A[26][22] * mat_B[22][8] +
                  mat_A[26][23] * mat_B[23][8] +
                  mat_A[26][24] * mat_B[24][8] +
                  mat_A[26][25] * mat_B[25][8] +
                  mat_A[26][26] * mat_B[26][8] +
                  mat_A[26][27] * mat_B[27][8] +
                  mat_A[26][28] * mat_B[28][8] +
                  mat_A[26][29] * mat_B[29][8] +
                  mat_A[26][30] * mat_B[30][8] +
                  mat_A[26][31] * mat_B[31][8];
    mat_C[26][9] <= 
                  mat_A[26][0] * mat_B[0][9] +
                  mat_A[26][1] * mat_B[1][9] +
                  mat_A[26][2] * mat_B[2][9] +
                  mat_A[26][3] * mat_B[3][9] +
                  mat_A[26][4] * mat_B[4][9] +
                  mat_A[26][5] * mat_B[5][9] +
                  mat_A[26][6] * mat_B[6][9] +
                  mat_A[26][7] * mat_B[7][9] +
                  mat_A[26][8] * mat_B[8][9] +
                  mat_A[26][9] * mat_B[9][9] +
                  mat_A[26][10] * mat_B[10][9] +
                  mat_A[26][11] * mat_B[11][9] +
                  mat_A[26][12] * mat_B[12][9] +
                  mat_A[26][13] * mat_B[13][9] +
                  mat_A[26][14] * mat_B[14][9] +
                  mat_A[26][15] * mat_B[15][9] +
                  mat_A[26][16] * mat_B[16][9] +
                  mat_A[26][17] * mat_B[17][9] +
                  mat_A[26][18] * mat_B[18][9] +
                  mat_A[26][19] * mat_B[19][9] +
                  mat_A[26][20] * mat_B[20][9] +
                  mat_A[26][21] * mat_B[21][9] +
                  mat_A[26][22] * mat_B[22][9] +
                  mat_A[26][23] * mat_B[23][9] +
                  mat_A[26][24] * mat_B[24][9] +
                  mat_A[26][25] * mat_B[25][9] +
                  mat_A[26][26] * mat_B[26][9] +
                  mat_A[26][27] * mat_B[27][9] +
                  mat_A[26][28] * mat_B[28][9] +
                  mat_A[26][29] * mat_B[29][9] +
                  mat_A[26][30] * mat_B[30][9] +
                  mat_A[26][31] * mat_B[31][9];
    mat_C[26][10] <= 
                  mat_A[26][0] * mat_B[0][10] +
                  mat_A[26][1] * mat_B[1][10] +
                  mat_A[26][2] * mat_B[2][10] +
                  mat_A[26][3] * mat_B[3][10] +
                  mat_A[26][4] * mat_B[4][10] +
                  mat_A[26][5] * mat_B[5][10] +
                  mat_A[26][6] * mat_B[6][10] +
                  mat_A[26][7] * mat_B[7][10] +
                  mat_A[26][8] * mat_B[8][10] +
                  mat_A[26][9] * mat_B[9][10] +
                  mat_A[26][10] * mat_B[10][10] +
                  mat_A[26][11] * mat_B[11][10] +
                  mat_A[26][12] * mat_B[12][10] +
                  mat_A[26][13] * mat_B[13][10] +
                  mat_A[26][14] * mat_B[14][10] +
                  mat_A[26][15] * mat_B[15][10] +
                  mat_A[26][16] * mat_B[16][10] +
                  mat_A[26][17] * mat_B[17][10] +
                  mat_A[26][18] * mat_B[18][10] +
                  mat_A[26][19] * mat_B[19][10] +
                  mat_A[26][20] * mat_B[20][10] +
                  mat_A[26][21] * mat_B[21][10] +
                  mat_A[26][22] * mat_B[22][10] +
                  mat_A[26][23] * mat_B[23][10] +
                  mat_A[26][24] * mat_B[24][10] +
                  mat_A[26][25] * mat_B[25][10] +
                  mat_A[26][26] * mat_B[26][10] +
                  mat_A[26][27] * mat_B[27][10] +
                  mat_A[26][28] * mat_B[28][10] +
                  mat_A[26][29] * mat_B[29][10] +
                  mat_A[26][30] * mat_B[30][10] +
                  mat_A[26][31] * mat_B[31][10];
    mat_C[26][11] <= 
                  mat_A[26][0] * mat_B[0][11] +
                  mat_A[26][1] * mat_B[1][11] +
                  mat_A[26][2] * mat_B[2][11] +
                  mat_A[26][3] * mat_B[3][11] +
                  mat_A[26][4] * mat_B[4][11] +
                  mat_A[26][5] * mat_B[5][11] +
                  mat_A[26][6] * mat_B[6][11] +
                  mat_A[26][7] * mat_B[7][11] +
                  mat_A[26][8] * mat_B[8][11] +
                  mat_A[26][9] * mat_B[9][11] +
                  mat_A[26][10] * mat_B[10][11] +
                  mat_A[26][11] * mat_B[11][11] +
                  mat_A[26][12] * mat_B[12][11] +
                  mat_A[26][13] * mat_B[13][11] +
                  mat_A[26][14] * mat_B[14][11] +
                  mat_A[26][15] * mat_B[15][11] +
                  mat_A[26][16] * mat_B[16][11] +
                  mat_A[26][17] * mat_B[17][11] +
                  mat_A[26][18] * mat_B[18][11] +
                  mat_A[26][19] * mat_B[19][11] +
                  mat_A[26][20] * mat_B[20][11] +
                  mat_A[26][21] * mat_B[21][11] +
                  mat_A[26][22] * mat_B[22][11] +
                  mat_A[26][23] * mat_B[23][11] +
                  mat_A[26][24] * mat_B[24][11] +
                  mat_A[26][25] * mat_B[25][11] +
                  mat_A[26][26] * mat_B[26][11] +
                  mat_A[26][27] * mat_B[27][11] +
                  mat_A[26][28] * mat_B[28][11] +
                  mat_A[26][29] * mat_B[29][11] +
                  mat_A[26][30] * mat_B[30][11] +
                  mat_A[26][31] * mat_B[31][11];
    mat_C[26][12] <= 
                  mat_A[26][0] * mat_B[0][12] +
                  mat_A[26][1] * mat_B[1][12] +
                  mat_A[26][2] * mat_B[2][12] +
                  mat_A[26][3] * mat_B[3][12] +
                  mat_A[26][4] * mat_B[4][12] +
                  mat_A[26][5] * mat_B[5][12] +
                  mat_A[26][6] * mat_B[6][12] +
                  mat_A[26][7] * mat_B[7][12] +
                  mat_A[26][8] * mat_B[8][12] +
                  mat_A[26][9] * mat_B[9][12] +
                  mat_A[26][10] * mat_B[10][12] +
                  mat_A[26][11] * mat_B[11][12] +
                  mat_A[26][12] * mat_B[12][12] +
                  mat_A[26][13] * mat_B[13][12] +
                  mat_A[26][14] * mat_B[14][12] +
                  mat_A[26][15] * mat_B[15][12] +
                  mat_A[26][16] * mat_B[16][12] +
                  mat_A[26][17] * mat_B[17][12] +
                  mat_A[26][18] * mat_B[18][12] +
                  mat_A[26][19] * mat_B[19][12] +
                  mat_A[26][20] * mat_B[20][12] +
                  mat_A[26][21] * mat_B[21][12] +
                  mat_A[26][22] * mat_B[22][12] +
                  mat_A[26][23] * mat_B[23][12] +
                  mat_A[26][24] * mat_B[24][12] +
                  mat_A[26][25] * mat_B[25][12] +
                  mat_A[26][26] * mat_B[26][12] +
                  mat_A[26][27] * mat_B[27][12] +
                  mat_A[26][28] * mat_B[28][12] +
                  mat_A[26][29] * mat_B[29][12] +
                  mat_A[26][30] * mat_B[30][12] +
                  mat_A[26][31] * mat_B[31][12];
    mat_C[26][13] <= 
                  mat_A[26][0] * mat_B[0][13] +
                  mat_A[26][1] * mat_B[1][13] +
                  mat_A[26][2] * mat_B[2][13] +
                  mat_A[26][3] * mat_B[3][13] +
                  mat_A[26][4] * mat_B[4][13] +
                  mat_A[26][5] * mat_B[5][13] +
                  mat_A[26][6] * mat_B[6][13] +
                  mat_A[26][7] * mat_B[7][13] +
                  mat_A[26][8] * mat_B[8][13] +
                  mat_A[26][9] * mat_B[9][13] +
                  mat_A[26][10] * mat_B[10][13] +
                  mat_A[26][11] * mat_B[11][13] +
                  mat_A[26][12] * mat_B[12][13] +
                  mat_A[26][13] * mat_B[13][13] +
                  mat_A[26][14] * mat_B[14][13] +
                  mat_A[26][15] * mat_B[15][13] +
                  mat_A[26][16] * mat_B[16][13] +
                  mat_A[26][17] * mat_B[17][13] +
                  mat_A[26][18] * mat_B[18][13] +
                  mat_A[26][19] * mat_B[19][13] +
                  mat_A[26][20] * mat_B[20][13] +
                  mat_A[26][21] * mat_B[21][13] +
                  mat_A[26][22] * mat_B[22][13] +
                  mat_A[26][23] * mat_B[23][13] +
                  mat_A[26][24] * mat_B[24][13] +
                  mat_A[26][25] * mat_B[25][13] +
                  mat_A[26][26] * mat_B[26][13] +
                  mat_A[26][27] * mat_B[27][13] +
                  mat_A[26][28] * mat_B[28][13] +
                  mat_A[26][29] * mat_B[29][13] +
                  mat_A[26][30] * mat_B[30][13] +
                  mat_A[26][31] * mat_B[31][13];
    mat_C[26][14] <= 
                  mat_A[26][0] * mat_B[0][14] +
                  mat_A[26][1] * mat_B[1][14] +
                  mat_A[26][2] * mat_B[2][14] +
                  mat_A[26][3] * mat_B[3][14] +
                  mat_A[26][4] * mat_B[4][14] +
                  mat_A[26][5] * mat_B[5][14] +
                  mat_A[26][6] * mat_B[6][14] +
                  mat_A[26][7] * mat_B[7][14] +
                  mat_A[26][8] * mat_B[8][14] +
                  mat_A[26][9] * mat_B[9][14] +
                  mat_A[26][10] * mat_B[10][14] +
                  mat_A[26][11] * mat_B[11][14] +
                  mat_A[26][12] * mat_B[12][14] +
                  mat_A[26][13] * mat_B[13][14] +
                  mat_A[26][14] * mat_B[14][14] +
                  mat_A[26][15] * mat_B[15][14] +
                  mat_A[26][16] * mat_B[16][14] +
                  mat_A[26][17] * mat_B[17][14] +
                  mat_A[26][18] * mat_B[18][14] +
                  mat_A[26][19] * mat_B[19][14] +
                  mat_A[26][20] * mat_B[20][14] +
                  mat_A[26][21] * mat_B[21][14] +
                  mat_A[26][22] * mat_B[22][14] +
                  mat_A[26][23] * mat_B[23][14] +
                  mat_A[26][24] * mat_B[24][14] +
                  mat_A[26][25] * mat_B[25][14] +
                  mat_A[26][26] * mat_B[26][14] +
                  mat_A[26][27] * mat_B[27][14] +
                  mat_A[26][28] * mat_B[28][14] +
                  mat_A[26][29] * mat_B[29][14] +
                  mat_A[26][30] * mat_B[30][14] +
                  mat_A[26][31] * mat_B[31][14];
    mat_C[26][15] <= 
                  mat_A[26][0] * mat_B[0][15] +
                  mat_A[26][1] * mat_B[1][15] +
                  mat_A[26][2] * mat_B[2][15] +
                  mat_A[26][3] * mat_B[3][15] +
                  mat_A[26][4] * mat_B[4][15] +
                  mat_A[26][5] * mat_B[5][15] +
                  mat_A[26][6] * mat_B[6][15] +
                  mat_A[26][7] * mat_B[7][15] +
                  mat_A[26][8] * mat_B[8][15] +
                  mat_A[26][9] * mat_B[9][15] +
                  mat_A[26][10] * mat_B[10][15] +
                  mat_A[26][11] * mat_B[11][15] +
                  mat_A[26][12] * mat_B[12][15] +
                  mat_A[26][13] * mat_B[13][15] +
                  mat_A[26][14] * mat_B[14][15] +
                  mat_A[26][15] * mat_B[15][15] +
                  mat_A[26][16] * mat_B[16][15] +
                  mat_A[26][17] * mat_B[17][15] +
                  mat_A[26][18] * mat_B[18][15] +
                  mat_A[26][19] * mat_B[19][15] +
                  mat_A[26][20] * mat_B[20][15] +
                  mat_A[26][21] * mat_B[21][15] +
                  mat_A[26][22] * mat_B[22][15] +
                  mat_A[26][23] * mat_B[23][15] +
                  mat_A[26][24] * mat_B[24][15] +
                  mat_A[26][25] * mat_B[25][15] +
                  mat_A[26][26] * mat_B[26][15] +
                  mat_A[26][27] * mat_B[27][15] +
                  mat_A[26][28] * mat_B[28][15] +
                  mat_A[26][29] * mat_B[29][15] +
                  mat_A[26][30] * mat_B[30][15] +
                  mat_A[26][31] * mat_B[31][15];
    mat_C[26][16] <= 
                  mat_A[26][0] * mat_B[0][16] +
                  mat_A[26][1] * mat_B[1][16] +
                  mat_A[26][2] * mat_B[2][16] +
                  mat_A[26][3] * mat_B[3][16] +
                  mat_A[26][4] * mat_B[4][16] +
                  mat_A[26][5] * mat_B[5][16] +
                  mat_A[26][6] * mat_B[6][16] +
                  mat_A[26][7] * mat_B[7][16] +
                  mat_A[26][8] * mat_B[8][16] +
                  mat_A[26][9] * mat_B[9][16] +
                  mat_A[26][10] * mat_B[10][16] +
                  mat_A[26][11] * mat_B[11][16] +
                  mat_A[26][12] * mat_B[12][16] +
                  mat_A[26][13] * mat_B[13][16] +
                  mat_A[26][14] * mat_B[14][16] +
                  mat_A[26][15] * mat_B[15][16] +
                  mat_A[26][16] * mat_B[16][16] +
                  mat_A[26][17] * mat_B[17][16] +
                  mat_A[26][18] * mat_B[18][16] +
                  mat_A[26][19] * mat_B[19][16] +
                  mat_A[26][20] * mat_B[20][16] +
                  mat_A[26][21] * mat_B[21][16] +
                  mat_A[26][22] * mat_B[22][16] +
                  mat_A[26][23] * mat_B[23][16] +
                  mat_A[26][24] * mat_B[24][16] +
                  mat_A[26][25] * mat_B[25][16] +
                  mat_A[26][26] * mat_B[26][16] +
                  mat_A[26][27] * mat_B[27][16] +
                  mat_A[26][28] * mat_B[28][16] +
                  mat_A[26][29] * mat_B[29][16] +
                  mat_A[26][30] * mat_B[30][16] +
                  mat_A[26][31] * mat_B[31][16];
    mat_C[26][17] <= 
                  mat_A[26][0] * mat_B[0][17] +
                  mat_A[26][1] * mat_B[1][17] +
                  mat_A[26][2] * mat_B[2][17] +
                  mat_A[26][3] * mat_B[3][17] +
                  mat_A[26][4] * mat_B[4][17] +
                  mat_A[26][5] * mat_B[5][17] +
                  mat_A[26][6] * mat_B[6][17] +
                  mat_A[26][7] * mat_B[7][17] +
                  mat_A[26][8] * mat_B[8][17] +
                  mat_A[26][9] * mat_B[9][17] +
                  mat_A[26][10] * mat_B[10][17] +
                  mat_A[26][11] * mat_B[11][17] +
                  mat_A[26][12] * mat_B[12][17] +
                  mat_A[26][13] * mat_B[13][17] +
                  mat_A[26][14] * mat_B[14][17] +
                  mat_A[26][15] * mat_B[15][17] +
                  mat_A[26][16] * mat_B[16][17] +
                  mat_A[26][17] * mat_B[17][17] +
                  mat_A[26][18] * mat_B[18][17] +
                  mat_A[26][19] * mat_B[19][17] +
                  mat_A[26][20] * mat_B[20][17] +
                  mat_A[26][21] * mat_B[21][17] +
                  mat_A[26][22] * mat_B[22][17] +
                  mat_A[26][23] * mat_B[23][17] +
                  mat_A[26][24] * mat_B[24][17] +
                  mat_A[26][25] * mat_B[25][17] +
                  mat_A[26][26] * mat_B[26][17] +
                  mat_A[26][27] * mat_B[27][17] +
                  mat_A[26][28] * mat_B[28][17] +
                  mat_A[26][29] * mat_B[29][17] +
                  mat_A[26][30] * mat_B[30][17] +
                  mat_A[26][31] * mat_B[31][17];
    mat_C[26][18] <= 
                  mat_A[26][0] * mat_B[0][18] +
                  mat_A[26][1] * mat_B[1][18] +
                  mat_A[26][2] * mat_B[2][18] +
                  mat_A[26][3] * mat_B[3][18] +
                  mat_A[26][4] * mat_B[4][18] +
                  mat_A[26][5] * mat_B[5][18] +
                  mat_A[26][6] * mat_B[6][18] +
                  mat_A[26][7] * mat_B[7][18] +
                  mat_A[26][8] * mat_B[8][18] +
                  mat_A[26][9] * mat_B[9][18] +
                  mat_A[26][10] * mat_B[10][18] +
                  mat_A[26][11] * mat_B[11][18] +
                  mat_A[26][12] * mat_B[12][18] +
                  mat_A[26][13] * mat_B[13][18] +
                  mat_A[26][14] * mat_B[14][18] +
                  mat_A[26][15] * mat_B[15][18] +
                  mat_A[26][16] * mat_B[16][18] +
                  mat_A[26][17] * mat_B[17][18] +
                  mat_A[26][18] * mat_B[18][18] +
                  mat_A[26][19] * mat_B[19][18] +
                  mat_A[26][20] * mat_B[20][18] +
                  mat_A[26][21] * mat_B[21][18] +
                  mat_A[26][22] * mat_B[22][18] +
                  mat_A[26][23] * mat_B[23][18] +
                  mat_A[26][24] * mat_B[24][18] +
                  mat_A[26][25] * mat_B[25][18] +
                  mat_A[26][26] * mat_B[26][18] +
                  mat_A[26][27] * mat_B[27][18] +
                  mat_A[26][28] * mat_B[28][18] +
                  mat_A[26][29] * mat_B[29][18] +
                  mat_A[26][30] * mat_B[30][18] +
                  mat_A[26][31] * mat_B[31][18];
    mat_C[26][19] <= 
                  mat_A[26][0] * mat_B[0][19] +
                  mat_A[26][1] * mat_B[1][19] +
                  mat_A[26][2] * mat_B[2][19] +
                  mat_A[26][3] * mat_B[3][19] +
                  mat_A[26][4] * mat_B[4][19] +
                  mat_A[26][5] * mat_B[5][19] +
                  mat_A[26][6] * mat_B[6][19] +
                  mat_A[26][7] * mat_B[7][19] +
                  mat_A[26][8] * mat_B[8][19] +
                  mat_A[26][9] * mat_B[9][19] +
                  mat_A[26][10] * mat_B[10][19] +
                  mat_A[26][11] * mat_B[11][19] +
                  mat_A[26][12] * mat_B[12][19] +
                  mat_A[26][13] * mat_B[13][19] +
                  mat_A[26][14] * mat_B[14][19] +
                  mat_A[26][15] * mat_B[15][19] +
                  mat_A[26][16] * mat_B[16][19] +
                  mat_A[26][17] * mat_B[17][19] +
                  mat_A[26][18] * mat_B[18][19] +
                  mat_A[26][19] * mat_B[19][19] +
                  mat_A[26][20] * mat_B[20][19] +
                  mat_A[26][21] * mat_B[21][19] +
                  mat_A[26][22] * mat_B[22][19] +
                  mat_A[26][23] * mat_B[23][19] +
                  mat_A[26][24] * mat_B[24][19] +
                  mat_A[26][25] * mat_B[25][19] +
                  mat_A[26][26] * mat_B[26][19] +
                  mat_A[26][27] * mat_B[27][19] +
                  mat_A[26][28] * mat_B[28][19] +
                  mat_A[26][29] * mat_B[29][19] +
                  mat_A[26][30] * mat_B[30][19] +
                  mat_A[26][31] * mat_B[31][19];
    mat_C[26][20] <= 
                  mat_A[26][0] * mat_B[0][20] +
                  mat_A[26][1] * mat_B[1][20] +
                  mat_A[26][2] * mat_B[2][20] +
                  mat_A[26][3] * mat_B[3][20] +
                  mat_A[26][4] * mat_B[4][20] +
                  mat_A[26][5] * mat_B[5][20] +
                  mat_A[26][6] * mat_B[6][20] +
                  mat_A[26][7] * mat_B[7][20] +
                  mat_A[26][8] * mat_B[8][20] +
                  mat_A[26][9] * mat_B[9][20] +
                  mat_A[26][10] * mat_B[10][20] +
                  mat_A[26][11] * mat_B[11][20] +
                  mat_A[26][12] * mat_B[12][20] +
                  mat_A[26][13] * mat_B[13][20] +
                  mat_A[26][14] * mat_B[14][20] +
                  mat_A[26][15] * mat_B[15][20] +
                  mat_A[26][16] * mat_B[16][20] +
                  mat_A[26][17] * mat_B[17][20] +
                  mat_A[26][18] * mat_B[18][20] +
                  mat_A[26][19] * mat_B[19][20] +
                  mat_A[26][20] * mat_B[20][20] +
                  mat_A[26][21] * mat_B[21][20] +
                  mat_A[26][22] * mat_B[22][20] +
                  mat_A[26][23] * mat_B[23][20] +
                  mat_A[26][24] * mat_B[24][20] +
                  mat_A[26][25] * mat_B[25][20] +
                  mat_A[26][26] * mat_B[26][20] +
                  mat_A[26][27] * mat_B[27][20] +
                  mat_A[26][28] * mat_B[28][20] +
                  mat_A[26][29] * mat_B[29][20] +
                  mat_A[26][30] * mat_B[30][20] +
                  mat_A[26][31] * mat_B[31][20];
    mat_C[26][21] <= 
                  mat_A[26][0] * mat_B[0][21] +
                  mat_A[26][1] * mat_B[1][21] +
                  mat_A[26][2] * mat_B[2][21] +
                  mat_A[26][3] * mat_B[3][21] +
                  mat_A[26][4] * mat_B[4][21] +
                  mat_A[26][5] * mat_B[5][21] +
                  mat_A[26][6] * mat_B[6][21] +
                  mat_A[26][7] * mat_B[7][21] +
                  mat_A[26][8] * mat_B[8][21] +
                  mat_A[26][9] * mat_B[9][21] +
                  mat_A[26][10] * mat_B[10][21] +
                  mat_A[26][11] * mat_B[11][21] +
                  mat_A[26][12] * mat_B[12][21] +
                  mat_A[26][13] * mat_B[13][21] +
                  mat_A[26][14] * mat_B[14][21] +
                  mat_A[26][15] * mat_B[15][21] +
                  mat_A[26][16] * mat_B[16][21] +
                  mat_A[26][17] * mat_B[17][21] +
                  mat_A[26][18] * mat_B[18][21] +
                  mat_A[26][19] * mat_B[19][21] +
                  mat_A[26][20] * mat_B[20][21] +
                  mat_A[26][21] * mat_B[21][21] +
                  mat_A[26][22] * mat_B[22][21] +
                  mat_A[26][23] * mat_B[23][21] +
                  mat_A[26][24] * mat_B[24][21] +
                  mat_A[26][25] * mat_B[25][21] +
                  mat_A[26][26] * mat_B[26][21] +
                  mat_A[26][27] * mat_B[27][21] +
                  mat_A[26][28] * mat_B[28][21] +
                  mat_A[26][29] * mat_B[29][21] +
                  mat_A[26][30] * mat_B[30][21] +
                  mat_A[26][31] * mat_B[31][21];
    mat_C[26][22] <= 
                  mat_A[26][0] * mat_B[0][22] +
                  mat_A[26][1] * mat_B[1][22] +
                  mat_A[26][2] * mat_B[2][22] +
                  mat_A[26][3] * mat_B[3][22] +
                  mat_A[26][4] * mat_B[4][22] +
                  mat_A[26][5] * mat_B[5][22] +
                  mat_A[26][6] * mat_B[6][22] +
                  mat_A[26][7] * mat_B[7][22] +
                  mat_A[26][8] * mat_B[8][22] +
                  mat_A[26][9] * mat_B[9][22] +
                  mat_A[26][10] * mat_B[10][22] +
                  mat_A[26][11] * mat_B[11][22] +
                  mat_A[26][12] * mat_B[12][22] +
                  mat_A[26][13] * mat_B[13][22] +
                  mat_A[26][14] * mat_B[14][22] +
                  mat_A[26][15] * mat_B[15][22] +
                  mat_A[26][16] * mat_B[16][22] +
                  mat_A[26][17] * mat_B[17][22] +
                  mat_A[26][18] * mat_B[18][22] +
                  mat_A[26][19] * mat_B[19][22] +
                  mat_A[26][20] * mat_B[20][22] +
                  mat_A[26][21] * mat_B[21][22] +
                  mat_A[26][22] * mat_B[22][22] +
                  mat_A[26][23] * mat_B[23][22] +
                  mat_A[26][24] * mat_B[24][22] +
                  mat_A[26][25] * mat_B[25][22] +
                  mat_A[26][26] * mat_B[26][22] +
                  mat_A[26][27] * mat_B[27][22] +
                  mat_A[26][28] * mat_B[28][22] +
                  mat_A[26][29] * mat_B[29][22] +
                  mat_A[26][30] * mat_B[30][22] +
                  mat_A[26][31] * mat_B[31][22];
    mat_C[26][23] <= 
                  mat_A[26][0] * mat_B[0][23] +
                  mat_A[26][1] * mat_B[1][23] +
                  mat_A[26][2] * mat_B[2][23] +
                  mat_A[26][3] * mat_B[3][23] +
                  mat_A[26][4] * mat_B[4][23] +
                  mat_A[26][5] * mat_B[5][23] +
                  mat_A[26][6] * mat_B[6][23] +
                  mat_A[26][7] * mat_B[7][23] +
                  mat_A[26][8] * mat_B[8][23] +
                  mat_A[26][9] * mat_B[9][23] +
                  mat_A[26][10] * mat_B[10][23] +
                  mat_A[26][11] * mat_B[11][23] +
                  mat_A[26][12] * mat_B[12][23] +
                  mat_A[26][13] * mat_B[13][23] +
                  mat_A[26][14] * mat_B[14][23] +
                  mat_A[26][15] * mat_B[15][23] +
                  mat_A[26][16] * mat_B[16][23] +
                  mat_A[26][17] * mat_B[17][23] +
                  mat_A[26][18] * mat_B[18][23] +
                  mat_A[26][19] * mat_B[19][23] +
                  mat_A[26][20] * mat_B[20][23] +
                  mat_A[26][21] * mat_B[21][23] +
                  mat_A[26][22] * mat_B[22][23] +
                  mat_A[26][23] * mat_B[23][23] +
                  mat_A[26][24] * mat_B[24][23] +
                  mat_A[26][25] * mat_B[25][23] +
                  mat_A[26][26] * mat_B[26][23] +
                  mat_A[26][27] * mat_B[27][23] +
                  mat_A[26][28] * mat_B[28][23] +
                  mat_A[26][29] * mat_B[29][23] +
                  mat_A[26][30] * mat_B[30][23] +
                  mat_A[26][31] * mat_B[31][23];
    mat_C[26][24] <= 
                  mat_A[26][0] * mat_B[0][24] +
                  mat_A[26][1] * mat_B[1][24] +
                  mat_A[26][2] * mat_B[2][24] +
                  mat_A[26][3] * mat_B[3][24] +
                  mat_A[26][4] * mat_B[4][24] +
                  mat_A[26][5] * mat_B[5][24] +
                  mat_A[26][6] * mat_B[6][24] +
                  mat_A[26][7] * mat_B[7][24] +
                  mat_A[26][8] * mat_B[8][24] +
                  mat_A[26][9] * mat_B[9][24] +
                  mat_A[26][10] * mat_B[10][24] +
                  mat_A[26][11] * mat_B[11][24] +
                  mat_A[26][12] * mat_B[12][24] +
                  mat_A[26][13] * mat_B[13][24] +
                  mat_A[26][14] * mat_B[14][24] +
                  mat_A[26][15] * mat_B[15][24] +
                  mat_A[26][16] * mat_B[16][24] +
                  mat_A[26][17] * mat_B[17][24] +
                  mat_A[26][18] * mat_B[18][24] +
                  mat_A[26][19] * mat_B[19][24] +
                  mat_A[26][20] * mat_B[20][24] +
                  mat_A[26][21] * mat_B[21][24] +
                  mat_A[26][22] * mat_B[22][24] +
                  mat_A[26][23] * mat_B[23][24] +
                  mat_A[26][24] * mat_B[24][24] +
                  mat_A[26][25] * mat_B[25][24] +
                  mat_A[26][26] * mat_B[26][24] +
                  mat_A[26][27] * mat_B[27][24] +
                  mat_A[26][28] * mat_B[28][24] +
                  mat_A[26][29] * mat_B[29][24] +
                  mat_A[26][30] * mat_B[30][24] +
                  mat_A[26][31] * mat_B[31][24];
    mat_C[26][25] <= 
                  mat_A[26][0] * mat_B[0][25] +
                  mat_A[26][1] * mat_B[1][25] +
                  mat_A[26][2] * mat_B[2][25] +
                  mat_A[26][3] * mat_B[3][25] +
                  mat_A[26][4] * mat_B[4][25] +
                  mat_A[26][5] * mat_B[5][25] +
                  mat_A[26][6] * mat_B[6][25] +
                  mat_A[26][7] * mat_B[7][25] +
                  mat_A[26][8] * mat_B[8][25] +
                  mat_A[26][9] * mat_B[9][25] +
                  mat_A[26][10] * mat_B[10][25] +
                  mat_A[26][11] * mat_B[11][25] +
                  mat_A[26][12] * mat_B[12][25] +
                  mat_A[26][13] * mat_B[13][25] +
                  mat_A[26][14] * mat_B[14][25] +
                  mat_A[26][15] * mat_B[15][25] +
                  mat_A[26][16] * mat_B[16][25] +
                  mat_A[26][17] * mat_B[17][25] +
                  mat_A[26][18] * mat_B[18][25] +
                  mat_A[26][19] * mat_B[19][25] +
                  mat_A[26][20] * mat_B[20][25] +
                  mat_A[26][21] * mat_B[21][25] +
                  mat_A[26][22] * mat_B[22][25] +
                  mat_A[26][23] * mat_B[23][25] +
                  mat_A[26][24] * mat_B[24][25] +
                  mat_A[26][25] * mat_B[25][25] +
                  mat_A[26][26] * mat_B[26][25] +
                  mat_A[26][27] * mat_B[27][25] +
                  mat_A[26][28] * mat_B[28][25] +
                  mat_A[26][29] * mat_B[29][25] +
                  mat_A[26][30] * mat_B[30][25] +
                  mat_A[26][31] * mat_B[31][25];
    mat_C[26][26] <= 
                  mat_A[26][0] * mat_B[0][26] +
                  mat_A[26][1] * mat_B[1][26] +
                  mat_A[26][2] * mat_B[2][26] +
                  mat_A[26][3] * mat_B[3][26] +
                  mat_A[26][4] * mat_B[4][26] +
                  mat_A[26][5] * mat_B[5][26] +
                  mat_A[26][6] * mat_B[6][26] +
                  mat_A[26][7] * mat_B[7][26] +
                  mat_A[26][8] * mat_B[8][26] +
                  mat_A[26][9] * mat_B[9][26] +
                  mat_A[26][10] * mat_B[10][26] +
                  mat_A[26][11] * mat_B[11][26] +
                  mat_A[26][12] * mat_B[12][26] +
                  mat_A[26][13] * mat_B[13][26] +
                  mat_A[26][14] * mat_B[14][26] +
                  mat_A[26][15] * mat_B[15][26] +
                  mat_A[26][16] * mat_B[16][26] +
                  mat_A[26][17] * mat_B[17][26] +
                  mat_A[26][18] * mat_B[18][26] +
                  mat_A[26][19] * mat_B[19][26] +
                  mat_A[26][20] * mat_B[20][26] +
                  mat_A[26][21] * mat_B[21][26] +
                  mat_A[26][22] * mat_B[22][26] +
                  mat_A[26][23] * mat_B[23][26] +
                  mat_A[26][24] * mat_B[24][26] +
                  mat_A[26][25] * mat_B[25][26] +
                  mat_A[26][26] * mat_B[26][26] +
                  mat_A[26][27] * mat_B[27][26] +
                  mat_A[26][28] * mat_B[28][26] +
                  mat_A[26][29] * mat_B[29][26] +
                  mat_A[26][30] * mat_B[30][26] +
                  mat_A[26][31] * mat_B[31][26];
    mat_C[26][27] <= 
                  mat_A[26][0] * mat_B[0][27] +
                  mat_A[26][1] * mat_B[1][27] +
                  mat_A[26][2] * mat_B[2][27] +
                  mat_A[26][3] * mat_B[3][27] +
                  mat_A[26][4] * mat_B[4][27] +
                  mat_A[26][5] * mat_B[5][27] +
                  mat_A[26][6] * mat_B[6][27] +
                  mat_A[26][7] * mat_B[7][27] +
                  mat_A[26][8] * mat_B[8][27] +
                  mat_A[26][9] * mat_B[9][27] +
                  mat_A[26][10] * mat_B[10][27] +
                  mat_A[26][11] * mat_B[11][27] +
                  mat_A[26][12] * mat_B[12][27] +
                  mat_A[26][13] * mat_B[13][27] +
                  mat_A[26][14] * mat_B[14][27] +
                  mat_A[26][15] * mat_B[15][27] +
                  mat_A[26][16] * mat_B[16][27] +
                  mat_A[26][17] * mat_B[17][27] +
                  mat_A[26][18] * mat_B[18][27] +
                  mat_A[26][19] * mat_B[19][27] +
                  mat_A[26][20] * mat_B[20][27] +
                  mat_A[26][21] * mat_B[21][27] +
                  mat_A[26][22] * mat_B[22][27] +
                  mat_A[26][23] * mat_B[23][27] +
                  mat_A[26][24] * mat_B[24][27] +
                  mat_A[26][25] * mat_B[25][27] +
                  mat_A[26][26] * mat_B[26][27] +
                  mat_A[26][27] * mat_B[27][27] +
                  mat_A[26][28] * mat_B[28][27] +
                  mat_A[26][29] * mat_B[29][27] +
                  mat_A[26][30] * mat_B[30][27] +
                  mat_A[26][31] * mat_B[31][27];
    mat_C[26][28] <= 
                  mat_A[26][0] * mat_B[0][28] +
                  mat_A[26][1] * mat_B[1][28] +
                  mat_A[26][2] * mat_B[2][28] +
                  mat_A[26][3] * mat_B[3][28] +
                  mat_A[26][4] * mat_B[4][28] +
                  mat_A[26][5] * mat_B[5][28] +
                  mat_A[26][6] * mat_B[6][28] +
                  mat_A[26][7] * mat_B[7][28] +
                  mat_A[26][8] * mat_B[8][28] +
                  mat_A[26][9] * mat_B[9][28] +
                  mat_A[26][10] * mat_B[10][28] +
                  mat_A[26][11] * mat_B[11][28] +
                  mat_A[26][12] * mat_B[12][28] +
                  mat_A[26][13] * mat_B[13][28] +
                  mat_A[26][14] * mat_B[14][28] +
                  mat_A[26][15] * mat_B[15][28] +
                  mat_A[26][16] * mat_B[16][28] +
                  mat_A[26][17] * mat_B[17][28] +
                  mat_A[26][18] * mat_B[18][28] +
                  mat_A[26][19] * mat_B[19][28] +
                  mat_A[26][20] * mat_B[20][28] +
                  mat_A[26][21] * mat_B[21][28] +
                  mat_A[26][22] * mat_B[22][28] +
                  mat_A[26][23] * mat_B[23][28] +
                  mat_A[26][24] * mat_B[24][28] +
                  mat_A[26][25] * mat_B[25][28] +
                  mat_A[26][26] * mat_B[26][28] +
                  mat_A[26][27] * mat_B[27][28] +
                  mat_A[26][28] * mat_B[28][28] +
                  mat_A[26][29] * mat_B[29][28] +
                  mat_A[26][30] * mat_B[30][28] +
                  mat_A[26][31] * mat_B[31][28];
    mat_C[26][29] <= 
                  mat_A[26][0] * mat_B[0][29] +
                  mat_A[26][1] * mat_B[1][29] +
                  mat_A[26][2] * mat_B[2][29] +
                  mat_A[26][3] * mat_B[3][29] +
                  mat_A[26][4] * mat_B[4][29] +
                  mat_A[26][5] * mat_B[5][29] +
                  mat_A[26][6] * mat_B[6][29] +
                  mat_A[26][7] * mat_B[7][29] +
                  mat_A[26][8] * mat_B[8][29] +
                  mat_A[26][9] * mat_B[9][29] +
                  mat_A[26][10] * mat_B[10][29] +
                  mat_A[26][11] * mat_B[11][29] +
                  mat_A[26][12] * mat_B[12][29] +
                  mat_A[26][13] * mat_B[13][29] +
                  mat_A[26][14] * mat_B[14][29] +
                  mat_A[26][15] * mat_B[15][29] +
                  mat_A[26][16] * mat_B[16][29] +
                  mat_A[26][17] * mat_B[17][29] +
                  mat_A[26][18] * mat_B[18][29] +
                  mat_A[26][19] * mat_B[19][29] +
                  mat_A[26][20] * mat_B[20][29] +
                  mat_A[26][21] * mat_B[21][29] +
                  mat_A[26][22] * mat_B[22][29] +
                  mat_A[26][23] * mat_B[23][29] +
                  mat_A[26][24] * mat_B[24][29] +
                  mat_A[26][25] * mat_B[25][29] +
                  mat_A[26][26] * mat_B[26][29] +
                  mat_A[26][27] * mat_B[27][29] +
                  mat_A[26][28] * mat_B[28][29] +
                  mat_A[26][29] * mat_B[29][29] +
                  mat_A[26][30] * mat_B[30][29] +
                  mat_A[26][31] * mat_B[31][29];
    mat_C[26][30] <= 
                  mat_A[26][0] * mat_B[0][30] +
                  mat_A[26][1] * mat_B[1][30] +
                  mat_A[26][2] * mat_B[2][30] +
                  mat_A[26][3] * mat_B[3][30] +
                  mat_A[26][4] * mat_B[4][30] +
                  mat_A[26][5] * mat_B[5][30] +
                  mat_A[26][6] * mat_B[6][30] +
                  mat_A[26][7] * mat_B[7][30] +
                  mat_A[26][8] * mat_B[8][30] +
                  mat_A[26][9] * mat_B[9][30] +
                  mat_A[26][10] * mat_B[10][30] +
                  mat_A[26][11] * mat_B[11][30] +
                  mat_A[26][12] * mat_B[12][30] +
                  mat_A[26][13] * mat_B[13][30] +
                  mat_A[26][14] * mat_B[14][30] +
                  mat_A[26][15] * mat_B[15][30] +
                  mat_A[26][16] * mat_B[16][30] +
                  mat_A[26][17] * mat_B[17][30] +
                  mat_A[26][18] * mat_B[18][30] +
                  mat_A[26][19] * mat_B[19][30] +
                  mat_A[26][20] * mat_B[20][30] +
                  mat_A[26][21] * mat_B[21][30] +
                  mat_A[26][22] * mat_B[22][30] +
                  mat_A[26][23] * mat_B[23][30] +
                  mat_A[26][24] * mat_B[24][30] +
                  mat_A[26][25] * mat_B[25][30] +
                  mat_A[26][26] * mat_B[26][30] +
                  mat_A[26][27] * mat_B[27][30] +
                  mat_A[26][28] * mat_B[28][30] +
                  mat_A[26][29] * mat_B[29][30] +
                  mat_A[26][30] * mat_B[30][30] +
                  mat_A[26][31] * mat_B[31][30];
    mat_C[26][31] <= 
                  mat_A[26][0] * mat_B[0][31] +
                  mat_A[26][1] * mat_B[1][31] +
                  mat_A[26][2] * mat_B[2][31] +
                  mat_A[26][3] * mat_B[3][31] +
                  mat_A[26][4] * mat_B[4][31] +
                  mat_A[26][5] * mat_B[5][31] +
                  mat_A[26][6] * mat_B[6][31] +
                  mat_A[26][7] * mat_B[7][31] +
                  mat_A[26][8] * mat_B[8][31] +
                  mat_A[26][9] * mat_B[9][31] +
                  mat_A[26][10] * mat_B[10][31] +
                  mat_A[26][11] * mat_B[11][31] +
                  mat_A[26][12] * mat_B[12][31] +
                  mat_A[26][13] * mat_B[13][31] +
                  mat_A[26][14] * mat_B[14][31] +
                  mat_A[26][15] * mat_B[15][31] +
                  mat_A[26][16] * mat_B[16][31] +
                  mat_A[26][17] * mat_B[17][31] +
                  mat_A[26][18] * mat_B[18][31] +
                  mat_A[26][19] * mat_B[19][31] +
                  mat_A[26][20] * mat_B[20][31] +
                  mat_A[26][21] * mat_B[21][31] +
                  mat_A[26][22] * mat_B[22][31] +
                  mat_A[26][23] * mat_B[23][31] +
                  mat_A[26][24] * mat_B[24][31] +
                  mat_A[26][25] * mat_B[25][31] +
                  mat_A[26][26] * mat_B[26][31] +
                  mat_A[26][27] * mat_B[27][31] +
                  mat_A[26][28] * mat_B[28][31] +
                  mat_A[26][29] * mat_B[29][31] +
                  mat_A[26][30] * mat_B[30][31] +
                  mat_A[26][31] * mat_B[31][31];
    mat_C[27][0] <= 
                  mat_A[27][0] * mat_B[0][0] +
                  mat_A[27][1] * mat_B[1][0] +
                  mat_A[27][2] * mat_B[2][0] +
                  mat_A[27][3] * mat_B[3][0] +
                  mat_A[27][4] * mat_B[4][0] +
                  mat_A[27][5] * mat_B[5][0] +
                  mat_A[27][6] * mat_B[6][0] +
                  mat_A[27][7] * mat_B[7][0] +
                  mat_A[27][8] * mat_B[8][0] +
                  mat_A[27][9] * mat_B[9][0] +
                  mat_A[27][10] * mat_B[10][0] +
                  mat_A[27][11] * mat_B[11][0] +
                  mat_A[27][12] * mat_B[12][0] +
                  mat_A[27][13] * mat_B[13][0] +
                  mat_A[27][14] * mat_B[14][0] +
                  mat_A[27][15] * mat_B[15][0] +
                  mat_A[27][16] * mat_B[16][0] +
                  mat_A[27][17] * mat_B[17][0] +
                  mat_A[27][18] * mat_B[18][0] +
                  mat_A[27][19] * mat_B[19][0] +
                  mat_A[27][20] * mat_B[20][0] +
                  mat_A[27][21] * mat_B[21][0] +
                  mat_A[27][22] * mat_B[22][0] +
                  mat_A[27][23] * mat_B[23][0] +
                  mat_A[27][24] * mat_B[24][0] +
                  mat_A[27][25] * mat_B[25][0] +
                  mat_A[27][26] * mat_B[26][0] +
                  mat_A[27][27] * mat_B[27][0] +
                  mat_A[27][28] * mat_B[28][0] +
                  mat_A[27][29] * mat_B[29][0] +
                  mat_A[27][30] * mat_B[30][0] +
                  mat_A[27][31] * mat_B[31][0];
    mat_C[27][1] <= 
                  mat_A[27][0] * mat_B[0][1] +
                  mat_A[27][1] * mat_B[1][1] +
                  mat_A[27][2] * mat_B[2][1] +
                  mat_A[27][3] * mat_B[3][1] +
                  mat_A[27][4] * mat_B[4][1] +
                  mat_A[27][5] * mat_B[5][1] +
                  mat_A[27][6] * mat_B[6][1] +
                  mat_A[27][7] * mat_B[7][1] +
                  mat_A[27][8] * mat_B[8][1] +
                  mat_A[27][9] * mat_B[9][1] +
                  mat_A[27][10] * mat_B[10][1] +
                  mat_A[27][11] * mat_B[11][1] +
                  mat_A[27][12] * mat_B[12][1] +
                  mat_A[27][13] * mat_B[13][1] +
                  mat_A[27][14] * mat_B[14][1] +
                  mat_A[27][15] * mat_B[15][1] +
                  mat_A[27][16] * mat_B[16][1] +
                  mat_A[27][17] * mat_B[17][1] +
                  mat_A[27][18] * mat_B[18][1] +
                  mat_A[27][19] * mat_B[19][1] +
                  mat_A[27][20] * mat_B[20][1] +
                  mat_A[27][21] * mat_B[21][1] +
                  mat_A[27][22] * mat_B[22][1] +
                  mat_A[27][23] * mat_B[23][1] +
                  mat_A[27][24] * mat_B[24][1] +
                  mat_A[27][25] * mat_B[25][1] +
                  mat_A[27][26] * mat_B[26][1] +
                  mat_A[27][27] * mat_B[27][1] +
                  mat_A[27][28] * mat_B[28][1] +
                  mat_A[27][29] * mat_B[29][1] +
                  mat_A[27][30] * mat_B[30][1] +
                  mat_A[27][31] * mat_B[31][1];
    mat_C[27][2] <= 
                  mat_A[27][0] * mat_B[0][2] +
                  mat_A[27][1] * mat_B[1][2] +
                  mat_A[27][2] * mat_B[2][2] +
                  mat_A[27][3] * mat_B[3][2] +
                  mat_A[27][4] * mat_B[4][2] +
                  mat_A[27][5] * mat_B[5][2] +
                  mat_A[27][6] * mat_B[6][2] +
                  mat_A[27][7] * mat_B[7][2] +
                  mat_A[27][8] * mat_B[8][2] +
                  mat_A[27][9] * mat_B[9][2] +
                  mat_A[27][10] * mat_B[10][2] +
                  mat_A[27][11] * mat_B[11][2] +
                  mat_A[27][12] * mat_B[12][2] +
                  mat_A[27][13] * mat_B[13][2] +
                  mat_A[27][14] * mat_B[14][2] +
                  mat_A[27][15] * mat_B[15][2] +
                  mat_A[27][16] * mat_B[16][2] +
                  mat_A[27][17] * mat_B[17][2] +
                  mat_A[27][18] * mat_B[18][2] +
                  mat_A[27][19] * mat_B[19][2] +
                  mat_A[27][20] * mat_B[20][2] +
                  mat_A[27][21] * mat_B[21][2] +
                  mat_A[27][22] * mat_B[22][2] +
                  mat_A[27][23] * mat_B[23][2] +
                  mat_A[27][24] * mat_B[24][2] +
                  mat_A[27][25] * mat_B[25][2] +
                  mat_A[27][26] * mat_B[26][2] +
                  mat_A[27][27] * mat_B[27][2] +
                  mat_A[27][28] * mat_B[28][2] +
                  mat_A[27][29] * mat_B[29][2] +
                  mat_A[27][30] * mat_B[30][2] +
                  mat_A[27][31] * mat_B[31][2];
    mat_C[27][3] <= 
                  mat_A[27][0] * mat_B[0][3] +
                  mat_A[27][1] * mat_B[1][3] +
                  mat_A[27][2] * mat_B[2][3] +
                  mat_A[27][3] * mat_B[3][3] +
                  mat_A[27][4] * mat_B[4][3] +
                  mat_A[27][5] * mat_B[5][3] +
                  mat_A[27][6] * mat_B[6][3] +
                  mat_A[27][7] * mat_B[7][3] +
                  mat_A[27][8] * mat_B[8][3] +
                  mat_A[27][9] * mat_B[9][3] +
                  mat_A[27][10] * mat_B[10][3] +
                  mat_A[27][11] * mat_B[11][3] +
                  mat_A[27][12] * mat_B[12][3] +
                  mat_A[27][13] * mat_B[13][3] +
                  mat_A[27][14] * mat_B[14][3] +
                  mat_A[27][15] * mat_B[15][3] +
                  mat_A[27][16] * mat_B[16][3] +
                  mat_A[27][17] * mat_B[17][3] +
                  mat_A[27][18] * mat_B[18][3] +
                  mat_A[27][19] * mat_B[19][3] +
                  mat_A[27][20] * mat_B[20][3] +
                  mat_A[27][21] * mat_B[21][3] +
                  mat_A[27][22] * mat_B[22][3] +
                  mat_A[27][23] * mat_B[23][3] +
                  mat_A[27][24] * mat_B[24][3] +
                  mat_A[27][25] * mat_B[25][3] +
                  mat_A[27][26] * mat_B[26][3] +
                  mat_A[27][27] * mat_B[27][3] +
                  mat_A[27][28] * mat_B[28][3] +
                  mat_A[27][29] * mat_B[29][3] +
                  mat_A[27][30] * mat_B[30][3] +
                  mat_A[27][31] * mat_B[31][3];
    mat_C[27][4] <= 
                  mat_A[27][0] * mat_B[0][4] +
                  mat_A[27][1] * mat_B[1][4] +
                  mat_A[27][2] * mat_B[2][4] +
                  mat_A[27][3] * mat_B[3][4] +
                  mat_A[27][4] * mat_B[4][4] +
                  mat_A[27][5] * mat_B[5][4] +
                  mat_A[27][6] * mat_B[6][4] +
                  mat_A[27][7] * mat_B[7][4] +
                  mat_A[27][8] * mat_B[8][4] +
                  mat_A[27][9] * mat_B[9][4] +
                  mat_A[27][10] * mat_B[10][4] +
                  mat_A[27][11] * mat_B[11][4] +
                  mat_A[27][12] * mat_B[12][4] +
                  mat_A[27][13] * mat_B[13][4] +
                  mat_A[27][14] * mat_B[14][4] +
                  mat_A[27][15] * mat_B[15][4] +
                  mat_A[27][16] * mat_B[16][4] +
                  mat_A[27][17] * mat_B[17][4] +
                  mat_A[27][18] * mat_B[18][4] +
                  mat_A[27][19] * mat_B[19][4] +
                  mat_A[27][20] * mat_B[20][4] +
                  mat_A[27][21] * mat_B[21][4] +
                  mat_A[27][22] * mat_B[22][4] +
                  mat_A[27][23] * mat_B[23][4] +
                  mat_A[27][24] * mat_B[24][4] +
                  mat_A[27][25] * mat_B[25][4] +
                  mat_A[27][26] * mat_B[26][4] +
                  mat_A[27][27] * mat_B[27][4] +
                  mat_A[27][28] * mat_B[28][4] +
                  mat_A[27][29] * mat_B[29][4] +
                  mat_A[27][30] * mat_B[30][4] +
                  mat_A[27][31] * mat_B[31][4];
    mat_C[27][5] <= 
                  mat_A[27][0] * mat_B[0][5] +
                  mat_A[27][1] * mat_B[1][5] +
                  mat_A[27][2] * mat_B[2][5] +
                  mat_A[27][3] * mat_B[3][5] +
                  mat_A[27][4] * mat_B[4][5] +
                  mat_A[27][5] * mat_B[5][5] +
                  mat_A[27][6] * mat_B[6][5] +
                  mat_A[27][7] * mat_B[7][5] +
                  mat_A[27][8] * mat_B[8][5] +
                  mat_A[27][9] * mat_B[9][5] +
                  mat_A[27][10] * mat_B[10][5] +
                  mat_A[27][11] * mat_B[11][5] +
                  mat_A[27][12] * mat_B[12][5] +
                  mat_A[27][13] * mat_B[13][5] +
                  mat_A[27][14] * mat_B[14][5] +
                  mat_A[27][15] * mat_B[15][5] +
                  mat_A[27][16] * mat_B[16][5] +
                  mat_A[27][17] * mat_B[17][5] +
                  mat_A[27][18] * mat_B[18][5] +
                  mat_A[27][19] * mat_B[19][5] +
                  mat_A[27][20] * mat_B[20][5] +
                  mat_A[27][21] * mat_B[21][5] +
                  mat_A[27][22] * mat_B[22][5] +
                  mat_A[27][23] * mat_B[23][5] +
                  mat_A[27][24] * mat_B[24][5] +
                  mat_A[27][25] * mat_B[25][5] +
                  mat_A[27][26] * mat_B[26][5] +
                  mat_A[27][27] * mat_B[27][5] +
                  mat_A[27][28] * mat_B[28][5] +
                  mat_A[27][29] * mat_B[29][5] +
                  mat_A[27][30] * mat_B[30][5] +
                  mat_A[27][31] * mat_B[31][5];
    mat_C[27][6] <= 
                  mat_A[27][0] * mat_B[0][6] +
                  mat_A[27][1] * mat_B[1][6] +
                  mat_A[27][2] * mat_B[2][6] +
                  mat_A[27][3] * mat_B[3][6] +
                  mat_A[27][4] * mat_B[4][6] +
                  mat_A[27][5] * mat_B[5][6] +
                  mat_A[27][6] * mat_B[6][6] +
                  mat_A[27][7] * mat_B[7][6] +
                  mat_A[27][8] * mat_B[8][6] +
                  mat_A[27][9] * mat_B[9][6] +
                  mat_A[27][10] * mat_B[10][6] +
                  mat_A[27][11] * mat_B[11][6] +
                  mat_A[27][12] * mat_B[12][6] +
                  mat_A[27][13] * mat_B[13][6] +
                  mat_A[27][14] * mat_B[14][6] +
                  mat_A[27][15] * mat_B[15][6] +
                  mat_A[27][16] * mat_B[16][6] +
                  mat_A[27][17] * mat_B[17][6] +
                  mat_A[27][18] * mat_B[18][6] +
                  mat_A[27][19] * mat_B[19][6] +
                  mat_A[27][20] * mat_B[20][6] +
                  mat_A[27][21] * mat_B[21][6] +
                  mat_A[27][22] * mat_B[22][6] +
                  mat_A[27][23] * mat_B[23][6] +
                  mat_A[27][24] * mat_B[24][6] +
                  mat_A[27][25] * mat_B[25][6] +
                  mat_A[27][26] * mat_B[26][6] +
                  mat_A[27][27] * mat_B[27][6] +
                  mat_A[27][28] * mat_B[28][6] +
                  mat_A[27][29] * mat_B[29][6] +
                  mat_A[27][30] * mat_B[30][6] +
                  mat_A[27][31] * mat_B[31][6];
    mat_C[27][7] <= 
                  mat_A[27][0] * mat_B[0][7] +
                  mat_A[27][1] * mat_B[1][7] +
                  mat_A[27][2] * mat_B[2][7] +
                  mat_A[27][3] * mat_B[3][7] +
                  mat_A[27][4] * mat_B[4][7] +
                  mat_A[27][5] * mat_B[5][7] +
                  mat_A[27][6] * mat_B[6][7] +
                  mat_A[27][7] * mat_B[7][7] +
                  mat_A[27][8] * mat_B[8][7] +
                  mat_A[27][9] * mat_B[9][7] +
                  mat_A[27][10] * mat_B[10][7] +
                  mat_A[27][11] * mat_B[11][7] +
                  mat_A[27][12] * mat_B[12][7] +
                  mat_A[27][13] * mat_B[13][7] +
                  mat_A[27][14] * mat_B[14][7] +
                  mat_A[27][15] * mat_B[15][7] +
                  mat_A[27][16] * mat_B[16][7] +
                  mat_A[27][17] * mat_B[17][7] +
                  mat_A[27][18] * mat_B[18][7] +
                  mat_A[27][19] * mat_B[19][7] +
                  mat_A[27][20] * mat_B[20][7] +
                  mat_A[27][21] * mat_B[21][7] +
                  mat_A[27][22] * mat_B[22][7] +
                  mat_A[27][23] * mat_B[23][7] +
                  mat_A[27][24] * mat_B[24][7] +
                  mat_A[27][25] * mat_B[25][7] +
                  mat_A[27][26] * mat_B[26][7] +
                  mat_A[27][27] * mat_B[27][7] +
                  mat_A[27][28] * mat_B[28][7] +
                  mat_A[27][29] * mat_B[29][7] +
                  mat_A[27][30] * mat_B[30][7] +
                  mat_A[27][31] * mat_B[31][7];
    mat_C[27][8] <= 
                  mat_A[27][0] * mat_B[0][8] +
                  mat_A[27][1] * mat_B[1][8] +
                  mat_A[27][2] * mat_B[2][8] +
                  mat_A[27][3] * mat_B[3][8] +
                  mat_A[27][4] * mat_B[4][8] +
                  mat_A[27][5] * mat_B[5][8] +
                  mat_A[27][6] * mat_B[6][8] +
                  mat_A[27][7] * mat_B[7][8] +
                  mat_A[27][8] * mat_B[8][8] +
                  mat_A[27][9] * mat_B[9][8] +
                  mat_A[27][10] * mat_B[10][8] +
                  mat_A[27][11] * mat_B[11][8] +
                  mat_A[27][12] * mat_B[12][8] +
                  mat_A[27][13] * mat_B[13][8] +
                  mat_A[27][14] * mat_B[14][8] +
                  mat_A[27][15] * mat_B[15][8] +
                  mat_A[27][16] * mat_B[16][8] +
                  mat_A[27][17] * mat_B[17][8] +
                  mat_A[27][18] * mat_B[18][8] +
                  mat_A[27][19] * mat_B[19][8] +
                  mat_A[27][20] * mat_B[20][8] +
                  mat_A[27][21] * mat_B[21][8] +
                  mat_A[27][22] * mat_B[22][8] +
                  mat_A[27][23] * mat_B[23][8] +
                  mat_A[27][24] * mat_B[24][8] +
                  mat_A[27][25] * mat_B[25][8] +
                  mat_A[27][26] * mat_B[26][8] +
                  mat_A[27][27] * mat_B[27][8] +
                  mat_A[27][28] * mat_B[28][8] +
                  mat_A[27][29] * mat_B[29][8] +
                  mat_A[27][30] * mat_B[30][8] +
                  mat_A[27][31] * mat_B[31][8];
    mat_C[27][9] <= 
                  mat_A[27][0] * mat_B[0][9] +
                  mat_A[27][1] * mat_B[1][9] +
                  mat_A[27][2] * mat_B[2][9] +
                  mat_A[27][3] * mat_B[3][9] +
                  mat_A[27][4] * mat_B[4][9] +
                  mat_A[27][5] * mat_B[5][9] +
                  mat_A[27][6] * mat_B[6][9] +
                  mat_A[27][7] * mat_B[7][9] +
                  mat_A[27][8] * mat_B[8][9] +
                  mat_A[27][9] * mat_B[9][9] +
                  mat_A[27][10] * mat_B[10][9] +
                  mat_A[27][11] * mat_B[11][9] +
                  mat_A[27][12] * mat_B[12][9] +
                  mat_A[27][13] * mat_B[13][9] +
                  mat_A[27][14] * mat_B[14][9] +
                  mat_A[27][15] * mat_B[15][9] +
                  mat_A[27][16] * mat_B[16][9] +
                  mat_A[27][17] * mat_B[17][9] +
                  mat_A[27][18] * mat_B[18][9] +
                  mat_A[27][19] * mat_B[19][9] +
                  mat_A[27][20] * mat_B[20][9] +
                  mat_A[27][21] * mat_B[21][9] +
                  mat_A[27][22] * mat_B[22][9] +
                  mat_A[27][23] * mat_B[23][9] +
                  mat_A[27][24] * mat_B[24][9] +
                  mat_A[27][25] * mat_B[25][9] +
                  mat_A[27][26] * mat_B[26][9] +
                  mat_A[27][27] * mat_B[27][9] +
                  mat_A[27][28] * mat_B[28][9] +
                  mat_A[27][29] * mat_B[29][9] +
                  mat_A[27][30] * mat_B[30][9] +
                  mat_A[27][31] * mat_B[31][9];
    mat_C[27][10] <= 
                  mat_A[27][0] * mat_B[0][10] +
                  mat_A[27][1] * mat_B[1][10] +
                  mat_A[27][2] * mat_B[2][10] +
                  mat_A[27][3] * mat_B[3][10] +
                  mat_A[27][4] * mat_B[4][10] +
                  mat_A[27][5] * mat_B[5][10] +
                  mat_A[27][6] * mat_B[6][10] +
                  mat_A[27][7] * mat_B[7][10] +
                  mat_A[27][8] * mat_B[8][10] +
                  mat_A[27][9] * mat_B[9][10] +
                  mat_A[27][10] * mat_B[10][10] +
                  mat_A[27][11] * mat_B[11][10] +
                  mat_A[27][12] * mat_B[12][10] +
                  mat_A[27][13] * mat_B[13][10] +
                  mat_A[27][14] * mat_B[14][10] +
                  mat_A[27][15] * mat_B[15][10] +
                  mat_A[27][16] * mat_B[16][10] +
                  mat_A[27][17] * mat_B[17][10] +
                  mat_A[27][18] * mat_B[18][10] +
                  mat_A[27][19] * mat_B[19][10] +
                  mat_A[27][20] * mat_B[20][10] +
                  mat_A[27][21] * mat_B[21][10] +
                  mat_A[27][22] * mat_B[22][10] +
                  mat_A[27][23] * mat_B[23][10] +
                  mat_A[27][24] * mat_B[24][10] +
                  mat_A[27][25] * mat_B[25][10] +
                  mat_A[27][26] * mat_B[26][10] +
                  mat_A[27][27] * mat_B[27][10] +
                  mat_A[27][28] * mat_B[28][10] +
                  mat_A[27][29] * mat_B[29][10] +
                  mat_A[27][30] * mat_B[30][10] +
                  mat_A[27][31] * mat_B[31][10];
    mat_C[27][11] <= 
                  mat_A[27][0] * mat_B[0][11] +
                  mat_A[27][1] * mat_B[1][11] +
                  mat_A[27][2] * mat_B[2][11] +
                  mat_A[27][3] * mat_B[3][11] +
                  mat_A[27][4] * mat_B[4][11] +
                  mat_A[27][5] * mat_B[5][11] +
                  mat_A[27][6] * mat_B[6][11] +
                  mat_A[27][7] * mat_B[7][11] +
                  mat_A[27][8] * mat_B[8][11] +
                  mat_A[27][9] * mat_B[9][11] +
                  mat_A[27][10] * mat_B[10][11] +
                  mat_A[27][11] * mat_B[11][11] +
                  mat_A[27][12] * mat_B[12][11] +
                  mat_A[27][13] * mat_B[13][11] +
                  mat_A[27][14] * mat_B[14][11] +
                  mat_A[27][15] * mat_B[15][11] +
                  mat_A[27][16] * mat_B[16][11] +
                  mat_A[27][17] * mat_B[17][11] +
                  mat_A[27][18] * mat_B[18][11] +
                  mat_A[27][19] * mat_B[19][11] +
                  mat_A[27][20] * mat_B[20][11] +
                  mat_A[27][21] * mat_B[21][11] +
                  mat_A[27][22] * mat_B[22][11] +
                  mat_A[27][23] * mat_B[23][11] +
                  mat_A[27][24] * mat_B[24][11] +
                  mat_A[27][25] * mat_B[25][11] +
                  mat_A[27][26] * mat_B[26][11] +
                  mat_A[27][27] * mat_B[27][11] +
                  mat_A[27][28] * mat_B[28][11] +
                  mat_A[27][29] * mat_B[29][11] +
                  mat_A[27][30] * mat_B[30][11] +
                  mat_A[27][31] * mat_B[31][11];
    mat_C[27][12] <= 
                  mat_A[27][0] * mat_B[0][12] +
                  mat_A[27][1] * mat_B[1][12] +
                  mat_A[27][2] * mat_B[2][12] +
                  mat_A[27][3] * mat_B[3][12] +
                  mat_A[27][4] * mat_B[4][12] +
                  mat_A[27][5] * mat_B[5][12] +
                  mat_A[27][6] * mat_B[6][12] +
                  mat_A[27][7] * mat_B[7][12] +
                  mat_A[27][8] * mat_B[8][12] +
                  mat_A[27][9] * mat_B[9][12] +
                  mat_A[27][10] * mat_B[10][12] +
                  mat_A[27][11] * mat_B[11][12] +
                  mat_A[27][12] * mat_B[12][12] +
                  mat_A[27][13] * mat_B[13][12] +
                  mat_A[27][14] * mat_B[14][12] +
                  mat_A[27][15] * mat_B[15][12] +
                  mat_A[27][16] * mat_B[16][12] +
                  mat_A[27][17] * mat_B[17][12] +
                  mat_A[27][18] * mat_B[18][12] +
                  mat_A[27][19] * mat_B[19][12] +
                  mat_A[27][20] * mat_B[20][12] +
                  mat_A[27][21] * mat_B[21][12] +
                  mat_A[27][22] * mat_B[22][12] +
                  mat_A[27][23] * mat_B[23][12] +
                  mat_A[27][24] * mat_B[24][12] +
                  mat_A[27][25] * mat_B[25][12] +
                  mat_A[27][26] * mat_B[26][12] +
                  mat_A[27][27] * mat_B[27][12] +
                  mat_A[27][28] * mat_B[28][12] +
                  mat_A[27][29] * mat_B[29][12] +
                  mat_A[27][30] * mat_B[30][12] +
                  mat_A[27][31] * mat_B[31][12];
    mat_C[27][13] <= 
                  mat_A[27][0] * mat_B[0][13] +
                  mat_A[27][1] * mat_B[1][13] +
                  mat_A[27][2] * mat_B[2][13] +
                  mat_A[27][3] * mat_B[3][13] +
                  mat_A[27][4] * mat_B[4][13] +
                  mat_A[27][5] * mat_B[5][13] +
                  mat_A[27][6] * mat_B[6][13] +
                  mat_A[27][7] * mat_B[7][13] +
                  mat_A[27][8] * mat_B[8][13] +
                  mat_A[27][9] * mat_B[9][13] +
                  mat_A[27][10] * mat_B[10][13] +
                  mat_A[27][11] * mat_B[11][13] +
                  mat_A[27][12] * mat_B[12][13] +
                  mat_A[27][13] * mat_B[13][13] +
                  mat_A[27][14] * mat_B[14][13] +
                  mat_A[27][15] * mat_B[15][13] +
                  mat_A[27][16] * mat_B[16][13] +
                  mat_A[27][17] * mat_B[17][13] +
                  mat_A[27][18] * mat_B[18][13] +
                  mat_A[27][19] * mat_B[19][13] +
                  mat_A[27][20] * mat_B[20][13] +
                  mat_A[27][21] * mat_B[21][13] +
                  mat_A[27][22] * mat_B[22][13] +
                  mat_A[27][23] * mat_B[23][13] +
                  mat_A[27][24] * mat_B[24][13] +
                  mat_A[27][25] * mat_B[25][13] +
                  mat_A[27][26] * mat_B[26][13] +
                  mat_A[27][27] * mat_B[27][13] +
                  mat_A[27][28] * mat_B[28][13] +
                  mat_A[27][29] * mat_B[29][13] +
                  mat_A[27][30] * mat_B[30][13] +
                  mat_A[27][31] * mat_B[31][13];
    mat_C[27][14] <= 
                  mat_A[27][0] * mat_B[0][14] +
                  mat_A[27][1] * mat_B[1][14] +
                  mat_A[27][2] * mat_B[2][14] +
                  mat_A[27][3] * mat_B[3][14] +
                  mat_A[27][4] * mat_B[4][14] +
                  mat_A[27][5] * mat_B[5][14] +
                  mat_A[27][6] * mat_B[6][14] +
                  mat_A[27][7] * mat_B[7][14] +
                  mat_A[27][8] * mat_B[8][14] +
                  mat_A[27][9] * mat_B[9][14] +
                  mat_A[27][10] * mat_B[10][14] +
                  mat_A[27][11] * mat_B[11][14] +
                  mat_A[27][12] * mat_B[12][14] +
                  mat_A[27][13] * mat_B[13][14] +
                  mat_A[27][14] * mat_B[14][14] +
                  mat_A[27][15] * mat_B[15][14] +
                  mat_A[27][16] * mat_B[16][14] +
                  mat_A[27][17] * mat_B[17][14] +
                  mat_A[27][18] * mat_B[18][14] +
                  mat_A[27][19] * mat_B[19][14] +
                  mat_A[27][20] * mat_B[20][14] +
                  mat_A[27][21] * mat_B[21][14] +
                  mat_A[27][22] * mat_B[22][14] +
                  mat_A[27][23] * mat_B[23][14] +
                  mat_A[27][24] * mat_B[24][14] +
                  mat_A[27][25] * mat_B[25][14] +
                  mat_A[27][26] * mat_B[26][14] +
                  mat_A[27][27] * mat_B[27][14] +
                  mat_A[27][28] * mat_B[28][14] +
                  mat_A[27][29] * mat_B[29][14] +
                  mat_A[27][30] * mat_B[30][14] +
                  mat_A[27][31] * mat_B[31][14];
    mat_C[27][15] <= 
                  mat_A[27][0] * mat_B[0][15] +
                  mat_A[27][1] * mat_B[1][15] +
                  mat_A[27][2] * mat_B[2][15] +
                  mat_A[27][3] * mat_B[3][15] +
                  mat_A[27][4] * mat_B[4][15] +
                  mat_A[27][5] * mat_B[5][15] +
                  mat_A[27][6] * mat_B[6][15] +
                  mat_A[27][7] * mat_B[7][15] +
                  mat_A[27][8] * mat_B[8][15] +
                  mat_A[27][9] * mat_B[9][15] +
                  mat_A[27][10] * mat_B[10][15] +
                  mat_A[27][11] * mat_B[11][15] +
                  mat_A[27][12] * mat_B[12][15] +
                  mat_A[27][13] * mat_B[13][15] +
                  mat_A[27][14] * mat_B[14][15] +
                  mat_A[27][15] * mat_B[15][15] +
                  mat_A[27][16] * mat_B[16][15] +
                  mat_A[27][17] * mat_B[17][15] +
                  mat_A[27][18] * mat_B[18][15] +
                  mat_A[27][19] * mat_B[19][15] +
                  mat_A[27][20] * mat_B[20][15] +
                  mat_A[27][21] * mat_B[21][15] +
                  mat_A[27][22] * mat_B[22][15] +
                  mat_A[27][23] * mat_B[23][15] +
                  mat_A[27][24] * mat_B[24][15] +
                  mat_A[27][25] * mat_B[25][15] +
                  mat_A[27][26] * mat_B[26][15] +
                  mat_A[27][27] * mat_B[27][15] +
                  mat_A[27][28] * mat_B[28][15] +
                  mat_A[27][29] * mat_B[29][15] +
                  mat_A[27][30] * mat_B[30][15] +
                  mat_A[27][31] * mat_B[31][15];
    mat_C[27][16] <= 
                  mat_A[27][0] * mat_B[0][16] +
                  mat_A[27][1] * mat_B[1][16] +
                  mat_A[27][2] * mat_B[2][16] +
                  mat_A[27][3] * mat_B[3][16] +
                  mat_A[27][4] * mat_B[4][16] +
                  mat_A[27][5] * mat_B[5][16] +
                  mat_A[27][6] * mat_B[6][16] +
                  mat_A[27][7] * mat_B[7][16] +
                  mat_A[27][8] * mat_B[8][16] +
                  mat_A[27][9] * mat_B[9][16] +
                  mat_A[27][10] * mat_B[10][16] +
                  mat_A[27][11] * mat_B[11][16] +
                  mat_A[27][12] * mat_B[12][16] +
                  mat_A[27][13] * mat_B[13][16] +
                  mat_A[27][14] * mat_B[14][16] +
                  mat_A[27][15] * mat_B[15][16] +
                  mat_A[27][16] * mat_B[16][16] +
                  mat_A[27][17] * mat_B[17][16] +
                  mat_A[27][18] * mat_B[18][16] +
                  mat_A[27][19] * mat_B[19][16] +
                  mat_A[27][20] * mat_B[20][16] +
                  mat_A[27][21] * mat_B[21][16] +
                  mat_A[27][22] * mat_B[22][16] +
                  mat_A[27][23] * mat_B[23][16] +
                  mat_A[27][24] * mat_B[24][16] +
                  mat_A[27][25] * mat_B[25][16] +
                  mat_A[27][26] * mat_B[26][16] +
                  mat_A[27][27] * mat_B[27][16] +
                  mat_A[27][28] * mat_B[28][16] +
                  mat_A[27][29] * mat_B[29][16] +
                  mat_A[27][30] * mat_B[30][16] +
                  mat_A[27][31] * mat_B[31][16];
    mat_C[27][17] <= 
                  mat_A[27][0] * mat_B[0][17] +
                  mat_A[27][1] * mat_B[1][17] +
                  mat_A[27][2] * mat_B[2][17] +
                  mat_A[27][3] * mat_B[3][17] +
                  mat_A[27][4] * mat_B[4][17] +
                  mat_A[27][5] * mat_B[5][17] +
                  mat_A[27][6] * mat_B[6][17] +
                  mat_A[27][7] * mat_B[7][17] +
                  mat_A[27][8] * mat_B[8][17] +
                  mat_A[27][9] * mat_B[9][17] +
                  mat_A[27][10] * mat_B[10][17] +
                  mat_A[27][11] * mat_B[11][17] +
                  mat_A[27][12] * mat_B[12][17] +
                  mat_A[27][13] * mat_B[13][17] +
                  mat_A[27][14] * mat_B[14][17] +
                  mat_A[27][15] * mat_B[15][17] +
                  mat_A[27][16] * mat_B[16][17] +
                  mat_A[27][17] * mat_B[17][17] +
                  mat_A[27][18] * mat_B[18][17] +
                  mat_A[27][19] * mat_B[19][17] +
                  mat_A[27][20] * mat_B[20][17] +
                  mat_A[27][21] * mat_B[21][17] +
                  mat_A[27][22] * mat_B[22][17] +
                  mat_A[27][23] * mat_B[23][17] +
                  mat_A[27][24] * mat_B[24][17] +
                  mat_A[27][25] * mat_B[25][17] +
                  mat_A[27][26] * mat_B[26][17] +
                  mat_A[27][27] * mat_B[27][17] +
                  mat_A[27][28] * mat_B[28][17] +
                  mat_A[27][29] * mat_B[29][17] +
                  mat_A[27][30] * mat_B[30][17] +
                  mat_A[27][31] * mat_B[31][17];
    mat_C[27][18] <= 
                  mat_A[27][0] * mat_B[0][18] +
                  mat_A[27][1] * mat_B[1][18] +
                  mat_A[27][2] * mat_B[2][18] +
                  mat_A[27][3] * mat_B[3][18] +
                  mat_A[27][4] * mat_B[4][18] +
                  mat_A[27][5] * mat_B[5][18] +
                  mat_A[27][6] * mat_B[6][18] +
                  mat_A[27][7] * mat_B[7][18] +
                  mat_A[27][8] * mat_B[8][18] +
                  mat_A[27][9] * mat_B[9][18] +
                  mat_A[27][10] * mat_B[10][18] +
                  mat_A[27][11] * mat_B[11][18] +
                  mat_A[27][12] * mat_B[12][18] +
                  mat_A[27][13] * mat_B[13][18] +
                  mat_A[27][14] * mat_B[14][18] +
                  mat_A[27][15] * mat_B[15][18] +
                  mat_A[27][16] * mat_B[16][18] +
                  mat_A[27][17] * mat_B[17][18] +
                  mat_A[27][18] * mat_B[18][18] +
                  mat_A[27][19] * mat_B[19][18] +
                  mat_A[27][20] * mat_B[20][18] +
                  mat_A[27][21] * mat_B[21][18] +
                  mat_A[27][22] * mat_B[22][18] +
                  mat_A[27][23] * mat_B[23][18] +
                  mat_A[27][24] * mat_B[24][18] +
                  mat_A[27][25] * mat_B[25][18] +
                  mat_A[27][26] * mat_B[26][18] +
                  mat_A[27][27] * mat_B[27][18] +
                  mat_A[27][28] * mat_B[28][18] +
                  mat_A[27][29] * mat_B[29][18] +
                  mat_A[27][30] * mat_B[30][18] +
                  mat_A[27][31] * mat_B[31][18];
    mat_C[27][19] <= 
                  mat_A[27][0] * mat_B[0][19] +
                  mat_A[27][1] * mat_B[1][19] +
                  mat_A[27][2] * mat_B[2][19] +
                  mat_A[27][3] * mat_B[3][19] +
                  mat_A[27][4] * mat_B[4][19] +
                  mat_A[27][5] * mat_B[5][19] +
                  mat_A[27][6] * mat_B[6][19] +
                  mat_A[27][7] * mat_B[7][19] +
                  mat_A[27][8] * mat_B[8][19] +
                  mat_A[27][9] * mat_B[9][19] +
                  mat_A[27][10] * mat_B[10][19] +
                  mat_A[27][11] * mat_B[11][19] +
                  mat_A[27][12] * mat_B[12][19] +
                  mat_A[27][13] * mat_B[13][19] +
                  mat_A[27][14] * mat_B[14][19] +
                  mat_A[27][15] * mat_B[15][19] +
                  mat_A[27][16] * mat_B[16][19] +
                  mat_A[27][17] * mat_B[17][19] +
                  mat_A[27][18] * mat_B[18][19] +
                  mat_A[27][19] * mat_B[19][19] +
                  mat_A[27][20] * mat_B[20][19] +
                  mat_A[27][21] * mat_B[21][19] +
                  mat_A[27][22] * mat_B[22][19] +
                  mat_A[27][23] * mat_B[23][19] +
                  mat_A[27][24] * mat_B[24][19] +
                  mat_A[27][25] * mat_B[25][19] +
                  mat_A[27][26] * mat_B[26][19] +
                  mat_A[27][27] * mat_B[27][19] +
                  mat_A[27][28] * mat_B[28][19] +
                  mat_A[27][29] * mat_B[29][19] +
                  mat_A[27][30] * mat_B[30][19] +
                  mat_A[27][31] * mat_B[31][19];
    mat_C[27][20] <= 
                  mat_A[27][0] * mat_B[0][20] +
                  mat_A[27][1] * mat_B[1][20] +
                  mat_A[27][2] * mat_B[2][20] +
                  mat_A[27][3] * mat_B[3][20] +
                  mat_A[27][4] * mat_B[4][20] +
                  mat_A[27][5] * mat_B[5][20] +
                  mat_A[27][6] * mat_B[6][20] +
                  mat_A[27][7] * mat_B[7][20] +
                  mat_A[27][8] * mat_B[8][20] +
                  mat_A[27][9] * mat_B[9][20] +
                  mat_A[27][10] * mat_B[10][20] +
                  mat_A[27][11] * mat_B[11][20] +
                  mat_A[27][12] * mat_B[12][20] +
                  mat_A[27][13] * mat_B[13][20] +
                  mat_A[27][14] * mat_B[14][20] +
                  mat_A[27][15] * mat_B[15][20] +
                  mat_A[27][16] * mat_B[16][20] +
                  mat_A[27][17] * mat_B[17][20] +
                  mat_A[27][18] * mat_B[18][20] +
                  mat_A[27][19] * mat_B[19][20] +
                  mat_A[27][20] * mat_B[20][20] +
                  mat_A[27][21] * mat_B[21][20] +
                  mat_A[27][22] * mat_B[22][20] +
                  mat_A[27][23] * mat_B[23][20] +
                  mat_A[27][24] * mat_B[24][20] +
                  mat_A[27][25] * mat_B[25][20] +
                  mat_A[27][26] * mat_B[26][20] +
                  mat_A[27][27] * mat_B[27][20] +
                  mat_A[27][28] * mat_B[28][20] +
                  mat_A[27][29] * mat_B[29][20] +
                  mat_A[27][30] * mat_B[30][20] +
                  mat_A[27][31] * mat_B[31][20];
    mat_C[27][21] <= 
                  mat_A[27][0] * mat_B[0][21] +
                  mat_A[27][1] * mat_B[1][21] +
                  mat_A[27][2] * mat_B[2][21] +
                  mat_A[27][3] * mat_B[3][21] +
                  mat_A[27][4] * mat_B[4][21] +
                  mat_A[27][5] * mat_B[5][21] +
                  mat_A[27][6] * mat_B[6][21] +
                  mat_A[27][7] * mat_B[7][21] +
                  mat_A[27][8] * mat_B[8][21] +
                  mat_A[27][9] * mat_B[9][21] +
                  mat_A[27][10] * mat_B[10][21] +
                  mat_A[27][11] * mat_B[11][21] +
                  mat_A[27][12] * mat_B[12][21] +
                  mat_A[27][13] * mat_B[13][21] +
                  mat_A[27][14] * mat_B[14][21] +
                  mat_A[27][15] * mat_B[15][21] +
                  mat_A[27][16] * mat_B[16][21] +
                  mat_A[27][17] * mat_B[17][21] +
                  mat_A[27][18] * mat_B[18][21] +
                  mat_A[27][19] * mat_B[19][21] +
                  mat_A[27][20] * mat_B[20][21] +
                  mat_A[27][21] * mat_B[21][21] +
                  mat_A[27][22] * mat_B[22][21] +
                  mat_A[27][23] * mat_B[23][21] +
                  mat_A[27][24] * mat_B[24][21] +
                  mat_A[27][25] * mat_B[25][21] +
                  mat_A[27][26] * mat_B[26][21] +
                  mat_A[27][27] * mat_B[27][21] +
                  mat_A[27][28] * mat_B[28][21] +
                  mat_A[27][29] * mat_B[29][21] +
                  mat_A[27][30] * mat_B[30][21] +
                  mat_A[27][31] * mat_B[31][21];
    mat_C[27][22] <= 
                  mat_A[27][0] * mat_B[0][22] +
                  mat_A[27][1] * mat_B[1][22] +
                  mat_A[27][2] * mat_B[2][22] +
                  mat_A[27][3] * mat_B[3][22] +
                  mat_A[27][4] * mat_B[4][22] +
                  mat_A[27][5] * mat_B[5][22] +
                  mat_A[27][6] * mat_B[6][22] +
                  mat_A[27][7] * mat_B[7][22] +
                  mat_A[27][8] * mat_B[8][22] +
                  mat_A[27][9] * mat_B[9][22] +
                  mat_A[27][10] * mat_B[10][22] +
                  mat_A[27][11] * mat_B[11][22] +
                  mat_A[27][12] * mat_B[12][22] +
                  mat_A[27][13] * mat_B[13][22] +
                  mat_A[27][14] * mat_B[14][22] +
                  mat_A[27][15] * mat_B[15][22] +
                  mat_A[27][16] * mat_B[16][22] +
                  mat_A[27][17] * mat_B[17][22] +
                  mat_A[27][18] * mat_B[18][22] +
                  mat_A[27][19] * mat_B[19][22] +
                  mat_A[27][20] * mat_B[20][22] +
                  mat_A[27][21] * mat_B[21][22] +
                  mat_A[27][22] * mat_B[22][22] +
                  mat_A[27][23] * mat_B[23][22] +
                  mat_A[27][24] * mat_B[24][22] +
                  mat_A[27][25] * mat_B[25][22] +
                  mat_A[27][26] * mat_B[26][22] +
                  mat_A[27][27] * mat_B[27][22] +
                  mat_A[27][28] * mat_B[28][22] +
                  mat_A[27][29] * mat_B[29][22] +
                  mat_A[27][30] * mat_B[30][22] +
                  mat_A[27][31] * mat_B[31][22];
    mat_C[27][23] <= 
                  mat_A[27][0] * mat_B[0][23] +
                  mat_A[27][1] * mat_B[1][23] +
                  mat_A[27][2] * mat_B[2][23] +
                  mat_A[27][3] * mat_B[3][23] +
                  mat_A[27][4] * mat_B[4][23] +
                  mat_A[27][5] * mat_B[5][23] +
                  mat_A[27][6] * mat_B[6][23] +
                  mat_A[27][7] * mat_B[7][23] +
                  mat_A[27][8] * mat_B[8][23] +
                  mat_A[27][9] * mat_B[9][23] +
                  mat_A[27][10] * mat_B[10][23] +
                  mat_A[27][11] * mat_B[11][23] +
                  mat_A[27][12] * mat_B[12][23] +
                  mat_A[27][13] * mat_B[13][23] +
                  mat_A[27][14] * mat_B[14][23] +
                  mat_A[27][15] * mat_B[15][23] +
                  mat_A[27][16] * mat_B[16][23] +
                  mat_A[27][17] * mat_B[17][23] +
                  mat_A[27][18] * mat_B[18][23] +
                  mat_A[27][19] * mat_B[19][23] +
                  mat_A[27][20] * mat_B[20][23] +
                  mat_A[27][21] * mat_B[21][23] +
                  mat_A[27][22] * mat_B[22][23] +
                  mat_A[27][23] * mat_B[23][23] +
                  mat_A[27][24] * mat_B[24][23] +
                  mat_A[27][25] * mat_B[25][23] +
                  mat_A[27][26] * mat_B[26][23] +
                  mat_A[27][27] * mat_B[27][23] +
                  mat_A[27][28] * mat_B[28][23] +
                  mat_A[27][29] * mat_B[29][23] +
                  mat_A[27][30] * mat_B[30][23] +
                  mat_A[27][31] * mat_B[31][23];
    mat_C[27][24] <= 
                  mat_A[27][0] * mat_B[0][24] +
                  mat_A[27][1] * mat_B[1][24] +
                  mat_A[27][2] * mat_B[2][24] +
                  mat_A[27][3] * mat_B[3][24] +
                  mat_A[27][4] * mat_B[4][24] +
                  mat_A[27][5] * mat_B[5][24] +
                  mat_A[27][6] * mat_B[6][24] +
                  mat_A[27][7] * mat_B[7][24] +
                  mat_A[27][8] * mat_B[8][24] +
                  mat_A[27][9] * mat_B[9][24] +
                  mat_A[27][10] * mat_B[10][24] +
                  mat_A[27][11] * mat_B[11][24] +
                  mat_A[27][12] * mat_B[12][24] +
                  mat_A[27][13] * mat_B[13][24] +
                  mat_A[27][14] * mat_B[14][24] +
                  mat_A[27][15] * mat_B[15][24] +
                  mat_A[27][16] * mat_B[16][24] +
                  mat_A[27][17] * mat_B[17][24] +
                  mat_A[27][18] * mat_B[18][24] +
                  mat_A[27][19] * mat_B[19][24] +
                  mat_A[27][20] * mat_B[20][24] +
                  mat_A[27][21] * mat_B[21][24] +
                  mat_A[27][22] * mat_B[22][24] +
                  mat_A[27][23] * mat_B[23][24] +
                  mat_A[27][24] * mat_B[24][24] +
                  mat_A[27][25] * mat_B[25][24] +
                  mat_A[27][26] * mat_B[26][24] +
                  mat_A[27][27] * mat_B[27][24] +
                  mat_A[27][28] * mat_B[28][24] +
                  mat_A[27][29] * mat_B[29][24] +
                  mat_A[27][30] * mat_B[30][24] +
                  mat_A[27][31] * mat_B[31][24];
    mat_C[27][25] <= 
                  mat_A[27][0] * mat_B[0][25] +
                  mat_A[27][1] * mat_B[1][25] +
                  mat_A[27][2] * mat_B[2][25] +
                  mat_A[27][3] * mat_B[3][25] +
                  mat_A[27][4] * mat_B[4][25] +
                  mat_A[27][5] * mat_B[5][25] +
                  mat_A[27][6] * mat_B[6][25] +
                  mat_A[27][7] * mat_B[7][25] +
                  mat_A[27][8] * mat_B[8][25] +
                  mat_A[27][9] * mat_B[9][25] +
                  mat_A[27][10] * mat_B[10][25] +
                  mat_A[27][11] * mat_B[11][25] +
                  mat_A[27][12] * mat_B[12][25] +
                  mat_A[27][13] * mat_B[13][25] +
                  mat_A[27][14] * mat_B[14][25] +
                  mat_A[27][15] * mat_B[15][25] +
                  mat_A[27][16] * mat_B[16][25] +
                  mat_A[27][17] * mat_B[17][25] +
                  mat_A[27][18] * mat_B[18][25] +
                  mat_A[27][19] * mat_B[19][25] +
                  mat_A[27][20] * mat_B[20][25] +
                  mat_A[27][21] * mat_B[21][25] +
                  mat_A[27][22] * mat_B[22][25] +
                  mat_A[27][23] * mat_B[23][25] +
                  mat_A[27][24] * mat_B[24][25] +
                  mat_A[27][25] * mat_B[25][25] +
                  mat_A[27][26] * mat_B[26][25] +
                  mat_A[27][27] * mat_B[27][25] +
                  mat_A[27][28] * mat_B[28][25] +
                  mat_A[27][29] * mat_B[29][25] +
                  mat_A[27][30] * mat_B[30][25] +
                  mat_A[27][31] * mat_B[31][25];
    mat_C[27][26] <= 
                  mat_A[27][0] * mat_B[0][26] +
                  mat_A[27][1] * mat_B[1][26] +
                  mat_A[27][2] * mat_B[2][26] +
                  mat_A[27][3] * mat_B[3][26] +
                  mat_A[27][4] * mat_B[4][26] +
                  mat_A[27][5] * mat_B[5][26] +
                  mat_A[27][6] * mat_B[6][26] +
                  mat_A[27][7] * mat_B[7][26] +
                  mat_A[27][8] * mat_B[8][26] +
                  mat_A[27][9] * mat_B[9][26] +
                  mat_A[27][10] * mat_B[10][26] +
                  mat_A[27][11] * mat_B[11][26] +
                  mat_A[27][12] * mat_B[12][26] +
                  mat_A[27][13] * mat_B[13][26] +
                  mat_A[27][14] * mat_B[14][26] +
                  mat_A[27][15] * mat_B[15][26] +
                  mat_A[27][16] * mat_B[16][26] +
                  mat_A[27][17] * mat_B[17][26] +
                  mat_A[27][18] * mat_B[18][26] +
                  mat_A[27][19] * mat_B[19][26] +
                  mat_A[27][20] * mat_B[20][26] +
                  mat_A[27][21] * mat_B[21][26] +
                  mat_A[27][22] * mat_B[22][26] +
                  mat_A[27][23] * mat_B[23][26] +
                  mat_A[27][24] * mat_B[24][26] +
                  mat_A[27][25] * mat_B[25][26] +
                  mat_A[27][26] * mat_B[26][26] +
                  mat_A[27][27] * mat_B[27][26] +
                  mat_A[27][28] * mat_B[28][26] +
                  mat_A[27][29] * mat_B[29][26] +
                  mat_A[27][30] * mat_B[30][26] +
                  mat_A[27][31] * mat_B[31][26];
    mat_C[27][27] <= 
                  mat_A[27][0] * mat_B[0][27] +
                  mat_A[27][1] * mat_B[1][27] +
                  mat_A[27][2] * mat_B[2][27] +
                  mat_A[27][3] * mat_B[3][27] +
                  mat_A[27][4] * mat_B[4][27] +
                  mat_A[27][5] * mat_B[5][27] +
                  mat_A[27][6] * mat_B[6][27] +
                  mat_A[27][7] * mat_B[7][27] +
                  mat_A[27][8] * mat_B[8][27] +
                  mat_A[27][9] * mat_B[9][27] +
                  mat_A[27][10] * mat_B[10][27] +
                  mat_A[27][11] * mat_B[11][27] +
                  mat_A[27][12] * mat_B[12][27] +
                  mat_A[27][13] * mat_B[13][27] +
                  mat_A[27][14] * mat_B[14][27] +
                  mat_A[27][15] * mat_B[15][27] +
                  mat_A[27][16] * mat_B[16][27] +
                  mat_A[27][17] * mat_B[17][27] +
                  mat_A[27][18] * mat_B[18][27] +
                  mat_A[27][19] * mat_B[19][27] +
                  mat_A[27][20] * mat_B[20][27] +
                  mat_A[27][21] * mat_B[21][27] +
                  mat_A[27][22] * mat_B[22][27] +
                  mat_A[27][23] * mat_B[23][27] +
                  mat_A[27][24] * mat_B[24][27] +
                  mat_A[27][25] * mat_B[25][27] +
                  mat_A[27][26] * mat_B[26][27] +
                  mat_A[27][27] * mat_B[27][27] +
                  mat_A[27][28] * mat_B[28][27] +
                  mat_A[27][29] * mat_B[29][27] +
                  mat_A[27][30] * mat_B[30][27] +
                  mat_A[27][31] * mat_B[31][27];
    mat_C[27][28] <= 
                  mat_A[27][0] * mat_B[0][28] +
                  mat_A[27][1] * mat_B[1][28] +
                  mat_A[27][2] * mat_B[2][28] +
                  mat_A[27][3] * mat_B[3][28] +
                  mat_A[27][4] * mat_B[4][28] +
                  mat_A[27][5] * mat_B[5][28] +
                  mat_A[27][6] * mat_B[6][28] +
                  mat_A[27][7] * mat_B[7][28] +
                  mat_A[27][8] * mat_B[8][28] +
                  mat_A[27][9] * mat_B[9][28] +
                  mat_A[27][10] * mat_B[10][28] +
                  mat_A[27][11] * mat_B[11][28] +
                  mat_A[27][12] * mat_B[12][28] +
                  mat_A[27][13] * mat_B[13][28] +
                  mat_A[27][14] * mat_B[14][28] +
                  mat_A[27][15] * mat_B[15][28] +
                  mat_A[27][16] * mat_B[16][28] +
                  mat_A[27][17] * mat_B[17][28] +
                  mat_A[27][18] * mat_B[18][28] +
                  mat_A[27][19] * mat_B[19][28] +
                  mat_A[27][20] * mat_B[20][28] +
                  mat_A[27][21] * mat_B[21][28] +
                  mat_A[27][22] * mat_B[22][28] +
                  mat_A[27][23] * mat_B[23][28] +
                  mat_A[27][24] * mat_B[24][28] +
                  mat_A[27][25] * mat_B[25][28] +
                  mat_A[27][26] * mat_B[26][28] +
                  mat_A[27][27] * mat_B[27][28] +
                  mat_A[27][28] * mat_B[28][28] +
                  mat_A[27][29] * mat_B[29][28] +
                  mat_A[27][30] * mat_B[30][28] +
                  mat_A[27][31] * mat_B[31][28];
    mat_C[27][29] <= 
                  mat_A[27][0] * mat_B[0][29] +
                  mat_A[27][1] * mat_B[1][29] +
                  mat_A[27][2] * mat_B[2][29] +
                  mat_A[27][3] * mat_B[3][29] +
                  mat_A[27][4] * mat_B[4][29] +
                  mat_A[27][5] * mat_B[5][29] +
                  mat_A[27][6] * mat_B[6][29] +
                  mat_A[27][7] * mat_B[7][29] +
                  mat_A[27][8] * mat_B[8][29] +
                  mat_A[27][9] * mat_B[9][29] +
                  mat_A[27][10] * mat_B[10][29] +
                  mat_A[27][11] * mat_B[11][29] +
                  mat_A[27][12] * mat_B[12][29] +
                  mat_A[27][13] * mat_B[13][29] +
                  mat_A[27][14] * mat_B[14][29] +
                  mat_A[27][15] * mat_B[15][29] +
                  mat_A[27][16] * mat_B[16][29] +
                  mat_A[27][17] * mat_B[17][29] +
                  mat_A[27][18] * mat_B[18][29] +
                  mat_A[27][19] * mat_B[19][29] +
                  mat_A[27][20] * mat_B[20][29] +
                  mat_A[27][21] * mat_B[21][29] +
                  mat_A[27][22] * mat_B[22][29] +
                  mat_A[27][23] * mat_B[23][29] +
                  mat_A[27][24] * mat_B[24][29] +
                  mat_A[27][25] * mat_B[25][29] +
                  mat_A[27][26] * mat_B[26][29] +
                  mat_A[27][27] * mat_B[27][29] +
                  mat_A[27][28] * mat_B[28][29] +
                  mat_A[27][29] * mat_B[29][29] +
                  mat_A[27][30] * mat_B[30][29] +
                  mat_A[27][31] * mat_B[31][29];
    mat_C[27][30] <= 
                  mat_A[27][0] * mat_B[0][30] +
                  mat_A[27][1] * mat_B[1][30] +
                  mat_A[27][2] * mat_B[2][30] +
                  mat_A[27][3] * mat_B[3][30] +
                  mat_A[27][4] * mat_B[4][30] +
                  mat_A[27][5] * mat_B[5][30] +
                  mat_A[27][6] * mat_B[6][30] +
                  mat_A[27][7] * mat_B[7][30] +
                  mat_A[27][8] * mat_B[8][30] +
                  mat_A[27][9] * mat_B[9][30] +
                  mat_A[27][10] * mat_B[10][30] +
                  mat_A[27][11] * mat_B[11][30] +
                  mat_A[27][12] * mat_B[12][30] +
                  mat_A[27][13] * mat_B[13][30] +
                  mat_A[27][14] * mat_B[14][30] +
                  mat_A[27][15] * mat_B[15][30] +
                  mat_A[27][16] * mat_B[16][30] +
                  mat_A[27][17] * mat_B[17][30] +
                  mat_A[27][18] * mat_B[18][30] +
                  mat_A[27][19] * mat_B[19][30] +
                  mat_A[27][20] * mat_B[20][30] +
                  mat_A[27][21] * mat_B[21][30] +
                  mat_A[27][22] * mat_B[22][30] +
                  mat_A[27][23] * mat_B[23][30] +
                  mat_A[27][24] * mat_B[24][30] +
                  mat_A[27][25] * mat_B[25][30] +
                  mat_A[27][26] * mat_B[26][30] +
                  mat_A[27][27] * mat_B[27][30] +
                  mat_A[27][28] * mat_B[28][30] +
                  mat_A[27][29] * mat_B[29][30] +
                  mat_A[27][30] * mat_B[30][30] +
                  mat_A[27][31] * mat_B[31][30];
    mat_C[27][31] <= 
                  mat_A[27][0] * mat_B[0][31] +
                  mat_A[27][1] * mat_B[1][31] +
                  mat_A[27][2] * mat_B[2][31] +
                  mat_A[27][3] * mat_B[3][31] +
                  mat_A[27][4] * mat_B[4][31] +
                  mat_A[27][5] * mat_B[5][31] +
                  mat_A[27][6] * mat_B[6][31] +
                  mat_A[27][7] * mat_B[7][31] +
                  mat_A[27][8] * mat_B[8][31] +
                  mat_A[27][9] * mat_B[9][31] +
                  mat_A[27][10] * mat_B[10][31] +
                  mat_A[27][11] * mat_B[11][31] +
                  mat_A[27][12] * mat_B[12][31] +
                  mat_A[27][13] * mat_B[13][31] +
                  mat_A[27][14] * mat_B[14][31] +
                  mat_A[27][15] * mat_B[15][31] +
                  mat_A[27][16] * mat_B[16][31] +
                  mat_A[27][17] * mat_B[17][31] +
                  mat_A[27][18] * mat_B[18][31] +
                  mat_A[27][19] * mat_B[19][31] +
                  mat_A[27][20] * mat_B[20][31] +
                  mat_A[27][21] * mat_B[21][31] +
                  mat_A[27][22] * mat_B[22][31] +
                  mat_A[27][23] * mat_B[23][31] +
                  mat_A[27][24] * mat_B[24][31] +
                  mat_A[27][25] * mat_B[25][31] +
                  mat_A[27][26] * mat_B[26][31] +
                  mat_A[27][27] * mat_B[27][31] +
                  mat_A[27][28] * mat_B[28][31] +
                  mat_A[27][29] * mat_B[29][31] +
                  mat_A[27][30] * mat_B[30][31] +
                  mat_A[27][31] * mat_B[31][31];
    mat_C[28][0] <= 
                  mat_A[28][0] * mat_B[0][0] +
                  mat_A[28][1] * mat_B[1][0] +
                  mat_A[28][2] * mat_B[2][0] +
                  mat_A[28][3] * mat_B[3][0] +
                  mat_A[28][4] * mat_B[4][0] +
                  mat_A[28][5] * mat_B[5][0] +
                  mat_A[28][6] * mat_B[6][0] +
                  mat_A[28][7] * mat_B[7][0] +
                  mat_A[28][8] * mat_B[8][0] +
                  mat_A[28][9] * mat_B[9][0] +
                  mat_A[28][10] * mat_B[10][0] +
                  mat_A[28][11] * mat_B[11][0] +
                  mat_A[28][12] * mat_B[12][0] +
                  mat_A[28][13] * mat_B[13][0] +
                  mat_A[28][14] * mat_B[14][0] +
                  mat_A[28][15] * mat_B[15][0] +
                  mat_A[28][16] * mat_B[16][0] +
                  mat_A[28][17] * mat_B[17][0] +
                  mat_A[28][18] * mat_B[18][0] +
                  mat_A[28][19] * mat_B[19][0] +
                  mat_A[28][20] * mat_B[20][0] +
                  mat_A[28][21] * mat_B[21][0] +
                  mat_A[28][22] * mat_B[22][0] +
                  mat_A[28][23] * mat_B[23][0] +
                  mat_A[28][24] * mat_B[24][0] +
                  mat_A[28][25] * mat_B[25][0] +
                  mat_A[28][26] * mat_B[26][0] +
                  mat_A[28][27] * mat_B[27][0] +
                  mat_A[28][28] * mat_B[28][0] +
                  mat_A[28][29] * mat_B[29][0] +
                  mat_A[28][30] * mat_B[30][0] +
                  mat_A[28][31] * mat_B[31][0];
    mat_C[28][1] <= 
                  mat_A[28][0] * mat_B[0][1] +
                  mat_A[28][1] * mat_B[1][1] +
                  mat_A[28][2] * mat_B[2][1] +
                  mat_A[28][3] * mat_B[3][1] +
                  mat_A[28][4] * mat_B[4][1] +
                  mat_A[28][5] * mat_B[5][1] +
                  mat_A[28][6] * mat_B[6][1] +
                  mat_A[28][7] * mat_B[7][1] +
                  mat_A[28][8] * mat_B[8][1] +
                  mat_A[28][9] * mat_B[9][1] +
                  mat_A[28][10] * mat_B[10][1] +
                  mat_A[28][11] * mat_B[11][1] +
                  mat_A[28][12] * mat_B[12][1] +
                  mat_A[28][13] * mat_B[13][1] +
                  mat_A[28][14] * mat_B[14][1] +
                  mat_A[28][15] * mat_B[15][1] +
                  mat_A[28][16] * mat_B[16][1] +
                  mat_A[28][17] * mat_B[17][1] +
                  mat_A[28][18] * mat_B[18][1] +
                  mat_A[28][19] * mat_B[19][1] +
                  mat_A[28][20] * mat_B[20][1] +
                  mat_A[28][21] * mat_B[21][1] +
                  mat_A[28][22] * mat_B[22][1] +
                  mat_A[28][23] * mat_B[23][1] +
                  mat_A[28][24] * mat_B[24][1] +
                  mat_A[28][25] * mat_B[25][1] +
                  mat_A[28][26] * mat_B[26][1] +
                  mat_A[28][27] * mat_B[27][1] +
                  mat_A[28][28] * mat_B[28][1] +
                  mat_A[28][29] * mat_B[29][1] +
                  mat_A[28][30] * mat_B[30][1] +
                  mat_A[28][31] * mat_B[31][1];
    mat_C[28][2] <= 
                  mat_A[28][0] * mat_B[0][2] +
                  mat_A[28][1] * mat_B[1][2] +
                  mat_A[28][2] * mat_B[2][2] +
                  mat_A[28][3] * mat_B[3][2] +
                  mat_A[28][4] * mat_B[4][2] +
                  mat_A[28][5] * mat_B[5][2] +
                  mat_A[28][6] * mat_B[6][2] +
                  mat_A[28][7] * mat_B[7][2] +
                  mat_A[28][8] * mat_B[8][2] +
                  mat_A[28][9] * mat_B[9][2] +
                  mat_A[28][10] * mat_B[10][2] +
                  mat_A[28][11] * mat_B[11][2] +
                  mat_A[28][12] * mat_B[12][2] +
                  mat_A[28][13] * mat_B[13][2] +
                  mat_A[28][14] * mat_B[14][2] +
                  mat_A[28][15] * mat_B[15][2] +
                  mat_A[28][16] * mat_B[16][2] +
                  mat_A[28][17] * mat_B[17][2] +
                  mat_A[28][18] * mat_B[18][2] +
                  mat_A[28][19] * mat_B[19][2] +
                  mat_A[28][20] * mat_B[20][2] +
                  mat_A[28][21] * mat_B[21][2] +
                  mat_A[28][22] * mat_B[22][2] +
                  mat_A[28][23] * mat_B[23][2] +
                  mat_A[28][24] * mat_B[24][2] +
                  mat_A[28][25] * mat_B[25][2] +
                  mat_A[28][26] * mat_B[26][2] +
                  mat_A[28][27] * mat_B[27][2] +
                  mat_A[28][28] * mat_B[28][2] +
                  mat_A[28][29] * mat_B[29][2] +
                  mat_A[28][30] * mat_B[30][2] +
                  mat_A[28][31] * mat_B[31][2];
    mat_C[28][3] <= 
                  mat_A[28][0] * mat_B[0][3] +
                  mat_A[28][1] * mat_B[1][3] +
                  mat_A[28][2] * mat_B[2][3] +
                  mat_A[28][3] * mat_B[3][3] +
                  mat_A[28][4] * mat_B[4][3] +
                  mat_A[28][5] * mat_B[5][3] +
                  mat_A[28][6] * mat_B[6][3] +
                  mat_A[28][7] * mat_B[7][3] +
                  mat_A[28][8] * mat_B[8][3] +
                  mat_A[28][9] * mat_B[9][3] +
                  mat_A[28][10] * mat_B[10][3] +
                  mat_A[28][11] * mat_B[11][3] +
                  mat_A[28][12] * mat_B[12][3] +
                  mat_A[28][13] * mat_B[13][3] +
                  mat_A[28][14] * mat_B[14][3] +
                  mat_A[28][15] * mat_B[15][3] +
                  mat_A[28][16] * mat_B[16][3] +
                  mat_A[28][17] * mat_B[17][3] +
                  mat_A[28][18] * mat_B[18][3] +
                  mat_A[28][19] * mat_B[19][3] +
                  mat_A[28][20] * mat_B[20][3] +
                  mat_A[28][21] * mat_B[21][3] +
                  mat_A[28][22] * mat_B[22][3] +
                  mat_A[28][23] * mat_B[23][3] +
                  mat_A[28][24] * mat_B[24][3] +
                  mat_A[28][25] * mat_B[25][3] +
                  mat_A[28][26] * mat_B[26][3] +
                  mat_A[28][27] * mat_B[27][3] +
                  mat_A[28][28] * mat_B[28][3] +
                  mat_A[28][29] * mat_B[29][3] +
                  mat_A[28][30] * mat_B[30][3] +
                  mat_A[28][31] * mat_B[31][3];
    mat_C[28][4] <= 
                  mat_A[28][0] * mat_B[0][4] +
                  mat_A[28][1] * mat_B[1][4] +
                  mat_A[28][2] * mat_B[2][4] +
                  mat_A[28][3] * mat_B[3][4] +
                  mat_A[28][4] * mat_B[4][4] +
                  mat_A[28][5] * mat_B[5][4] +
                  mat_A[28][6] * mat_B[6][4] +
                  mat_A[28][7] * mat_B[7][4] +
                  mat_A[28][8] * mat_B[8][4] +
                  mat_A[28][9] * mat_B[9][4] +
                  mat_A[28][10] * mat_B[10][4] +
                  mat_A[28][11] * mat_B[11][4] +
                  mat_A[28][12] * mat_B[12][4] +
                  mat_A[28][13] * mat_B[13][4] +
                  mat_A[28][14] * mat_B[14][4] +
                  mat_A[28][15] * mat_B[15][4] +
                  mat_A[28][16] * mat_B[16][4] +
                  mat_A[28][17] * mat_B[17][4] +
                  mat_A[28][18] * mat_B[18][4] +
                  mat_A[28][19] * mat_B[19][4] +
                  mat_A[28][20] * mat_B[20][4] +
                  mat_A[28][21] * mat_B[21][4] +
                  mat_A[28][22] * mat_B[22][4] +
                  mat_A[28][23] * mat_B[23][4] +
                  mat_A[28][24] * mat_B[24][4] +
                  mat_A[28][25] * mat_B[25][4] +
                  mat_A[28][26] * mat_B[26][4] +
                  mat_A[28][27] * mat_B[27][4] +
                  mat_A[28][28] * mat_B[28][4] +
                  mat_A[28][29] * mat_B[29][4] +
                  mat_A[28][30] * mat_B[30][4] +
                  mat_A[28][31] * mat_B[31][4];
    mat_C[28][5] <= 
                  mat_A[28][0] * mat_B[0][5] +
                  mat_A[28][1] * mat_B[1][5] +
                  mat_A[28][2] * mat_B[2][5] +
                  mat_A[28][3] * mat_B[3][5] +
                  mat_A[28][4] * mat_B[4][5] +
                  mat_A[28][5] * mat_B[5][5] +
                  mat_A[28][6] * mat_B[6][5] +
                  mat_A[28][7] * mat_B[7][5] +
                  mat_A[28][8] * mat_B[8][5] +
                  mat_A[28][9] * mat_B[9][5] +
                  mat_A[28][10] * mat_B[10][5] +
                  mat_A[28][11] * mat_B[11][5] +
                  mat_A[28][12] * mat_B[12][5] +
                  mat_A[28][13] * mat_B[13][5] +
                  mat_A[28][14] * mat_B[14][5] +
                  mat_A[28][15] * mat_B[15][5] +
                  mat_A[28][16] * mat_B[16][5] +
                  mat_A[28][17] * mat_B[17][5] +
                  mat_A[28][18] * mat_B[18][5] +
                  mat_A[28][19] * mat_B[19][5] +
                  mat_A[28][20] * mat_B[20][5] +
                  mat_A[28][21] * mat_B[21][5] +
                  mat_A[28][22] * mat_B[22][5] +
                  mat_A[28][23] * mat_B[23][5] +
                  mat_A[28][24] * mat_B[24][5] +
                  mat_A[28][25] * mat_B[25][5] +
                  mat_A[28][26] * mat_B[26][5] +
                  mat_A[28][27] * mat_B[27][5] +
                  mat_A[28][28] * mat_B[28][5] +
                  mat_A[28][29] * mat_B[29][5] +
                  mat_A[28][30] * mat_B[30][5] +
                  mat_A[28][31] * mat_B[31][5];
    mat_C[28][6] <= 
                  mat_A[28][0] * mat_B[0][6] +
                  mat_A[28][1] * mat_B[1][6] +
                  mat_A[28][2] * mat_B[2][6] +
                  mat_A[28][3] * mat_B[3][6] +
                  mat_A[28][4] * mat_B[4][6] +
                  mat_A[28][5] * mat_B[5][6] +
                  mat_A[28][6] * mat_B[6][6] +
                  mat_A[28][7] * mat_B[7][6] +
                  mat_A[28][8] * mat_B[8][6] +
                  mat_A[28][9] * mat_B[9][6] +
                  mat_A[28][10] * mat_B[10][6] +
                  mat_A[28][11] * mat_B[11][6] +
                  mat_A[28][12] * mat_B[12][6] +
                  mat_A[28][13] * mat_B[13][6] +
                  mat_A[28][14] * mat_B[14][6] +
                  mat_A[28][15] * mat_B[15][6] +
                  mat_A[28][16] * mat_B[16][6] +
                  mat_A[28][17] * mat_B[17][6] +
                  mat_A[28][18] * mat_B[18][6] +
                  mat_A[28][19] * mat_B[19][6] +
                  mat_A[28][20] * mat_B[20][6] +
                  mat_A[28][21] * mat_B[21][6] +
                  mat_A[28][22] * mat_B[22][6] +
                  mat_A[28][23] * mat_B[23][6] +
                  mat_A[28][24] * mat_B[24][6] +
                  mat_A[28][25] * mat_B[25][6] +
                  mat_A[28][26] * mat_B[26][6] +
                  mat_A[28][27] * mat_B[27][6] +
                  mat_A[28][28] * mat_B[28][6] +
                  mat_A[28][29] * mat_B[29][6] +
                  mat_A[28][30] * mat_B[30][6] +
                  mat_A[28][31] * mat_B[31][6];
    mat_C[28][7] <= 
                  mat_A[28][0] * mat_B[0][7] +
                  mat_A[28][1] * mat_B[1][7] +
                  mat_A[28][2] * mat_B[2][7] +
                  mat_A[28][3] * mat_B[3][7] +
                  mat_A[28][4] * mat_B[4][7] +
                  mat_A[28][5] * mat_B[5][7] +
                  mat_A[28][6] * mat_B[6][7] +
                  mat_A[28][7] * mat_B[7][7] +
                  mat_A[28][8] * mat_B[8][7] +
                  mat_A[28][9] * mat_B[9][7] +
                  mat_A[28][10] * mat_B[10][7] +
                  mat_A[28][11] * mat_B[11][7] +
                  mat_A[28][12] * mat_B[12][7] +
                  mat_A[28][13] * mat_B[13][7] +
                  mat_A[28][14] * mat_B[14][7] +
                  mat_A[28][15] * mat_B[15][7] +
                  mat_A[28][16] * mat_B[16][7] +
                  mat_A[28][17] * mat_B[17][7] +
                  mat_A[28][18] * mat_B[18][7] +
                  mat_A[28][19] * mat_B[19][7] +
                  mat_A[28][20] * mat_B[20][7] +
                  mat_A[28][21] * mat_B[21][7] +
                  mat_A[28][22] * mat_B[22][7] +
                  mat_A[28][23] * mat_B[23][7] +
                  mat_A[28][24] * mat_B[24][7] +
                  mat_A[28][25] * mat_B[25][7] +
                  mat_A[28][26] * mat_B[26][7] +
                  mat_A[28][27] * mat_B[27][7] +
                  mat_A[28][28] * mat_B[28][7] +
                  mat_A[28][29] * mat_B[29][7] +
                  mat_A[28][30] * mat_B[30][7] +
                  mat_A[28][31] * mat_B[31][7];
    mat_C[28][8] <= 
                  mat_A[28][0] * mat_B[0][8] +
                  mat_A[28][1] * mat_B[1][8] +
                  mat_A[28][2] * mat_B[2][8] +
                  mat_A[28][3] * mat_B[3][8] +
                  mat_A[28][4] * mat_B[4][8] +
                  mat_A[28][5] * mat_B[5][8] +
                  mat_A[28][6] * mat_B[6][8] +
                  mat_A[28][7] * mat_B[7][8] +
                  mat_A[28][8] * mat_B[8][8] +
                  mat_A[28][9] * mat_B[9][8] +
                  mat_A[28][10] * mat_B[10][8] +
                  mat_A[28][11] * mat_B[11][8] +
                  mat_A[28][12] * mat_B[12][8] +
                  mat_A[28][13] * mat_B[13][8] +
                  mat_A[28][14] * mat_B[14][8] +
                  mat_A[28][15] * mat_B[15][8] +
                  mat_A[28][16] * mat_B[16][8] +
                  mat_A[28][17] * mat_B[17][8] +
                  mat_A[28][18] * mat_B[18][8] +
                  mat_A[28][19] * mat_B[19][8] +
                  mat_A[28][20] * mat_B[20][8] +
                  mat_A[28][21] * mat_B[21][8] +
                  mat_A[28][22] * mat_B[22][8] +
                  mat_A[28][23] * mat_B[23][8] +
                  mat_A[28][24] * mat_B[24][8] +
                  mat_A[28][25] * mat_B[25][8] +
                  mat_A[28][26] * mat_B[26][8] +
                  mat_A[28][27] * mat_B[27][8] +
                  mat_A[28][28] * mat_B[28][8] +
                  mat_A[28][29] * mat_B[29][8] +
                  mat_A[28][30] * mat_B[30][8] +
                  mat_A[28][31] * mat_B[31][8];
    mat_C[28][9] <= 
                  mat_A[28][0] * mat_B[0][9] +
                  mat_A[28][1] * mat_B[1][9] +
                  mat_A[28][2] * mat_B[2][9] +
                  mat_A[28][3] * mat_B[3][9] +
                  mat_A[28][4] * mat_B[4][9] +
                  mat_A[28][5] * mat_B[5][9] +
                  mat_A[28][6] * mat_B[6][9] +
                  mat_A[28][7] * mat_B[7][9] +
                  mat_A[28][8] * mat_B[8][9] +
                  mat_A[28][9] * mat_B[9][9] +
                  mat_A[28][10] * mat_B[10][9] +
                  mat_A[28][11] * mat_B[11][9] +
                  mat_A[28][12] * mat_B[12][9] +
                  mat_A[28][13] * mat_B[13][9] +
                  mat_A[28][14] * mat_B[14][9] +
                  mat_A[28][15] * mat_B[15][9] +
                  mat_A[28][16] * mat_B[16][9] +
                  mat_A[28][17] * mat_B[17][9] +
                  mat_A[28][18] * mat_B[18][9] +
                  mat_A[28][19] * mat_B[19][9] +
                  mat_A[28][20] * mat_B[20][9] +
                  mat_A[28][21] * mat_B[21][9] +
                  mat_A[28][22] * mat_B[22][9] +
                  mat_A[28][23] * mat_B[23][9] +
                  mat_A[28][24] * mat_B[24][9] +
                  mat_A[28][25] * mat_B[25][9] +
                  mat_A[28][26] * mat_B[26][9] +
                  mat_A[28][27] * mat_B[27][9] +
                  mat_A[28][28] * mat_B[28][9] +
                  mat_A[28][29] * mat_B[29][9] +
                  mat_A[28][30] * mat_B[30][9] +
                  mat_A[28][31] * mat_B[31][9];
    mat_C[28][10] <= 
                  mat_A[28][0] * mat_B[0][10] +
                  mat_A[28][1] * mat_B[1][10] +
                  mat_A[28][2] * mat_B[2][10] +
                  mat_A[28][3] * mat_B[3][10] +
                  mat_A[28][4] * mat_B[4][10] +
                  mat_A[28][5] * mat_B[5][10] +
                  mat_A[28][6] * mat_B[6][10] +
                  mat_A[28][7] * mat_B[7][10] +
                  mat_A[28][8] * mat_B[8][10] +
                  mat_A[28][9] * mat_B[9][10] +
                  mat_A[28][10] * mat_B[10][10] +
                  mat_A[28][11] * mat_B[11][10] +
                  mat_A[28][12] * mat_B[12][10] +
                  mat_A[28][13] * mat_B[13][10] +
                  mat_A[28][14] * mat_B[14][10] +
                  mat_A[28][15] * mat_B[15][10] +
                  mat_A[28][16] * mat_B[16][10] +
                  mat_A[28][17] * mat_B[17][10] +
                  mat_A[28][18] * mat_B[18][10] +
                  mat_A[28][19] * mat_B[19][10] +
                  mat_A[28][20] * mat_B[20][10] +
                  mat_A[28][21] * mat_B[21][10] +
                  mat_A[28][22] * mat_B[22][10] +
                  mat_A[28][23] * mat_B[23][10] +
                  mat_A[28][24] * mat_B[24][10] +
                  mat_A[28][25] * mat_B[25][10] +
                  mat_A[28][26] * mat_B[26][10] +
                  mat_A[28][27] * mat_B[27][10] +
                  mat_A[28][28] * mat_B[28][10] +
                  mat_A[28][29] * mat_B[29][10] +
                  mat_A[28][30] * mat_B[30][10] +
                  mat_A[28][31] * mat_B[31][10];
    mat_C[28][11] <= 
                  mat_A[28][0] * mat_B[0][11] +
                  mat_A[28][1] * mat_B[1][11] +
                  mat_A[28][2] * mat_B[2][11] +
                  mat_A[28][3] * mat_B[3][11] +
                  mat_A[28][4] * mat_B[4][11] +
                  mat_A[28][5] * mat_B[5][11] +
                  mat_A[28][6] * mat_B[6][11] +
                  mat_A[28][7] * mat_B[7][11] +
                  mat_A[28][8] * mat_B[8][11] +
                  mat_A[28][9] * mat_B[9][11] +
                  mat_A[28][10] * mat_B[10][11] +
                  mat_A[28][11] * mat_B[11][11] +
                  mat_A[28][12] * mat_B[12][11] +
                  mat_A[28][13] * mat_B[13][11] +
                  mat_A[28][14] * mat_B[14][11] +
                  mat_A[28][15] * mat_B[15][11] +
                  mat_A[28][16] * mat_B[16][11] +
                  mat_A[28][17] * mat_B[17][11] +
                  mat_A[28][18] * mat_B[18][11] +
                  mat_A[28][19] * mat_B[19][11] +
                  mat_A[28][20] * mat_B[20][11] +
                  mat_A[28][21] * mat_B[21][11] +
                  mat_A[28][22] * mat_B[22][11] +
                  mat_A[28][23] * mat_B[23][11] +
                  mat_A[28][24] * mat_B[24][11] +
                  mat_A[28][25] * mat_B[25][11] +
                  mat_A[28][26] * mat_B[26][11] +
                  mat_A[28][27] * mat_B[27][11] +
                  mat_A[28][28] * mat_B[28][11] +
                  mat_A[28][29] * mat_B[29][11] +
                  mat_A[28][30] * mat_B[30][11] +
                  mat_A[28][31] * mat_B[31][11];
    mat_C[28][12] <= 
                  mat_A[28][0] * mat_B[0][12] +
                  mat_A[28][1] * mat_B[1][12] +
                  mat_A[28][2] * mat_B[2][12] +
                  mat_A[28][3] * mat_B[3][12] +
                  mat_A[28][4] * mat_B[4][12] +
                  mat_A[28][5] * mat_B[5][12] +
                  mat_A[28][6] * mat_B[6][12] +
                  mat_A[28][7] * mat_B[7][12] +
                  mat_A[28][8] * mat_B[8][12] +
                  mat_A[28][9] * mat_B[9][12] +
                  mat_A[28][10] * mat_B[10][12] +
                  mat_A[28][11] * mat_B[11][12] +
                  mat_A[28][12] * mat_B[12][12] +
                  mat_A[28][13] * mat_B[13][12] +
                  mat_A[28][14] * mat_B[14][12] +
                  mat_A[28][15] * mat_B[15][12] +
                  mat_A[28][16] * mat_B[16][12] +
                  mat_A[28][17] * mat_B[17][12] +
                  mat_A[28][18] * mat_B[18][12] +
                  mat_A[28][19] * mat_B[19][12] +
                  mat_A[28][20] * mat_B[20][12] +
                  mat_A[28][21] * mat_B[21][12] +
                  mat_A[28][22] * mat_B[22][12] +
                  mat_A[28][23] * mat_B[23][12] +
                  mat_A[28][24] * mat_B[24][12] +
                  mat_A[28][25] * mat_B[25][12] +
                  mat_A[28][26] * mat_B[26][12] +
                  mat_A[28][27] * mat_B[27][12] +
                  mat_A[28][28] * mat_B[28][12] +
                  mat_A[28][29] * mat_B[29][12] +
                  mat_A[28][30] * mat_B[30][12] +
                  mat_A[28][31] * mat_B[31][12];
    mat_C[28][13] <= 
                  mat_A[28][0] * mat_B[0][13] +
                  mat_A[28][1] * mat_B[1][13] +
                  mat_A[28][2] * mat_B[2][13] +
                  mat_A[28][3] * mat_B[3][13] +
                  mat_A[28][4] * mat_B[4][13] +
                  mat_A[28][5] * mat_B[5][13] +
                  mat_A[28][6] * mat_B[6][13] +
                  mat_A[28][7] * mat_B[7][13] +
                  mat_A[28][8] * mat_B[8][13] +
                  mat_A[28][9] * mat_B[9][13] +
                  mat_A[28][10] * mat_B[10][13] +
                  mat_A[28][11] * mat_B[11][13] +
                  mat_A[28][12] * mat_B[12][13] +
                  mat_A[28][13] * mat_B[13][13] +
                  mat_A[28][14] * mat_B[14][13] +
                  mat_A[28][15] * mat_B[15][13] +
                  mat_A[28][16] * mat_B[16][13] +
                  mat_A[28][17] * mat_B[17][13] +
                  mat_A[28][18] * mat_B[18][13] +
                  mat_A[28][19] * mat_B[19][13] +
                  mat_A[28][20] * mat_B[20][13] +
                  mat_A[28][21] * mat_B[21][13] +
                  mat_A[28][22] * mat_B[22][13] +
                  mat_A[28][23] * mat_B[23][13] +
                  mat_A[28][24] * mat_B[24][13] +
                  mat_A[28][25] * mat_B[25][13] +
                  mat_A[28][26] * mat_B[26][13] +
                  mat_A[28][27] * mat_B[27][13] +
                  mat_A[28][28] * mat_B[28][13] +
                  mat_A[28][29] * mat_B[29][13] +
                  mat_A[28][30] * mat_B[30][13] +
                  mat_A[28][31] * mat_B[31][13];
    mat_C[28][14] <= 
                  mat_A[28][0] * mat_B[0][14] +
                  mat_A[28][1] * mat_B[1][14] +
                  mat_A[28][2] * mat_B[2][14] +
                  mat_A[28][3] * mat_B[3][14] +
                  mat_A[28][4] * mat_B[4][14] +
                  mat_A[28][5] * mat_B[5][14] +
                  mat_A[28][6] * mat_B[6][14] +
                  mat_A[28][7] * mat_B[7][14] +
                  mat_A[28][8] * mat_B[8][14] +
                  mat_A[28][9] * mat_B[9][14] +
                  mat_A[28][10] * mat_B[10][14] +
                  mat_A[28][11] * mat_B[11][14] +
                  mat_A[28][12] * mat_B[12][14] +
                  mat_A[28][13] * mat_B[13][14] +
                  mat_A[28][14] * mat_B[14][14] +
                  mat_A[28][15] * mat_B[15][14] +
                  mat_A[28][16] * mat_B[16][14] +
                  mat_A[28][17] * mat_B[17][14] +
                  mat_A[28][18] * mat_B[18][14] +
                  mat_A[28][19] * mat_B[19][14] +
                  mat_A[28][20] * mat_B[20][14] +
                  mat_A[28][21] * mat_B[21][14] +
                  mat_A[28][22] * mat_B[22][14] +
                  mat_A[28][23] * mat_B[23][14] +
                  mat_A[28][24] * mat_B[24][14] +
                  mat_A[28][25] * mat_B[25][14] +
                  mat_A[28][26] * mat_B[26][14] +
                  mat_A[28][27] * mat_B[27][14] +
                  mat_A[28][28] * mat_B[28][14] +
                  mat_A[28][29] * mat_B[29][14] +
                  mat_A[28][30] * mat_B[30][14] +
                  mat_A[28][31] * mat_B[31][14];
    mat_C[28][15] <= 
                  mat_A[28][0] * mat_B[0][15] +
                  mat_A[28][1] * mat_B[1][15] +
                  mat_A[28][2] * mat_B[2][15] +
                  mat_A[28][3] * mat_B[3][15] +
                  mat_A[28][4] * mat_B[4][15] +
                  mat_A[28][5] * mat_B[5][15] +
                  mat_A[28][6] * mat_B[6][15] +
                  mat_A[28][7] * mat_B[7][15] +
                  mat_A[28][8] * mat_B[8][15] +
                  mat_A[28][9] * mat_B[9][15] +
                  mat_A[28][10] * mat_B[10][15] +
                  mat_A[28][11] * mat_B[11][15] +
                  mat_A[28][12] * mat_B[12][15] +
                  mat_A[28][13] * mat_B[13][15] +
                  mat_A[28][14] * mat_B[14][15] +
                  mat_A[28][15] * mat_B[15][15] +
                  mat_A[28][16] * mat_B[16][15] +
                  mat_A[28][17] * mat_B[17][15] +
                  mat_A[28][18] * mat_B[18][15] +
                  mat_A[28][19] * mat_B[19][15] +
                  mat_A[28][20] * mat_B[20][15] +
                  mat_A[28][21] * mat_B[21][15] +
                  mat_A[28][22] * mat_B[22][15] +
                  mat_A[28][23] * mat_B[23][15] +
                  mat_A[28][24] * mat_B[24][15] +
                  mat_A[28][25] * mat_B[25][15] +
                  mat_A[28][26] * mat_B[26][15] +
                  mat_A[28][27] * mat_B[27][15] +
                  mat_A[28][28] * mat_B[28][15] +
                  mat_A[28][29] * mat_B[29][15] +
                  mat_A[28][30] * mat_B[30][15] +
                  mat_A[28][31] * mat_B[31][15];
    mat_C[28][16] <= 
                  mat_A[28][0] * mat_B[0][16] +
                  mat_A[28][1] * mat_B[1][16] +
                  mat_A[28][2] * mat_B[2][16] +
                  mat_A[28][3] * mat_B[3][16] +
                  mat_A[28][4] * mat_B[4][16] +
                  mat_A[28][5] * mat_B[5][16] +
                  mat_A[28][6] * mat_B[6][16] +
                  mat_A[28][7] * mat_B[7][16] +
                  mat_A[28][8] * mat_B[8][16] +
                  mat_A[28][9] * mat_B[9][16] +
                  mat_A[28][10] * mat_B[10][16] +
                  mat_A[28][11] * mat_B[11][16] +
                  mat_A[28][12] * mat_B[12][16] +
                  mat_A[28][13] * mat_B[13][16] +
                  mat_A[28][14] * mat_B[14][16] +
                  mat_A[28][15] * mat_B[15][16] +
                  mat_A[28][16] * mat_B[16][16] +
                  mat_A[28][17] * mat_B[17][16] +
                  mat_A[28][18] * mat_B[18][16] +
                  mat_A[28][19] * mat_B[19][16] +
                  mat_A[28][20] * mat_B[20][16] +
                  mat_A[28][21] * mat_B[21][16] +
                  mat_A[28][22] * mat_B[22][16] +
                  mat_A[28][23] * mat_B[23][16] +
                  mat_A[28][24] * mat_B[24][16] +
                  mat_A[28][25] * mat_B[25][16] +
                  mat_A[28][26] * mat_B[26][16] +
                  mat_A[28][27] * mat_B[27][16] +
                  mat_A[28][28] * mat_B[28][16] +
                  mat_A[28][29] * mat_B[29][16] +
                  mat_A[28][30] * mat_B[30][16] +
                  mat_A[28][31] * mat_B[31][16];
    mat_C[28][17] <= 
                  mat_A[28][0] * mat_B[0][17] +
                  mat_A[28][1] * mat_B[1][17] +
                  mat_A[28][2] * mat_B[2][17] +
                  mat_A[28][3] * mat_B[3][17] +
                  mat_A[28][4] * mat_B[4][17] +
                  mat_A[28][5] * mat_B[5][17] +
                  mat_A[28][6] * mat_B[6][17] +
                  mat_A[28][7] * mat_B[7][17] +
                  mat_A[28][8] * mat_B[8][17] +
                  mat_A[28][9] * mat_B[9][17] +
                  mat_A[28][10] * mat_B[10][17] +
                  mat_A[28][11] * mat_B[11][17] +
                  mat_A[28][12] * mat_B[12][17] +
                  mat_A[28][13] * mat_B[13][17] +
                  mat_A[28][14] * mat_B[14][17] +
                  mat_A[28][15] * mat_B[15][17] +
                  mat_A[28][16] * mat_B[16][17] +
                  mat_A[28][17] * mat_B[17][17] +
                  mat_A[28][18] * mat_B[18][17] +
                  mat_A[28][19] * mat_B[19][17] +
                  mat_A[28][20] * mat_B[20][17] +
                  mat_A[28][21] * mat_B[21][17] +
                  mat_A[28][22] * mat_B[22][17] +
                  mat_A[28][23] * mat_B[23][17] +
                  mat_A[28][24] * mat_B[24][17] +
                  mat_A[28][25] * mat_B[25][17] +
                  mat_A[28][26] * mat_B[26][17] +
                  mat_A[28][27] * mat_B[27][17] +
                  mat_A[28][28] * mat_B[28][17] +
                  mat_A[28][29] * mat_B[29][17] +
                  mat_A[28][30] * mat_B[30][17] +
                  mat_A[28][31] * mat_B[31][17];
    mat_C[28][18] <= 
                  mat_A[28][0] * mat_B[0][18] +
                  mat_A[28][1] * mat_B[1][18] +
                  mat_A[28][2] * mat_B[2][18] +
                  mat_A[28][3] * mat_B[3][18] +
                  mat_A[28][4] * mat_B[4][18] +
                  mat_A[28][5] * mat_B[5][18] +
                  mat_A[28][6] * mat_B[6][18] +
                  mat_A[28][7] * mat_B[7][18] +
                  mat_A[28][8] * mat_B[8][18] +
                  mat_A[28][9] * mat_B[9][18] +
                  mat_A[28][10] * mat_B[10][18] +
                  mat_A[28][11] * mat_B[11][18] +
                  mat_A[28][12] * mat_B[12][18] +
                  mat_A[28][13] * mat_B[13][18] +
                  mat_A[28][14] * mat_B[14][18] +
                  mat_A[28][15] * mat_B[15][18] +
                  mat_A[28][16] * mat_B[16][18] +
                  mat_A[28][17] * mat_B[17][18] +
                  mat_A[28][18] * mat_B[18][18] +
                  mat_A[28][19] * mat_B[19][18] +
                  mat_A[28][20] * mat_B[20][18] +
                  mat_A[28][21] * mat_B[21][18] +
                  mat_A[28][22] * mat_B[22][18] +
                  mat_A[28][23] * mat_B[23][18] +
                  mat_A[28][24] * mat_B[24][18] +
                  mat_A[28][25] * mat_B[25][18] +
                  mat_A[28][26] * mat_B[26][18] +
                  mat_A[28][27] * mat_B[27][18] +
                  mat_A[28][28] * mat_B[28][18] +
                  mat_A[28][29] * mat_B[29][18] +
                  mat_A[28][30] * mat_B[30][18] +
                  mat_A[28][31] * mat_B[31][18];
    mat_C[28][19] <= 
                  mat_A[28][0] * mat_B[0][19] +
                  mat_A[28][1] * mat_B[1][19] +
                  mat_A[28][2] * mat_B[2][19] +
                  mat_A[28][3] * mat_B[3][19] +
                  mat_A[28][4] * mat_B[4][19] +
                  mat_A[28][5] * mat_B[5][19] +
                  mat_A[28][6] * mat_B[6][19] +
                  mat_A[28][7] * mat_B[7][19] +
                  mat_A[28][8] * mat_B[8][19] +
                  mat_A[28][9] * mat_B[9][19] +
                  mat_A[28][10] * mat_B[10][19] +
                  mat_A[28][11] * mat_B[11][19] +
                  mat_A[28][12] * mat_B[12][19] +
                  mat_A[28][13] * mat_B[13][19] +
                  mat_A[28][14] * mat_B[14][19] +
                  mat_A[28][15] * mat_B[15][19] +
                  mat_A[28][16] * mat_B[16][19] +
                  mat_A[28][17] * mat_B[17][19] +
                  mat_A[28][18] * mat_B[18][19] +
                  mat_A[28][19] * mat_B[19][19] +
                  mat_A[28][20] * mat_B[20][19] +
                  mat_A[28][21] * mat_B[21][19] +
                  mat_A[28][22] * mat_B[22][19] +
                  mat_A[28][23] * mat_B[23][19] +
                  mat_A[28][24] * mat_B[24][19] +
                  mat_A[28][25] * mat_B[25][19] +
                  mat_A[28][26] * mat_B[26][19] +
                  mat_A[28][27] * mat_B[27][19] +
                  mat_A[28][28] * mat_B[28][19] +
                  mat_A[28][29] * mat_B[29][19] +
                  mat_A[28][30] * mat_B[30][19] +
                  mat_A[28][31] * mat_B[31][19];
    mat_C[28][20] <= 
                  mat_A[28][0] * mat_B[0][20] +
                  mat_A[28][1] * mat_B[1][20] +
                  mat_A[28][2] * mat_B[2][20] +
                  mat_A[28][3] * mat_B[3][20] +
                  mat_A[28][4] * mat_B[4][20] +
                  mat_A[28][5] * mat_B[5][20] +
                  mat_A[28][6] * mat_B[6][20] +
                  mat_A[28][7] * mat_B[7][20] +
                  mat_A[28][8] * mat_B[8][20] +
                  mat_A[28][9] * mat_B[9][20] +
                  mat_A[28][10] * mat_B[10][20] +
                  mat_A[28][11] * mat_B[11][20] +
                  mat_A[28][12] * mat_B[12][20] +
                  mat_A[28][13] * mat_B[13][20] +
                  mat_A[28][14] * mat_B[14][20] +
                  mat_A[28][15] * mat_B[15][20] +
                  mat_A[28][16] * mat_B[16][20] +
                  mat_A[28][17] * mat_B[17][20] +
                  mat_A[28][18] * mat_B[18][20] +
                  mat_A[28][19] * mat_B[19][20] +
                  mat_A[28][20] * mat_B[20][20] +
                  mat_A[28][21] * mat_B[21][20] +
                  mat_A[28][22] * mat_B[22][20] +
                  mat_A[28][23] * mat_B[23][20] +
                  mat_A[28][24] * mat_B[24][20] +
                  mat_A[28][25] * mat_B[25][20] +
                  mat_A[28][26] * mat_B[26][20] +
                  mat_A[28][27] * mat_B[27][20] +
                  mat_A[28][28] * mat_B[28][20] +
                  mat_A[28][29] * mat_B[29][20] +
                  mat_A[28][30] * mat_B[30][20] +
                  mat_A[28][31] * mat_B[31][20];
    mat_C[28][21] <= 
                  mat_A[28][0] * mat_B[0][21] +
                  mat_A[28][1] * mat_B[1][21] +
                  mat_A[28][2] * mat_B[2][21] +
                  mat_A[28][3] * mat_B[3][21] +
                  mat_A[28][4] * mat_B[4][21] +
                  mat_A[28][5] * mat_B[5][21] +
                  mat_A[28][6] * mat_B[6][21] +
                  mat_A[28][7] * mat_B[7][21] +
                  mat_A[28][8] * mat_B[8][21] +
                  mat_A[28][9] * mat_B[9][21] +
                  mat_A[28][10] * mat_B[10][21] +
                  mat_A[28][11] * mat_B[11][21] +
                  mat_A[28][12] * mat_B[12][21] +
                  mat_A[28][13] * mat_B[13][21] +
                  mat_A[28][14] * mat_B[14][21] +
                  mat_A[28][15] * mat_B[15][21] +
                  mat_A[28][16] * mat_B[16][21] +
                  mat_A[28][17] * mat_B[17][21] +
                  mat_A[28][18] * mat_B[18][21] +
                  mat_A[28][19] * mat_B[19][21] +
                  mat_A[28][20] * mat_B[20][21] +
                  mat_A[28][21] * mat_B[21][21] +
                  mat_A[28][22] * mat_B[22][21] +
                  mat_A[28][23] * mat_B[23][21] +
                  mat_A[28][24] * mat_B[24][21] +
                  mat_A[28][25] * mat_B[25][21] +
                  mat_A[28][26] * mat_B[26][21] +
                  mat_A[28][27] * mat_B[27][21] +
                  mat_A[28][28] * mat_B[28][21] +
                  mat_A[28][29] * mat_B[29][21] +
                  mat_A[28][30] * mat_B[30][21] +
                  mat_A[28][31] * mat_B[31][21];
    mat_C[28][22] <= 
                  mat_A[28][0] * mat_B[0][22] +
                  mat_A[28][1] * mat_B[1][22] +
                  mat_A[28][2] * mat_B[2][22] +
                  mat_A[28][3] * mat_B[3][22] +
                  mat_A[28][4] * mat_B[4][22] +
                  mat_A[28][5] * mat_B[5][22] +
                  mat_A[28][6] * mat_B[6][22] +
                  mat_A[28][7] * mat_B[7][22] +
                  mat_A[28][8] * mat_B[8][22] +
                  mat_A[28][9] * mat_B[9][22] +
                  mat_A[28][10] * mat_B[10][22] +
                  mat_A[28][11] * mat_B[11][22] +
                  mat_A[28][12] * mat_B[12][22] +
                  mat_A[28][13] * mat_B[13][22] +
                  mat_A[28][14] * mat_B[14][22] +
                  mat_A[28][15] * mat_B[15][22] +
                  mat_A[28][16] * mat_B[16][22] +
                  mat_A[28][17] * mat_B[17][22] +
                  mat_A[28][18] * mat_B[18][22] +
                  mat_A[28][19] * mat_B[19][22] +
                  mat_A[28][20] * mat_B[20][22] +
                  mat_A[28][21] * mat_B[21][22] +
                  mat_A[28][22] * mat_B[22][22] +
                  mat_A[28][23] * mat_B[23][22] +
                  mat_A[28][24] * mat_B[24][22] +
                  mat_A[28][25] * mat_B[25][22] +
                  mat_A[28][26] * mat_B[26][22] +
                  mat_A[28][27] * mat_B[27][22] +
                  mat_A[28][28] * mat_B[28][22] +
                  mat_A[28][29] * mat_B[29][22] +
                  mat_A[28][30] * mat_B[30][22] +
                  mat_A[28][31] * mat_B[31][22];
    mat_C[28][23] <= 
                  mat_A[28][0] * mat_B[0][23] +
                  mat_A[28][1] * mat_B[1][23] +
                  mat_A[28][2] * mat_B[2][23] +
                  mat_A[28][3] * mat_B[3][23] +
                  mat_A[28][4] * mat_B[4][23] +
                  mat_A[28][5] * mat_B[5][23] +
                  mat_A[28][6] * mat_B[6][23] +
                  mat_A[28][7] * mat_B[7][23] +
                  mat_A[28][8] * mat_B[8][23] +
                  mat_A[28][9] * mat_B[9][23] +
                  mat_A[28][10] * mat_B[10][23] +
                  mat_A[28][11] * mat_B[11][23] +
                  mat_A[28][12] * mat_B[12][23] +
                  mat_A[28][13] * mat_B[13][23] +
                  mat_A[28][14] * mat_B[14][23] +
                  mat_A[28][15] * mat_B[15][23] +
                  mat_A[28][16] * mat_B[16][23] +
                  mat_A[28][17] * mat_B[17][23] +
                  mat_A[28][18] * mat_B[18][23] +
                  mat_A[28][19] * mat_B[19][23] +
                  mat_A[28][20] * mat_B[20][23] +
                  mat_A[28][21] * mat_B[21][23] +
                  mat_A[28][22] * mat_B[22][23] +
                  mat_A[28][23] * mat_B[23][23] +
                  mat_A[28][24] * mat_B[24][23] +
                  mat_A[28][25] * mat_B[25][23] +
                  mat_A[28][26] * mat_B[26][23] +
                  mat_A[28][27] * mat_B[27][23] +
                  mat_A[28][28] * mat_B[28][23] +
                  mat_A[28][29] * mat_B[29][23] +
                  mat_A[28][30] * mat_B[30][23] +
                  mat_A[28][31] * mat_B[31][23];
    mat_C[28][24] <= 
                  mat_A[28][0] * mat_B[0][24] +
                  mat_A[28][1] * mat_B[1][24] +
                  mat_A[28][2] * mat_B[2][24] +
                  mat_A[28][3] * mat_B[3][24] +
                  mat_A[28][4] * mat_B[4][24] +
                  mat_A[28][5] * mat_B[5][24] +
                  mat_A[28][6] * mat_B[6][24] +
                  mat_A[28][7] * mat_B[7][24] +
                  mat_A[28][8] * mat_B[8][24] +
                  mat_A[28][9] * mat_B[9][24] +
                  mat_A[28][10] * mat_B[10][24] +
                  mat_A[28][11] * mat_B[11][24] +
                  mat_A[28][12] * mat_B[12][24] +
                  mat_A[28][13] * mat_B[13][24] +
                  mat_A[28][14] * mat_B[14][24] +
                  mat_A[28][15] * mat_B[15][24] +
                  mat_A[28][16] * mat_B[16][24] +
                  mat_A[28][17] * mat_B[17][24] +
                  mat_A[28][18] * mat_B[18][24] +
                  mat_A[28][19] * mat_B[19][24] +
                  mat_A[28][20] * mat_B[20][24] +
                  mat_A[28][21] * mat_B[21][24] +
                  mat_A[28][22] * mat_B[22][24] +
                  mat_A[28][23] * mat_B[23][24] +
                  mat_A[28][24] * mat_B[24][24] +
                  mat_A[28][25] * mat_B[25][24] +
                  mat_A[28][26] * mat_B[26][24] +
                  mat_A[28][27] * mat_B[27][24] +
                  mat_A[28][28] * mat_B[28][24] +
                  mat_A[28][29] * mat_B[29][24] +
                  mat_A[28][30] * mat_B[30][24] +
                  mat_A[28][31] * mat_B[31][24];
    mat_C[28][25] <= 
                  mat_A[28][0] * mat_B[0][25] +
                  mat_A[28][1] * mat_B[1][25] +
                  mat_A[28][2] * mat_B[2][25] +
                  mat_A[28][3] * mat_B[3][25] +
                  mat_A[28][4] * mat_B[4][25] +
                  mat_A[28][5] * mat_B[5][25] +
                  mat_A[28][6] * mat_B[6][25] +
                  mat_A[28][7] * mat_B[7][25] +
                  mat_A[28][8] * mat_B[8][25] +
                  mat_A[28][9] * mat_B[9][25] +
                  mat_A[28][10] * mat_B[10][25] +
                  mat_A[28][11] * mat_B[11][25] +
                  mat_A[28][12] * mat_B[12][25] +
                  mat_A[28][13] * mat_B[13][25] +
                  mat_A[28][14] * mat_B[14][25] +
                  mat_A[28][15] * mat_B[15][25] +
                  mat_A[28][16] * mat_B[16][25] +
                  mat_A[28][17] * mat_B[17][25] +
                  mat_A[28][18] * mat_B[18][25] +
                  mat_A[28][19] * mat_B[19][25] +
                  mat_A[28][20] * mat_B[20][25] +
                  mat_A[28][21] * mat_B[21][25] +
                  mat_A[28][22] * mat_B[22][25] +
                  mat_A[28][23] * mat_B[23][25] +
                  mat_A[28][24] * mat_B[24][25] +
                  mat_A[28][25] * mat_B[25][25] +
                  mat_A[28][26] * mat_B[26][25] +
                  mat_A[28][27] * mat_B[27][25] +
                  mat_A[28][28] * mat_B[28][25] +
                  mat_A[28][29] * mat_B[29][25] +
                  mat_A[28][30] * mat_B[30][25] +
                  mat_A[28][31] * mat_B[31][25];
    mat_C[28][26] <= 
                  mat_A[28][0] * mat_B[0][26] +
                  mat_A[28][1] * mat_B[1][26] +
                  mat_A[28][2] * mat_B[2][26] +
                  mat_A[28][3] * mat_B[3][26] +
                  mat_A[28][4] * mat_B[4][26] +
                  mat_A[28][5] * mat_B[5][26] +
                  mat_A[28][6] * mat_B[6][26] +
                  mat_A[28][7] * mat_B[7][26] +
                  mat_A[28][8] * mat_B[8][26] +
                  mat_A[28][9] * mat_B[9][26] +
                  mat_A[28][10] * mat_B[10][26] +
                  mat_A[28][11] * mat_B[11][26] +
                  mat_A[28][12] * mat_B[12][26] +
                  mat_A[28][13] * mat_B[13][26] +
                  mat_A[28][14] * mat_B[14][26] +
                  mat_A[28][15] * mat_B[15][26] +
                  mat_A[28][16] * mat_B[16][26] +
                  mat_A[28][17] * mat_B[17][26] +
                  mat_A[28][18] * mat_B[18][26] +
                  mat_A[28][19] * mat_B[19][26] +
                  mat_A[28][20] * mat_B[20][26] +
                  mat_A[28][21] * mat_B[21][26] +
                  mat_A[28][22] * mat_B[22][26] +
                  mat_A[28][23] * mat_B[23][26] +
                  mat_A[28][24] * mat_B[24][26] +
                  mat_A[28][25] * mat_B[25][26] +
                  mat_A[28][26] * mat_B[26][26] +
                  mat_A[28][27] * mat_B[27][26] +
                  mat_A[28][28] * mat_B[28][26] +
                  mat_A[28][29] * mat_B[29][26] +
                  mat_A[28][30] * mat_B[30][26] +
                  mat_A[28][31] * mat_B[31][26];
    mat_C[28][27] <= 
                  mat_A[28][0] * mat_B[0][27] +
                  mat_A[28][1] * mat_B[1][27] +
                  mat_A[28][2] * mat_B[2][27] +
                  mat_A[28][3] * mat_B[3][27] +
                  mat_A[28][4] * mat_B[4][27] +
                  mat_A[28][5] * mat_B[5][27] +
                  mat_A[28][6] * mat_B[6][27] +
                  mat_A[28][7] * mat_B[7][27] +
                  mat_A[28][8] * mat_B[8][27] +
                  mat_A[28][9] * mat_B[9][27] +
                  mat_A[28][10] * mat_B[10][27] +
                  mat_A[28][11] * mat_B[11][27] +
                  mat_A[28][12] * mat_B[12][27] +
                  mat_A[28][13] * mat_B[13][27] +
                  mat_A[28][14] * mat_B[14][27] +
                  mat_A[28][15] * mat_B[15][27] +
                  mat_A[28][16] * mat_B[16][27] +
                  mat_A[28][17] * mat_B[17][27] +
                  mat_A[28][18] * mat_B[18][27] +
                  mat_A[28][19] * mat_B[19][27] +
                  mat_A[28][20] * mat_B[20][27] +
                  mat_A[28][21] * mat_B[21][27] +
                  mat_A[28][22] * mat_B[22][27] +
                  mat_A[28][23] * mat_B[23][27] +
                  mat_A[28][24] * mat_B[24][27] +
                  mat_A[28][25] * mat_B[25][27] +
                  mat_A[28][26] * mat_B[26][27] +
                  mat_A[28][27] * mat_B[27][27] +
                  mat_A[28][28] * mat_B[28][27] +
                  mat_A[28][29] * mat_B[29][27] +
                  mat_A[28][30] * mat_B[30][27] +
                  mat_A[28][31] * mat_B[31][27];
    mat_C[28][28] <= 
                  mat_A[28][0] * mat_B[0][28] +
                  mat_A[28][1] * mat_B[1][28] +
                  mat_A[28][2] * mat_B[2][28] +
                  mat_A[28][3] * mat_B[3][28] +
                  mat_A[28][4] * mat_B[4][28] +
                  mat_A[28][5] * mat_B[5][28] +
                  mat_A[28][6] * mat_B[6][28] +
                  mat_A[28][7] * mat_B[7][28] +
                  mat_A[28][8] * mat_B[8][28] +
                  mat_A[28][9] * mat_B[9][28] +
                  mat_A[28][10] * mat_B[10][28] +
                  mat_A[28][11] * mat_B[11][28] +
                  mat_A[28][12] * mat_B[12][28] +
                  mat_A[28][13] * mat_B[13][28] +
                  mat_A[28][14] * mat_B[14][28] +
                  mat_A[28][15] * mat_B[15][28] +
                  mat_A[28][16] * mat_B[16][28] +
                  mat_A[28][17] * mat_B[17][28] +
                  mat_A[28][18] * mat_B[18][28] +
                  mat_A[28][19] * mat_B[19][28] +
                  mat_A[28][20] * mat_B[20][28] +
                  mat_A[28][21] * mat_B[21][28] +
                  mat_A[28][22] * mat_B[22][28] +
                  mat_A[28][23] * mat_B[23][28] +
                  mat_A[28][24] * mat_B[24][28] +
                  mat_A[28][25] * mat_B[25][28] +
                  mat_A[28][26] * mat_B[26][28] +
                  mat_A[28][27] * mat_B[27][28] +
                  mat_A[28][28] * mat_B[28][28] +
                  mat_A[28][29] * mat_B[29][28] +
                  mat_A[28][30] * mat_B[30][28] +
                  mat_A[28][31] * mat_B[31][28];
    mat_C[28][29] <= 
                  mat_A[28][0] * mat_B[0][29] +
                  mat_A[28][1] * mat_B[1][29] +
                  mat_A[28][2] * mat_B[2][29] +
                  mat_A[28][3] * mat_B[3][29] +
                  mat_A[28][4] * mat_B[4][29] +
                  mat_A[28][5] * mat_B[5][29] +
                  mat_A[28][6] * mat_B[6][29] +
                  mat_A[28][7] * mat_B[7][29] +
                  mat_A[28][8] * mat_B[8][29] +
                  mat_A[28][9] * mat_B[9][29] +
                  mat_A[28][10] * mat_B[10][29] +
                  mat_A[28][11] * mat_B[11][29] +
                  mat_A[28][12] * mat_B[12][29] +
                  mat_A[28][13] * mat_B[13][29] +
                  mat_A[28][14] * mat_B[14][29] +
                  mat_A[28][15] * mat_B[15][29] +
                  mat_A[28][16] * mat_B[16][29] +
                  mat_A[28][17] * mat_B[17][29] +
                  mat_A[28][18] * mat_B[18][29] +
                  mat_A[28][19] * mat_B[19][29] +
                  mat_A[28][20] * mat_B[20][29] +
                  mat_A[28][21] * mat_B[21][29] +
                  mat_A[28][22] * mat_B[22][29] +
                  mat_A[28][23] * mat_B[23][29] +
                  mat_A[28][24] * mat_B[24][29] +
                  mat_A[28][25] * mat_B[25][29] +
                  mat_A[28][26] * mat_B[26][29] +
                  mat_A[28][27] * mat_B[27][29] +
                  mat_A[28][28] * mat_B[28][29] +
                  mat_A[28][29] * mat_B[29][29] +
                  mat_A[28][30] * mat_B[30][29] +
                  mat_A[28][31] * mat_B[31][29];
    mat_C[28][30] <= 
                  mat_A[28][0] * mat_B[0][30] +
                  mat_A[28][1] * mat_B[1][30] +
                  mat_A[28][2] * mat_B[2][30] +
                  mat_A[28][3] * mat_B[3][30] +
                  mat_A[28][4] * mat_B[4][30] +
                  mat_A[28][5] * mat_B[5][30] +
                  mat_A[28][6] * mat_B[6][30] +
                  mat_A[28][7] * mat_B[7][30] +
                  mat_A[28][8] * mat_B[8][30] +
                  mat_A[28][9] * mat_B[9][30] +
                  mat_A[28][10] * mat_B[10][30] +
                  mat_A[28][11] * mat_B[11][30] +
                  mat_A[28][12] * mat_B[12][30] +
                  mat_A[28][13] * mat_B[13][30] +
                  mat_A[28][14] * mat_B[14][30] +
                  mat_A[28][15] * mat_B[15][30] +
                  mat_A[28][16] * mat_B[16][30] +
                  mat_A[28][17] * mat_B[17][30] +
                  mat_A[28][18] * mat_B[18][30] +
                  mat_A[28][19] * mat_B[19][30] +
                  mat_A[28][20] * mat_B[20][30] +
                  mat_A[28][21] * mat_B[21][30] +
                  mat_A[28][22] * mat_B[22][30] +
                  mat_A[28][23] * mat_B[23][30] +
                  mat_A[28][24] * mat_B[24][30] +
                  mat_A[28][25] * mat_B[25][30] +
                  mat_A[28][26] * mat_B[26][30] +
                  mat_A[28][27] * mat_B[27][30] +
                  mat_A[28][28] * mat_B[28][30] +
                  mat_A[28][29] * mat_B[29][30] +
                  mat_A[28][30] * mat_B[30][30] +
                  mat_A[28][31] * mat_B[31][30];
    mat_C[28][31] <= 
                  mat_A[28][0] * mat_B[0][31] +
                  mat_A[28][1] * mat_B[1][31] +
                  mat_A[28][2] * mat_B[2][31] +
                  mat_A[28][3] * mat_B[3][31] +
                  mat_A[28][4] * mat_B[4][31] +
                  mat_A[28][5] * mat_B[5][31] +
                  mat_A[28][6] * mat_B[6][31] +
                  mat_A[28][7] * mat_B[7][31] +
                  mat_A[28][8] * mat_B[8][31] +
                  mat_A[28][9] * mat_B[9][31] +
                  mat_A[28][10] * mat_B[10][31] +
                  mat_A[28][11] * mat_B[11][31] +
                  mat_A[28][12] * mat_B[12][31] +
                  mat_A[28][13] * mat_B[13][31] +
                  mat_A[28][14] * mat_B[14][31] +
                  mat_A[28][15] * mat_B[15][31] +
                  mat_A[28][16] * mat_B[16][31] +
                  mat_A[28][17] * mat_B[17][31] +
                  mat_A[28][18] * mat_B[18][31] +
                  mat_A[28][19] * mat_B[19][31] +
                  mat_A[28][20] * mat_B[20][31] +
                  mat_A[28][21] * mat_B[21][31] +
                  mat_A[28][22] * mat_B[22][31] +
                  mat_A[28][23] * mat_B[23][31] +
                  mat_A[28][24] * mat_B[24][31] +
                  mat_A[28][25] * mat_B[25][31] +
                  mat_A[28][26] * mat_B[26][31] +
                  mat_A[28][27] * mat_B[27][31] +
                  mat_A[28][28] * mat_B[28][31] +
                  mat_A[28][29] * mat_B[29][31] +
                  mat_A[28][30] * mat_B[30][31] +
                  mat_A[28][31] * mat_B[31][31];
    mat_C[29][0] <= 
                  mat_A[29][0] * mat_B[0][0] +
                  mat_A[29][1] * mat_B[1][0] +
                  mat_A[29][2] * mat_B[2][0] +
                  mat_A[29][3] * mat_B[3][0] +
                  mat_A[29][4] * mat_B[4][0] +
                  mat_A[29][5] * mat_B[5][0] +
                  mat_A[29][6] * mat_B[6][0] +
                  mat_A[29][7] * mat_B[7][0] +
                  mat_A[29][8] * mat_B[8][0] +
                  mat_A[29][9] * mat_B[9][0] +
                  mat_A[29][10] * mat_B[10][0] +
                  mat_A[29][11] * mat_B[11][0] +
                  mat_A[29][12] * mat_B[12][0] +
                  mat_A[29][13] * mat_B[13][0] +
                  mat_A[29][14] * mat_B[14][0] +
                  mat_A[29][15] * mat_B[15][0] +
                  mat_A[29][16] * mat_B[16][0] +
                  mat_A[29][17] * mat_B[17][0] +
                  mat_A[29][18] * mat_B[18][0] +
                  mat_A[29][19] * mat_B[19][0] +
                  mat_A[29][20] * mat_B[20][0] +
                  mat_A[29][21] * mat_B[21][0] +
                  mat_A[29][22] * mat_B[22][0] +
                  mat_A[29][23] * mat_B[23][0] +
                  mat_A[29][24] * mat_B[24][0] +
                  mat_A[29][25] * mat_B[25][0] +
                  mat_A[29][26] * mat_B[26][0] +
                  mat_A[29][27] * mat_B[27][0] +
                  mat_A[29][28] * mat_B[28][0] +
                  mat_A[29][29] * mat_B[29][0] +
                  mat_A[29][30] * mat_B[30][0] +
                  mat_A[29][31] * mat_B[31][0];
    mat_C[29][1] <= 
                  mat_A[29][0] * mat_B[0][1] +
                  mat_A[29][1] * mat_B[1][1] +
                  mat_A[29][2] * mat_B[2][1] +
                  mat_A[29][3] * mat_B[3][1] +
                  mat_A[29][4] * mat_B[4][1] +
                  mat_A[29][5] * mat_B[5][1] +
                  mat_A[29][6] * mat_B[6][1] +
                  mat_A[29][7] * mat_B[7][1] +
                  mat_A[29][8] * mat_B[8][1] +
                  mat_A[29][9] * mat_B[9][1] +
                  mat_A[29][10] * mat_B[10][1] +
                  mat_A[29][11] * mat_B[11][1] +
                  mat_A[29][12] * mat_B[12][1] +
                  mat_A[29][13] * mat_B[13][1] +
                  mat_A[29][14] * mat_B[14][1] +
                  mat_A[29][15] * mat_B[15][1] +
                  mat_A[29][16] * mat_B[16][1] +
                  mat_A[29][17] * mat_B[17][1] +
                  mat_A[29][18] * mat_B[18][1] +
                  mat_A[29][19] * mat_B[19][1] +
                  mat_A[29][20] * mat_B[20][1] +
                  mat_A[29][21] * mat_B[21][1] +
                  mat_A[29][22] * mat_B[22][1] +
                  mat_A[29][23] * mat_B[23][1] +
                  mat_A[29][24] * mat_B[24][1] +
                  mat_A[29][25] * mat_B[25][1] +
                  mat_A[29][26] * mat_B[26][1] +
                  mat_A[29][27] * mat_B[27][1] +
                  mat_A[29][28] * mat_B[28][1] +
                  mat_A[29][29] * mat_B[29][1] +
                  mat_A[29][30] * mat_B[30][1] +
                  mat_A[29][31] * mat_B[31][1];
    mat_C[29][2] <= 
                  mat_A[29][0] * mat_B[0][2] +
                  mat_A[29][1] * mat_B[1][2] +
                  mat_A[29][2] * mat_B[2][2] +
                  mat_A[29][3] * mat_B[3][2] +
                  mat_A[29][4] * mat_B[4][2] +
                  mat_A[29][5] * mat_B[5][2] +
                  mat_A[29][6] * mat_B[6][2] +
                  mat_A[29][7] * mat_B[7][2] +
                  mat_A[29][8] * mat_B[8][2] +
                  mat_A[29][9] * mat_B[9][2] +
                  mat_A[29][10] * mat_B[10][2] +
                  mat_A[29][11] * mat_B[11][2] +
                  mat_A[29][12] * mat_B[12][2] +
                  mat_A[29][13] * mat_B[13][2] +
                  mat_A[29][14] * mat_B[14][2] +
                  mat_A[29][15] * mat_B[15][2] +
                  mat_A[29][16] * mat_B[16][2] +
                  mat_A[29][17] * mat_B[17][2] +
                  mat_A[29][18] * mat_B[18][2] +
                  mat_A[29][19] * mat_B[19][2] +
                  mat_A[29][20] * mat_B[20][2] +
                  mat_A[29][21] * mat_B[21][2] +
                  mat_A[29][22] * mat_B[22][2] +
                  mat_A[29][23] * mat_B[23][2] +
                  mat_A[29][24] * mat_B[24][2] +
                  mat_A[29][25] * mat_B[25][2] +
                  mat_A[29][26] * mat_B[26][2] +
                  mat_A[29][27] * mat_B[27][2] +
                  mat_A[29][28] * mat_B[28][2] +
                  mat_A[29][29] * mat_B[29][2] +
                  mat_A[29][30] * mat_B[30][2] +
                  mat_A[29][31] * mat_B[31][2];
    mat_C[29][3] <= 
                  mat_A[29][0] * mat_B[0][3] +
                  mat_A[29][1] * mat_B[1][3] +
                  mat_A[29][2] * mat_B[2][3] +
                  mat_A[29][3] * mat_B[3][3] +
                  mat_A[29][4] * mat_B[4][3] +
                  mat_A[29][5] * mat_B[5][3] +
                  mat_A[29][6] * mat_B[6][3] +
                  mat_A[29][7] * mat_B[7][3] +
                  mat_A[29][8] * mat_B[8][3] +
                  mat_A[29][9] * mat_B[9][3] +
                  mat_A[29][10] * mat_B[10][3] +
                  mat_A[29][11] * mat_B[11][3] +
                  mat_A[29][12] * mat_B[12][3] +
                  mat_A[29][13] * mat_B[13][3] +
                  mat_A[29][14] * mat_B[14][3] +
                  mat_A[29][15] * mat_B[15][3] +
                  mat_A[29][16] * mat_B[16][3] +
                  mat_A[29][17] * mat_B[17][3] +
                  mat_A[29][18] * mat_B[18][3] +
                  mat_A[29][19] * mat_B[19][3] +
                  mat_A[29][20] * mat_B[20][3] +
                  mat_A[29][21] * mat_B[21][3] +
                  mat_A[29][22] * mat_B[22][3] +
                  mat_A[29][23] * mat_B[23][3] +
                  mat_A[29][24] * mat_B[24][3] +
                  mat_A[29][25] * mat_B[25][3] +
                  mat_A[29][26] * mat_B[26][3] +
                  mat_A[29][27] * mat_B[27][3] +
                  mat_A[29][28] * mat_B[28][3] +
                  mat_A[29][29] * mat_B[29][3] +
                  mat_A[29][30] * mat_B[30][3] +
                  mat_A[29][31] * mat_B[31][3];
    mat_C[29][4] <= 
                  mat_A[29][0] * mat_B[0][4] +
                  mat_A[29][1] * mat_B[1][4] +
                  mat_A[29][2] * mat_B[2][4] +
                  mat_A[29][3] * mat_B[3][4] +
                  mat_A[29][4] * mat_B[4][4] +
                  mat_A[29][5] * mat_B[5][4] +
                  mat_A[29][6] * mat_B[6][4] +
                  mat_A[29][7] * mat_B[7][4] +
                  mat_A[29][8] * mat_B[8][4] +
                  mat_A[29][9] * mat_B[9][4] +
                  mat_A[29][10] * mat_B[10][4] +
                  mat_A[29][11] * mat_B[11][4] +
                  mat_A[29][12] * mat_B[12][4] +
                  mat_A[29][13] * mat_B[13][4] +
                  mat_A[29][14] * mat_B[14][4] +
                  mat_A[29][15] * mat_B[15][4] +
                  mat_A[29][16] * mat_B[16][4] +
                  mat_A[29][17] * mat_B[17][4] +
                  mat_A[29][18] * mat_B[18][4] +
                  mat_A[29][19] * mat_B[19][4] +
                  mat_A[29][20] * mat_B[20][4] +
                  mat_A[29][21] * mat_B[21][4] +
                  mat_A[29][22] * mat_B[22][4] +
                  mat_A[29][23] * mat_B[23][4] +
                  mat_A[29][24] * mat_B[24][4] +
                  mat_A[29][25] * mat_B[25][4] +
                  mat_A[29][26] * mat_B[26][4] +
                  mat_A[29][27] * mat_B[27][4] +
                  mat_A[29][28] * mat_B[28][4] +
                  mat_A[29][29] * mat_B[29][4] +
                  mat_A[29][30] * mat_B[30][4] +
                  mat_A[29][31] * mat_B[31][4];
    mat_C[29][5] <= 
                  mat_A[29][0] * mat_B[0][5] +
                  mat_A[29][1] * mat_B[1][5] +
                  mat_A[29][2] * mat_B[2][5] +
                  mat_A[29][3] * mat_B[3][5] +
                  mat_A[29][4] * mat_B[4][5] +
                  mat_A[29][5] * mat_B[5][5] +
                  mat_A[29][6] * mat_B[6][5] +
                  mat_A[29][7] * mat_B[7][5] +
                  mat_A[29][8] * mat_B[8][5] +
                  mat_A[29][9] * mat_B[9][5] +
                  mat_A[29][10] * mat_B[10][5] +
                  mat_A[29][11] * mat_B[11][5] +
                  mat_A[29][12] * mat_B[12][5] +
                  mat_A[29][13] * mat_B[13][5] +
                  mat_A[29][14] * mat_B[14][5] +
                  mat_A[29][15] * mat_B[15][5] +
                  mat_A[29][16] * mat_B[16][5] +
                  mat_A[29][17] * mat_B[17][5] +
                  mat_A[29][18] * mat_B[18][5] +
                  mat_A[29][19] * mat_B[19][5] +
                  mat_A[29][20] * mat_B[20][5] +
                  mat_A[29][21] * mat_B[21][5] +
                  mat_A[29][22] * mat_B[22][5] +
                  mat_A[29][23] * mat_B[23][5] +
                  mat_A[29][24] * mat_B[24][5] +
                  mat_A[29][25] * mat_B[25][5] +
                  mat_A[29][26] * mat_B[26][5] +
                  mat_A[29][27] * mat_B[27][5] +
                  mat_A[29][28] * mat_B[28][5] +
                  mat_A[29][29] * mat_B[29][5] +
                  mat_A[29][30] * mat_B[30][5] +
                  mat_A[29][31] * mat_B[31][5];
    mat_C[29][6] <= 
                  mat_A[29][0] * mat_B[0][6] +
                  mat_A[29][1] * mat_B[1][6] +
                  mat_A[29][2] * mat_B[2][6] +
                  mat_A[29][3] * mat_B[3][6] +
                  mat_A[29][4] * mat_B[4][6] +
                  mat_A[29][5] * mat_B[5][6] +
                  mat_A[29][6] * mat_B[6][6] +
                  mat_A[29][7] * mat_B[7][6] +
                  mat_A[29][8] * mat_B[8][6] +
                  mat_A[29][9] * mat_B[9][6] +
                  mat_A[29][10] * mat_B[10][6] +
                  mat_A[29][11] * mat_B[11][6] +
                  mat_A[29][12] * mat_B[12][6] +
                  mat_A[29][13] * mat_B[13][6] +
                  mat_A[29][14] * mat_B[14][6] +
                  mat_A[29][15] * mat_B[15][6] +
                  mat_A[29][16] * mat_B[16][6] +
                  mat_A[29][17] * mat_B[17][6] +
                  mat_A[29][18] * mat_B[18][6] +
                  mat_A[29][19] * mat_B[19][6] +
                  mat_A[29][20] * mat_B[20][6] +
                  mat_A[29][21] * mat_B[21][6] +
                  mat_A[29][22] * mat_B[22][6] +
                  mat_A[29][23] * mat_B[23][6] +
                  mat_A[29][24] * mat_B[24][6] +
                  mat_A[29][25] * mat_B[25][6] +
                  mat_A[29][26] * mat_B[26][6] +
                  mat_A[29][27] * mat_B[27][6] +
                  mat_A[29][28] * mat_B[28][6] +
                  mat_A[29][29] * mat_B[29][6] +
                  mat_A[29][30] * mat_B[30][6] +
                  mat_A[29][31] * mat_B[31][6];
    mat_C[29][7] <= 
                  mat_A[29][0] * mat_B[0][7] +
                  mat_A[29][1] * mat_B[1][7] +
                  mat_A[29][2] * mat_B[2][7] +
                  mat_A[29][3] * mat_B[3][7] +
                  mat_A[29][4] * mat_B[4][7] +
                  mat_A[29][5] * mat_B[5][7] +
                  mat_A[29][6] * mat_B[6][7] +
                  mat_A[29][7] * mat_B[7][7] +
                  mat_A[29][8] * mat_B[8][7] +
                  mat_A[29][9] * mat_B[9][7] +
                  mat_A[29][10] * mat_B[10][7] +
                  mat_A[29][11] * mat_B[11][7] +
                  mat_A[29][12] * mat_B[12][7] +
                  mat_A[29][13] * mat_B[13][7] +
                  mat_A[29][14] * mat_B[14][7] +
                  mat_A[29][15] * mat_B[15][7] +
                  mat_A[29][16] * mat_B[16][7] +
                  mat_A[29][17] * mat_B[17][7] +
                  mat_A[29][18] * mat_B[18][7] +
                  mat_A[29][19] * mat_B[19][7] +
                  mat_A[29][20] * mat_B[20][7] +
                  mat_A[29][21] * mat_B[21][7] +
                  mat_A[29][22] * mat_B[22][7] +
                  mat_A[29][23] * mat_B[23][7] +
                  mat_A[29][24] * mat_B[24][7] +
                  mat_A[29][25] * mat_B[25][7] +
                  mat_A[29][26] * mat_B[26][7] +
                  mat_A[29][27] * mat_B[27][7] +
                  mat_A[29][28] * mat_B[28][7] +
                  mat_A[29][29] * mat_B[29][7] +
                  mat_A[29][30] * mat_B[30][7] +
                  mat_A[29][31] * mat_B[31][7];
    mat_C[29][8] <= 
                  mat_A[29][0] * mat_B[0][8] +
                  mat_A[29][1] * mat_B[1][8] +
                  mat_A[29][2] * mat_B[2][8] +
                  mat_A[29][3] * mat_B[3][8] +
                  mat_A[29][4] * mat_B[4][8] +
                  mat_A[29][5] * mat_B[5][8] +
                  mat_A[29][6] * mat_B[6][8] +
                  mat_A[29][7] * mat_B[7][8] +
                  mat_A[29][8] * mat_B[8][8] +
                  mat_A[29][9] * mat_B[9][8] +
                  mat_A[29][10] * mat_B[10][8] +
                  mat_A[29][11] * mat_B[11][8] +
                  mat_A[29][12] * mat_B[12][8] +
                  mat_A[29][13] * mat_B[13][8] +
                  mat_A[29][14] * mat_B[14][8] +
                  mat_A[29][15] * mat_B[15][8] +
                  mat_A[29][16] * mat_B[16][8] +
                  mat_A[29][17] * mat_B[17][8] +
                  mat_A[29][18] * mat_B[18][8] +
                  mat_A[29][19] * mat_B[19][8] +
                  mat_A[29][20] * mat_B[20][8] +
                  mat_A[29][21] * mat_B[21][8] +
                  mat_A[29][22] * mat_B[22][8] +
                  mat_A[29][23] * mat_B[23][8] +
                  mat_A[29][24] * mat_B[24][8] +
                  mat_A[29][25] * mat_B[25][8] +
                  mat_A[29][26] * mat_B[26][8] +
                  mat_A[29][27] * mat_B[27][8] +
                  mat_A[29][28] * mat_B[28][8] +
                  mat_A[29][29] * mat_B[29][8] +
                  mat_A[29][30] * mat_B[30][8] +
                  mat_A[29][31] * mat_B[31][8];
    mat_C[29][9] <= 
                  mat_A[29][0] * mat_B[0][9] +
                  mat_A[29][1] * mat_B[1][9] +
                  mat_A[29][2] * mat_B[2][9] +
                  mat_A[29][3] * mat_B[3][9] +
                  mat_A[29][4] * mat_B[4][9] +
                  mat_A[29][5] * mat_B[5][9] +
                  mat_A[29][6] * mat_B[6][9] +
                  mat_A[29][7] * mat_B[7][9] +
                  mat_A[29][8] * mat_B[8][9] +
                  mat_A[29][9] * mat_B[9][9] +
                  mat_A[29][10] * mat_B[10][9] +
                  mat_A[29][11] * mat_B[11][9] +
                  mat_A[29][12] * mat_B[12][9] +
                  mat_A[29][13] * mat_B[13][9] +
                  mat_A[29][14] * mat_B[14][9] +
                  mat_A[29][15] * mat_B[15][9] +
                  mat_A[29][16] * mat_B[16][9] +
                  mat_A[29][17] * mat_B[17][9] +
                  mat_A[29][18] * mat_B[18][9] +
                  mat_A[29][19] * mat_B[19][9] +
                  mat_A[29][20] * mat_B[20][9] +
                  mat_A[29][21] * mat_B[21][9] +
                  mat_A[29][22] * mat_B[22][9] +
                  mat_A[29][23] * mat_B[23][9] +
                  mat_A[29][24] * mat_B[24][9] +
                  mat_A[29][25] * mat_B[25][9] +
                  mat_A[29][26] * mat_B[26][9] +
                  mat_A[29][27] * mat_B[27][9] +
                  mat_A[29][28] * mat_B[28][9] +
                  mat_A[29][29] * mat_B[29][9] +
                  mat_A[29][30] * mat_B[30][9] +
                  mat_A[29][31] * mat_B[31][9];
    mat_C[29][10] <= 
                  mat_A[29][0] * mat_B[0][10] +
                  mat_A[29][1] * mat_B[1][10] +
                  mat_A[29][2] * mat_B[2][10] +
                  mat_A[29][3] * mat_B[3][10] +
                  mat_A[29][4] * mat_B[4][10] +
                  mat_A[29][5] * mat_B[5][10] +
                  mat_A[29][6] * mat_B[6][10] +
                  mat_A[29][7] * mat_B[7][10] +
                  mat_A[29][8] * mat_B[8][10] +
                  mat_A[29][9] * mat_B[9][10] +
                  mat_A[29][10] * mat_B[10][10] +
                  mat_A[29][11] * mat_B[11][10] +
                  mat_A[29][12] * mat_B[12][10] +
                  mat_A[29][13] * mat_B[13][10] +
                  mat_A[29][14] * mat_B[14][10] +
                  mat_A[29][15] * mat_B[15][10] +
                  mat_A[29][16] * mat_B[16][10] +
                  mat_A[29][17] * mat_B[17][10] +
                  mat_A[29][18] * mat_B[18][10] +
                  mat_A[29][19] * mat_B[19][10] +
                  mat_A[29][20] * mat_B[20][10] +
                  mat_A[29][21] * mat_B[21][10] +
                  mat_A[29][22] * mat_B[22][10] +
                  mat_A[29][23] * mat_B[23][10] +
                  mat_A[29][24] * mat_B[24][10] +
                  mat_A[29][25] * mat_B[25][10] +
                  mat_A[29][26] * mat_B[26][10] +
                  mat_A[29][27] * mat_B[27][10] +
                  mat_A[29][28] * mat_B[28][10] +
                  mat_A[29][29] * mat_B[29][10] +
                  mat_A[29][30] * mat_B[30][10] +
                  mat_A[29][31] * mat_B[31][10];
    mat_C[29][11] <= 
                  mat_A[29][0] * mat_B[0][11] +
                  mat_A[29][1] * mat_B[1][11] +
                  mat_A[29][2] * mat_B[2][11] +
                  mat_A[29][3] * mat_B[3][11] +
                  mat_A[29][4] * mat_B[4][11] +
                  mat_A[29][5] * mat_B[5][11] +
                  mat_A[29][6] * mat_B[6][11] +
                  mat_A[29][7] * mat_B[7][11] +
                  mat_A[29][8] * mat_B[8][11] +
                  mat_A[29][9] * mat_B[9][11] +
                  mat_A[29][10] * mat_B[10][11] +
                  mat_A[29][11] * mat_B[11][11] +
                  mat_A[29][12] * mat_B[12][11] +
                  mat_A[29][13] * mat_B[13][11] +
                  mat_A[29][14] * mat_B[14][11] +
                  mat_A[29][15] * mat_B[15][11] +
                  mat_A[29][16] * mat_B[16][11] +
                  mat_A[29][17] * mat_B[17][11] +
                  mat_A[29][18] * mat_B[18][11] +
                  mat_A[29][19] * mat_B[19][11] +
                  mat_A[29][20] * mat_B[20][11] +
                  mat_A[29][21] * mat_B[21][11] +
                  mat_A[29][22] * mat_B[22][11] +
                  mat_A[29][23] * mat_B[23][11] +
                  mat_A[29][24] * mat_B[24][11] +
                  mat_A[29][25] * mat_B[25][11] +
                  mat_A[29][26] * mat_B[26][11] +
                  mat_A[29][27] * mat_B[27][11] +
                  mat_A[29][28] * mat_B[28][11] +
                  mat_A[29][29] * mat_B[29][11] +
                  mat_A[29][30] * mat_B[30][11] +
                  mat_A[29][31] * mat_B[31][11];
    mat_C[29][12] <= 
                  mat_A[29][0] * mat_B[0][12] +
                  mat_A[29][1] * mat_B[1][12] +
                  mat_A[29][2] * mat_B[2][12] +
                  mat_A[29][3] * mat_B[3][12] +
                  mat_A[29][4] * mat_B[4][12] +
                  mat_A[29][5] * mat_B[5][12] +
                  mat_A[29][6] * mat_B[6][12] +
                  mat_A[29][7] * mat_B[7][12] +
                  mat_A[29][8] * mat_B[8][12] +
                  mat_A[29][9] * mat_B[9][12] +
                  mat_A[29][10] * mat_B[10][12] +
                  mat_A[29][11] * mat_B[11][12] +
                  mat_A[29][12] * mat_B[12][12] +
                  mat_A[29][13] * mat_B[13][12] +
                  mat_A[29][14] * mat_B[14][12] +
                  mat_A[29][15] * mat_B[15][12] +
                  mat_A[29][16] * mat_B[16][12] +
                  mat_A[29][17] * mat_B[17][12] +
                  mat_A[29][18] * mat_B[18][12] +
                  mat_A[29][19] * mat_B[19][12] +
                  mat_A[29][20] * mat_B[20][12] +
                  mat_A[29][21] * mat_B[21][12] +
                  mat_A[29][22] * mat_B[22][12] +
                  mat_A[29][23] * mat_B[23][12] +
                  mat_A[29][24] * mat_B[24][12] +
                  mat_A[29][25] * mat_B[25][12] +
                  mat_A[29][26] * mat_B[26][12] +
                  mat_A[29][27] * mat_B[27][12] +
                  mat_A[29][28] * mat_B[28][12] +
                  mat_A[29][29] * mat_B[29][12] +
                  mat_A[29][30] * mat_B[30][12] +
                  mat_A[29][31] * mat_B[31][12];
    mat_C[29][13] <= 
                  mat_A[29][0] * mat_B[0][13] +
                  mat_A[29][1] * mat_B[1][13] +
                  mat_A[29][2] * mat_B[2][13] +
                  mat_A[29][3] * mat_B[3][13] +
                  mat_A[29][4] * mat_B[4][13] +
                  mat_A[29][5] * mat_B[5][13] +
                  mat_A[29][6] * mat_B[6][13] +
                  mat_A[29][7] * mat_B[7][13] +
                  mat_A[29][8] * mat_B[8][13] +
                  mat_A[29][9] * mat_B[9][13] +
                  mat_A[29][10] * mat_B[10][13] +
                  mat_A[29][11] * mat_B[11][13] +
                  mat_A[29][12] * mat_B[12][13] +
                  mat_A[29][13] * mat_B[13][13] +
                  mat_A[29][14] * mat_B[14][13] +
                  mat_A[29][15] * mat_B[15][13] +
                  mat_A[29][16] * mat_B[16][13] +
                  mat_A[29][17] * mat_B[17][13] +
                  mat_A[29][18] * mat_B[18][13] +
                  mat_A[29][19] * mat_B[19][13] +
                  mat_A[29][20] * mat_B[20][13] +
                  mat_A[29][21] * mat_B[21][13] +
                  mat_A[29][22] * mat_B[22][13] +
                  mat_A[29][23] * mat_B[23][13] +
                  mat_A[29][24] * mat_B[24][13] +
                  mat_A[29][25] * mat_B[25][13] +
                  mat_A[29][26] * mat_B[26][13] +
                  mat_A[29][27] * mat_B[27][13] +
                  mat_A[29][28] * mat_B[28][13] +
                  mat_A[29][29] * mat_B[29][13] +
                  mat_A[29][30] * mat_B[30][13] +
                  mat_A[29][31] * mat_B[31][13];
    mat_C[29][14] <= 
                  mat_A[29][0] * mat_B[0][14] +
                  mat_A[29][1] * mat_B[1][14] +
                  mat_A[29][2] * mat_B[2][14] +
                  mat_A[29][3] * mat_B[3][14] +
                  mat_A[29][4] * mat_B[4][14] +
                  mat_A[29][5] * mat_B[5][14] +
                  mat_A[29][6] * mat_B[6][14] +
                  mat_A[29][7] * mat_B[7][14] +
                  mat_A[29][8] * mat_B[8][14] +
                  mat_A[29][9] * mat_B[9][14] +
                  mat_A[29][10] * mat_B[10][14] +
                  mat_A[29][11] * mat_B[11][14] +
                  mat_A[29][12] * mat_B[12][14] +
                  mat_A[29][13] * mat_B[13][14] +
                  mat_A[29][14] * mat_B[14][14] +
                  mat_A[29][15] * mat_B[15][14] +
                  mat_A[29][16] * mat_B[16][14] +
                  mat_A[29][17] * mat_B[17][14] +
                  mat_A[29][18] * mat_B[18][14] +
                  mat_A[29][19] * mat_B[19][14] +
                  mat_A[29][20] * mat_B[20][14] +
                  mat_A[29][21] * mat_B[21][14] +
                  mat_A[29][22] * mat_B[22][14] +
                  mat_A[29][23] * mat_B[23][14] +
                  mat_A[29][24] * mat_B[24][14] +
                  mat_A[29][25] * mat_B[25][14] +
                  mat_A[29][26] * mat_B[26][14] +
                  mat_A[29][27] * mat_B[27][14] +
                  mat_A[29][28] * mat_B[28][14] +
                  mat_A[29][29] * mat_B[29][14] +
                  mat_A[29][30] * mat_B[30][14] +
                  mat_A[29][31] * mat_B[31][14];
    mat_C[29][15] <= 
                  mat_A[29][0] * mat_B[0][15] +
                  mat_A[29][1] * mat_B[1][15] +
                  mat_A[29][2] * mat_B[2][15] +
                  mat_A[29][3] * mat_B[3][15] +
                  mat_A[29][4] * mat_B[4][15] +
                  mat_A[29][5] * mat_B[5][15] +
                  mat_A[29][6] * mat_B[6][15] +
                  mat_A[29][7] * mat_B[7][15] +
                  mat_A[29][8] * mat_B[8][15] +
                  mat_A[29][9] * mat_B[9][15] +
                  mat_A[29][10] * mat_B[10][15] +
                  mat_A[29][11] * mat_B[11][15] +
                  mat_A[29][12] * mat_B[12][15] +
                  mat_A[29][13] * mat_B[13][15] +
                  mat_A[29][14] * mat_B[14][15] +
                  mat_A[29][15] * mat_B[15][15] +
                  mat_A[29][16] * mat_B[16][15] +
                  mat_A[29][17] * mat_B[17][15] +
                  mat_A[29][18] * mat_B[18][15] +
                  mat_A[29][19] * mat_B[19][15] +
                  mat_A[29][20] * mat_B[20][15] +
                  mat_A[29][21] * mat_B[21][15] +
                  mat_A[29][22] * mat_B[22][15] +
                  mat_A[29][23] * mat_B[23][15] +
                  mat_A[29][24] * mat_B[24][15] +
                  mat_A[29][25] * mat_B[25][15] +
                  mat_A[29][26] * mat_B[26][15] +
                  mat_A[29][27] * mat_B[27][15] +
                  mat_A[29][28] * mat_B[28][15] +
                  mat_A[29][29] * mat_B[29][15] +
                  mat_A[29][30] * mat_B[30][15] +
                  mat_A[29][31] * mat_B[31][15];
    mat_C[29][16] <= 
                  mat_A[29][0] * mat_B[0][16] +
                  mat_A[29][1] * mat_B[1][16] +
                  mat_A[29][2] * mat_B[2][16] +
                  mat_A[29][3] * mat_B[3][16] +
                  mat_A[29][4] * mat_B[4][16] +
                  mat_A[29][5] * mat_B[5][16] +
                  mat_A[29][6] * mat_B[6][16] +
                  mat_A[29][7] * mat_B[7][16] +
                  mat_A[29][8] * mat_B[8][16] +
                  mat_A[29][9] * mat_B[9][16] +
                  mat_A[29][10] * mat_B[10][16] +
                  mat_A[29][11] * mat_B[11][16] +
                  mat_A[29][12] * mat_B[12][16] +
                  mat_A[29][13] * mat_B[13][16] +
                  mat_A[29][14] * mat_B[14][16] +
                  mat_A[29][15] * mat_B[15][16] +
                  mat_A[29][16] * mat_B[16][16] +
                  mat_A[29][17] * mat_B[17][16] +
                  mat_A[29][18] * mat_B[18][16] +
                  mat_A[29][19] * mat_B[19][16] +
                  mat_A[29][20] * mat_B[20][16] +
                  mat_A[29][21] * mat_B[21][16] +
                  mat_A[29][22] * mat_B[22][16] +
                  mat_A[29][23] * mat_B[23][16] +
                  mat_A[29][24] * mat_B[24][16] +
                  mat_A[29][25] * mat_B[25][16] +
                  mat_A[29][26] * mat_B[26][16] +
                  mat_A[29][27] * mat_B[27][16] +
                  mat_A[29][28] * mat_B[28][16] +
                  mat_A[29][29] * mat_B[29][16] +
                  mat_A[29][30] * mat_B[30][16] +
                  mat_A[29][31] * mat_B[31][16];
    mat_C[29][17] <= 
                  mat_A[29][0] * mat_B[0][17] +
                  mat_A[29][1] * mat_B[1][17] +
                  mat_A[29][2] * mat_B[2][17] +
                  mat_A[29][3] * mat_B[3][17] +
                  mat_A[29][4] * mat_B[4][17] +
                  mat_A[29][5] * mat_B[5][17] +
                  mat_A[29][6] * mat_B[6][17] +
                  mat_A[29][7] * mat_B[7][17] +
                  mat_A[29][8] * mat_B[8][17] +
                  mat_A[29][9] * mat_B[9][17] +
                  mat_A[29][10] * mat_B[10][17] +
                  mat_A[29][11] * mat_B[11][17] +
                  mat_A[29][12] * mat_B[12][17] +
                  mat_A[29][13] * mat_B[13][17] +
                  mat_A[29][14] * mat_B[14][17] +
                  mat_A[29][15] * mat_B[15][17] +
                  mat_A[29][16] * mat_B[16][17] +
                  mat_A[29][17] * mat_B[17][17] +
                  mat_A[29][18] * mat_B[18][17] +
                  mat_A[29][19] * mat_B[19][17] +
                  mat_A[29][20] * mat_B[20][17] +
                  mat_A[29][21] * mat_B[21][17] +
                  mat_A[29][22] * mat_B[22][17] +
                  mat_A[29][23] * mat_B[23][17] +
                  mat_A[29][24] * mat_B[24][17] +
                  mat_A[29][25] * mat_B[25][17] +
                  mat_A[29][26] * mat_B[26][17] +
                  mat_A[29][27] * mat_B[27][17] +
                  mat_A[29][28] * mat_B[28][17] +
                  mat_A[29][29] * mat_B[29][17] +
                  mat_A[29][30] * mat_B[30][17] +
                  mat_A[29][31] * mat_B[31][17];
    mat_C[29][18] <= 
                  mat_A[29][0] * mat_B[0][18] +
                  mat_A[29][1] * mat_B[1][18] +
                  mat_A[29][2] * mat_B[2][18] +
                  mat_A[29][3] * mat_B[3][18] +
                  mat_A[29][4] * mat_B[4][18] +
                  mat_A[29][5] * mat_B[5][18] +
                  mat_A[29][6] * mat_B[6][18] +
                  mat_A[29][7] * mat_B[7][18] +
                  mat_A[29][8] * mat_B[8][18] +
                  mat_A[29][9] * mat_B[9][18] +
                  mat_A[29][10] * mat_B[10][18] +
                  mat_A[29][11] * mat_B[11][18] +
                  mat_A[29][12] * mat_B[12][18] +
                  mat_A[29][13] * mat_B[13][18] +
                  mat_A[29][14] * mat_B[14][18] +
                  mat_A[29][15] * mat_B[15][18] +
                  mat_A[29][16] * mat_B[16][18] +
                  mat_A[29][17] * mat_B[17][18] +
                  mat_A[29][18] * mat_B[18][18] +
                  mat_A[29][19] * mat_B[19][18] +
                  mat_A[29][20] * mat_B[20][18] +
                  mat_A[29][21] * mat_B[21][18] +
                  mat_A[29][22] * mat_B[22][18] +
                  mat_A[29][23] * mat_B[23][18] +
                  mat_A[29][24] * mat_B[24][18] +
                  mat_A[29][25] * mat_B[25][18] +
                  mat_A[29][26] * mat_B[26][18] +
                  mat_A[29][27] * mat_B[27][18] +
                  mat_A[29][28] * mat_B[28][18] +
                  mat_A[29][29] * mat_B[29][18] +
                  mat_A[29][30] * mat_B[30][18] +
                  mat_A[29][31] * mat_B[31][18];
    mat_C[29][19] <= 
                  mat_A[29][0] * mat_B[0][19] +
                  mat_A[29][1] * mat_B[1][19] +
                  mat_A[29][2] * mat_B[2][19] +
                  mat_A[29][3] * mat_B[3][19] +
                  mat_A[29][4] * mat_B[4][19] +
                  mat_A[29][5] * mat_B[5][19] +
                  mat_A[29][6] * mat_B[6][19] +
                  mat_A[29][7] * mat_B[7][19] +
                  mat_A[29][8] * mat_B[8][19] +
                  mat_A[29][9] * mat_B[9][19] +
                  mat_A[29][10] * mat_B[10][19] +
                  mat_A[29][11] * mat_B[11][19] +
                  mat_A[29][12] * mat_B[12][19] +
                  mat_A[29][13] * mat_B[13][19] +
                  mat_A[29][14] * mat_B[14][19] +
                  mat_A[29][15] * mat_B[15][19] +
                  mat_A[29][16] * mat_B[16][19] +
                  mat_A[29][17] * mat_B[17][19] +
                  mat_A[29][18] * mat_B[18][19] +
                  mat_A[29][19] * mat_B[19][19] +
                  mat_A[29][20] * mat_B[20][19] +
                  mat_A[29][21] * mat_B[21][19] +
                  mat_A[29][22] * mat_B[22][19] +
                  mat_A[29][23] * mat_B[23][19] +
                  mat_A[29][24] * mat_B[24][19] +
                  mat_A[29][25] * mat_B[25][19] +
                  mat_A[29][26] * mat_B[26][19] +
                  mat_A[29][27] * mat_B[27][19] +
                  mat_A[29][28] * mat_B[28][19] +
                  mat_A[29][29] * mat_B[29][19] +
                  mat_A[29][30] * mat_B[30][19] +
                  mat_A[29][31] * mat_B[31][19];
    mat_C[29][20] <= 
                  mat_A[29][0] * mat_B[0][20] +
                  mat_A[29][1] * mat_B[1][20] +
                  mat_A[29][2] * mat_B[2][20] +
                  mat_A[29][3] * mat_B[3][20] +
                  mat_A[29][4] * mat_B[4][20] +
                  mat_A[29][5] * mat_B[5][20] +
                  mat_A[29][6] * mat_B[6][20] +
                  mat_A[29][7] * mat_B[7][20] +
                  mat_A[29][8] * mat_B[8][20] +
                  mat_A[29][9] * mat_B[9][20] +
                  mat_A[29][10] * mat_B[10][20] +
                  mat_A[29][11] * mat_B[11][20] +
                  mat_A[29][12] * mat_B[12][20] +
                  mat_A[29][13] * mat_B[13][20] +
                  mat_A[29][14] * mat_B[14][20] +
                  mat_A[29][15] * mat_B[15][20] +
                  mat_A[29][16] * mat_B[16][20] +
                  mat_A[29][17] * mat_B[17][20] +
                  mat_A[29][18] * mat_B[18][20] +
                  mat_A[29][19] * mat_B[19][20] +
                  mat_A[29][20] * mat_B[20][20] +
                  mat_A[29][21] * mat_B[21][20] +
                  mat_A[29][22] * mat_B[22][20] +
                  mat_A[29][23] * mat_B[23][20] +
                  mat_A[29][24] * mat_B[24][20] +
                  mat_A[29][25] * mat_B[25][20] +
                  mat_A[29][26] * mat_B[26][20] +
                  mat_A[29][27] * mat_B[27][20] +
                  mat_A[29][28] * mat_B[28][20] +
                  mat_A[29][29] * mat_B[29][20] +
                  mat_A[29][30] * mat_B[30][20] +
                  mat_A[29][31] * mat_B[31][20];
    mat_C[29][21] <= 
                  mat_A[29][0] * mat_B[0][21] +
                  mat_A[29][1] * mat_B[1][21] +
                  mat_A[29][2] * mat_B[2][21] +
                  mat_A[29][3] * mat_B[3][21] +
                  mat_A[29][4] * mat_B[4][21] +
                  mat_A[29][5] * mat_B[5][21] +
                  mat_A[29][6] * mat_B[6][21] +
                  mat_A[29][7] * mat_B[7][21] +
                  mat_A[29][8] * mat_B[8][21] +
                  mat_A[29][9] * mat_B[9][21] +
                  mat_A[29][10] * mat_B[10][21] +
                  mat_A[29][11] * mat_B[11][21] +
                  mat_A[29][12] * mat_B[12][21] +
                  mat_A[29][13] * mat_B[13][21] +
                  mat_A[29][14] * mat_B[14][21] +
                  mat_A[29][15] * mat_B[15][21] +
                  mat_A[29][16] * mat_B[16][21] +
                  mat_A[29][17] * mat_B[17][21] +
                  mat_A[29][18] * mat_B[18][21] +
                  mat_A[29][19] * mat_B[19][21] +
                  mat_A[29][20] * mat_B[20][21] +
                  mat_A[29][21] * mat_B[21][21] +
                  mat_A[29][22] * mat_B[22][21] +
                  mat_A[29][23] * mat_B[23][21] +
                  mat_A[29][24] * mat_B[24][21] +
                  mat_A[29][25] * mat_B[25][21] +
                  mat_A[29][26] * mat_B[26][21] +
                  mat_A[29][27] * mat_B[27][21] +
                  mat_A[29][28] * mat_B[28][21] +
                  mat_A[29][29] * mat_B[29][21] +
                  mat_A[29][30] * mat_B[30][21] +
                  mat_A[29][31] * mat_B[31][21];
    mat_C[29][22] <= 
                  mat_A[29][0] * mat_B[0][22] +
                  mat_A[29][1] * mat_B[1][22] +
                  mat_A[29][2] * mat_B[2][22] +
                  mat_A[29][3] * mat_B[3][22] +
                  mat_A[29][4] * mat_B[4][22] +
                  mat_A[29][5] * mat_B[5][22] +
                  mat_A[29][6] * mat_B[6][22] +
                  mat_A[29][7] * mat_B[7][22] +
                  mat_A[29][8] * mat_B[8][22] +
                  mat_A[29][9] * mat_B[9][22] +
                  mat_A[29][10] * mat_B[10][22] +
                  mat_A[29][11] * mat_B[11][22] +
                  mat_A[29][12] * mat_B[12][22] +
                  mat_A[29][13] * mat_B[13][22] +
                  mat_A[29][14] * mat_B[14][22] +
                  mat_A[29][15] * mat_B[15][22] +
                  mat_A[29][16] * mat_B[16][22] +
                  mat_A[29][17] * mat_B[17][22] +
                  mat_A[29][18] * mat_B[18][22] +
                  mat_A[29][19] * mat_B[19][22] +
                  mat_A[29][20] * mat_B[20][22] +
                  mat_A[29][21] * mat_B[21][22] +
                  mat_A[29][22] * mat_B[22][22] +
                  mat_A[29][23] * mat_B[23][22] +
                  mat_A[29][24] * mat_B[24][22] +
                  mat_A[29][25] * mat_B[25][22] +
                  mat_A[29][26] * mat_B[26][22] +
                  mat_A[29][27] * mat_B[27][22] +
                  mat_A[29][28] * mat_B[28][22] +
                  mat_A[29][29] * mat_B[29][22] +
                  mat_A[29][30] * mat_B[30][22] +
                  mat_A[29][31] * mat_B[31][22];
    mat_C[29][23] <= 
                  mat_A[29][0] * mat_B[0][23] +
                  mat_A[29][1] * mat_B[1][23] +
                  mat_A[29][2] * mat_B[2][23] +
                  mat_A[29][3] * mat_B[3][23] +
                  mat_A[29][4] * mat_B[4][23] +
                  mat_A[29][5] * mat_B[5][23] +
                  mat_A[29][6] * mat_B[6][23] +
                  mat_A[29][7] * mat_B[7][23] +
                  mat_A[29][8] * mat_B[8][23] +
                  mat_A[29][9] * mat_B[9][23] +
                  mat_A[29][10] * mat_B[10][23] +
                  mat_A[29][11] * mat_B[11][23] +
                  mat_A[29][12] * mat_B[12][23] +
                  mat_A[29][13] * mat_B[13][23] +
                  mat_A[29][14] * mat_B[14][23] +
                  mat_A[29][15] * mat_B[15][23] +
                  mat_A[29][16] * mat_B[16][23] +
                  mat_A[29][17] * mat_B[17][23] +
                  mat_A[29][18] * mat_B[18][23] +
                  mat_A[29][19] * mat_B[19][23] +
                  mat_A[29][20] * mat_B[20][23] +
                  mat_A[29][21] * mat_B[21][23] +
                  mat_A[29][22] * mat_B[22][23] +
                  mat_A[29][23] * mat_B[23][23] +
                  mat_A[29][24] * mat_B[24][23] +
                  mat_A[29][25] * mat_B[25][23] +
                  mat_A[29][26] * mat_B[26][23] +
                  mat_A[29][27] * mat_B[27][23] +
                  mat_A[29][28] * mat_B[28][23] +
                  mat_A[29][29] * mat_B[29][23] +
                  mat_A[29][30] * mat_B[30][23] +
                  mat_A[29][31] * mat_B[31][23];
    mat_C[29][24] <= 
                  mat_A[29][0] * mat_B[0][24] +
                  mat_A[29][1] * mat_B[1][24] +
                  mat_A[29][2] * mat_B[2][24] +
                  mat_A[29][3] * mat_B[3][24] +
                  mat_A[29][4] * mat_B[4][24] +
                  mat_A[29][5] * mat_B[5][24] +
                  mat_A[29][6] * mat_B[6][24] +
                  mat_A[29][7] * mat_B[7][24] +
                  mat_A[29][8] * mat_B[8][24] +
                  mat_A[29][9] * mat_B[9][24] +
                  mat_A[29][10] * mat_B[10][24] +
                  mat_A[29][11] * mat_B[11][24] +
                  mat_A[29][12] * mat_B[12][24] +
                  mat_A[29][13] * mat_B[13][24] +
                  mat_A[29][14] * mat_B[14][24] +
                  mat_A[29][15] * mat_B[15][24] +
                  mat_A[29][16] * mat_B[16][24] +
                  mat_A[29][17] * mat_B[17][24] +
                  mat_A[29][18] * mat_B[18][24] +
                  mat_A[29][19] * mat_B[19][24] +
                  mat_A[29][20] * mat_B[20][24] +
                  mat_A[29][21] * mat_B[21][24] +
                  mat_A[29][22] * mat_B[22][24] +
                  mat_A[29][23] * mat_B[23][24] +
                  mat_A[29][24] * mat_B[24][24] +
                  mat_A[29][25] * mat_B[25][24] +
                  mat_A[29][26] * mat_B[26][24] +
                  mat_A[29][27] * mat_B[27][24] +
                  mat_A[29][28] * mat_B[28][24] +
                  mat_A[29][29] * mat_B[29][24] +
                  mat_A[29][30] * mat_B[30][24] +
                  mat_A[29][31] * mat_B[31][24];
    mat_C[29][25] <= 
                  mat_A[29][0] * mat_B[0][25] +
                  mat_A[29][1] * mat_B[1][25] +
                  mat_A[29][2] * mat_B[2][25] +
                  mat_A[29][3] * mat_B[3][25] +
                  mat_A[29][4] * mat_B[4][25] +
                  mat_A[29][5] * mat_B[5][25] +
                  mat_A[29][6] * mat_B[6][25] +
                  mat_A[29][7] * mat_B[7][25] +
                  mat_A[29][8] * mat_B[8][25] +
                  mat_A[29][9] * mat_B[9][25] +
                  mat_A[29][10] * mat_B[10][25] +
                  mat_A[29][11] * mat_B[11][25] +
                  mat_A[29][12] * mat_B[12][25] +
                  mat_A[29][13] * mat_B[13][25] +
                  mat_A[29][14] * mat_B[14][25] +
                  mat_A[29][15] * mat_B[15][25] +
                  mat_A[29][16] * mat_B[16][25] +
                  mat_A[29][17] * mat_B[17][25] +
                  mat_A[29][18] * mat_B[18][25] +
                  mat_A[29][19] * mat_B[19][25] +
                  mat_A[29][20] * mat_B[20][25] +
                  mat_A[29][21] * mat_B[21][25] +
                  mat_A[29][22] * mat_B[22][25] +
                  mat_A[29][23] * mat_B[23][25] +
                  mat_A[29][24] * mat_B[24][25] +
                  mat_A[29][25] * mat_B[25][25] +
                  mat_A[29][26] * mat_B[26][25] +
                  mat_A[29][27] * mat_B[27][25] +
                  mat_A[29][28] * mat_B[28][25] +
                  mat_A[29][29] * mat_B[29][25] +
                  mat_A[29][30] * mat_B[30][25] +
                  mat_A[29][31] * mat_B[31][25];
    mat_C[29][26] <= 
                  mat_A[29][0] * mat_B[0][26] +
                  mat_A[29][1] * mat_B[1][26] +
                  mat_A[29][2] * mat_B[2][26] +
                  mat_A[29][3] * mat_B[3][26] +
                  mat_A[29][4] * mat_B[4][26] +
                  mat_A[29][5] * mat_B[5][26] +
                  mat_A[29][6] * mat_B[6][26] +
                  mat_A[29][7] * mat_B[7][26] +
                  mat_A[29][8] * mat_B[8][26] +
                  mat_A[29][9] * mat_B[9][26] +
                  mat_A[29][10] * mat_B[10][26] +
                  mat_A[29][11] * mat_B[11][26] +
                  mat_A[29][12] * mat_B[12][26] +
                  mat_A[29][13] * mat_B[13][26] +
                  mat_A[29][14] * mat_B[14][26] +
                  mat_A[29][15] * mat_B[15][26] +
                  mat_A[29][16] * mat_B[16][26] +
                  mat_A[29][17] * mat_B[17][26] +
                  mat_A[29][18] * mat_B[18][26] +
                  mat_A[29][19] * mat_B[19][26] +
                  mat_A[29][20] * mat_B[20][26] +
                  mat_A[29][21] * mat_B[21][26] +
                  mat_A[29][22] * mat_B[22][26] +
                  mat_A[29][23] * mat_B[23][26] +
                  mat_A[29][24] * mat_B[24][26] +
                  mat_A[29][25] * mat_B[25][26] +
                  mat_A[29][26] * mat_B[26][26] +
                  mat_A[29][27] * mat_B[27][26] +
                  mat_A[29][28] * mat_B[28][26] +
                  mat_A[29][29] * mat_B[29][26] +
                  mat_A[29][30] * mat_B[30][26] +
                  mat_A[29][31] * mat_B[31][26];
    mat_C[29][27] <= 
                  mat_A[29][0] * mat_B[0][27] +
                  mat_A[29][1] * mat_B[1][27] +
                  mat_A[29][2] * mat_B[2][27] +
                  mat_A[29][3] * mat_B[3][27] +
                  mat_A[29][4] * mat_B[4][27] +
                  mat_A[29][5] * mat_B[5][27] +
                  mat_A[29][6] * mat_B[6][27] +
                  mat_A[29][7] * mat_B[7][27] +
                  mat_A[29][8] * mat_B[8][27] +
                  mat_A[29][9] * mat_B[9][27] +
                  mat_A[29][10] * mat_B[10][27] +
                  mat_A[29][11] * mat_B[11][27] +
                  mat_A[29][12] * mat_B[12][27] +
                  mat_A[29][13] * mat_B[13][27] +
                  mat_A[29][14] * mat_B[14][27] +
                  mat_A[29][15] * mat_B[15][27] +
                  mat_A[29][16] * mat_B[16][27] +
                  mat_A[29][17] * mat_B[17][27] +
                  mat_A[29][18] * mat_B[18][27] +
                  mat_A[29][19] * mat_B[19][27] +
                  mat_A[29][20] * mat_B[20][27] +
                  mat_A[29][21] * mat_B[21][27] +
                  mat_A[29][22] * mat_B[22][27] +
                  mat_A[29][23] * mat_B[23][27] +
                  mat_A[29][24] * mat_B[24][27] +
                  mat_A[29][25] * mat_B[25][27] +
                  mat_A[29][26] * mat_B[26][27] +
                  mat_A[29][27] * mat_B[27][27] +
                  mat_A[29][28] * mat_B[28][27] +
                  mat_A[29][29] * mat_B[29][27] +
                  mat_A[29][30] * mat_B[30][27] +
                  mat_A[29][31] * mat_B[31][27];
    mat_C[29][28] <= 
                  mat_A[29][0] * mat_B[0][28] +
                  mat_A[29][1] * mat_B[1][28] +
                  mat_A[29][2] * mat_B[2][28] +
                  mat_A[29][3] * mat_B[3][28] +
                  mat_A[29][4] * mat_B[4][28] +
                  mat_A[29][5] * mat_B[5][28] +
                  mat_A[29][6] * mat_B[6][28] +
                  mat_A[29][7] * mat_B[7][28] +
                  mat_A[29][8] * mat_B[8][28] +
                  mat_A[29][9] * mat_B[9][28] +
                  mat_A[29][10] * mat_B[10][28] +
                  mat_A[29][11] * mat_B[11][28] +
                  mat_A[29][12] * mat_B[12][28] +
                  mat_A[29][13] * mat_B[13][28] +
                  mat_A[29][14] * mat_B[14][28] +
                  mat_A[29][15] * mat_B[15][28] +
                  mat_A[29][16] * mat_B[16][28] +
                  mat_A[29][17] * mat_B[17][28] +
                  mat_A[29][18] * mat_B[18][28] +
                  mat_A[29][19] * mat_B[19][28] +
                  mat_A[29][20] * mat_B[20][28] +
                  mat_A[29][21] * mat_B[21][28] +
                  mat_A[29][22] * mat_B[22][28] +
                  mat_A[29][23] * mat_B[23][28] +
                  mat_A[29][24] * mat_B[24][28] +
                  mat_A[29][25] * mat_B[25][28] +
                  mat_A[29][26] * mat_B[26][28] +
                  mat_A[29][27] * mat_B[27][28] +
                  mat_A[29][28] * mat_B[28][28] +
                  mat_A[29][29] * mat_B[29][28] +
                  mat_A[29][30] * mat_B[30][28] +
                  mat_A[29][31] * mat_B[31][28];
    mat_C[29][29] <= 
                  mat_A[29][0] * mat_B[0][29] +
                  mat_A[29][1] * mat_B[1][29] +
                  mat_A[29][2] * mat_B[2][29] +
                  mat_A[29][3] * mat_B[3][29] +
                  mat_A[29][4] * mat_B[4][29] +
                  mat_A[29][5] * mat_B[5][29] +
                  mat_A[29][6] * mat_B[6][29] +
                  mat_A[29][7] * mat_B[7][29] +
                  mat_A[29][8] * mat_B[8][29] +
                  mat_A[29][9] * mat_B[9][29] +
                  mat_A[29][10] * mat_B[10][29] +
                  mat_A[29][11] * mat_B[11][29] +
                  mat_A[29][12] * mat_B[12][29] +
                  mat_A[29][13] * mat_B[13][29] +
                  mat_A[29][14] * mat_B[14][29] +
                  mat_A[29][15] * mat_B[15][29] +
                  mat_A[29][16] * mat_B[16][29] +
                  mat_A[29][17] * mat_B[17][29] +
                  mat_A[29][18] * mat_B[18][29] +
                  mat_A[29][19] * mat_B[19][29] +
                  mat_A[29][20] * mat_B[20][29] +
                  mat_A[29][21] * mat_B[21][29] +
                  mat_A[29][22] * mat_B[22][29] +
                  mat_A[29][23] * mat_B[23][29] +
                  mat_A[29][24] * mat_B[24][29] +
                  mat_A[29][25] * mat_B[25][29] +
                  mat_A[29][26] * mat_B[26][29] +
                  mat_A[29][27] * mat_B[27][29] +
                  mat_A[29][28] * mat_B[28][29] +
                  mat_A[29][29] * mat_B[29][29] +
                  mat_A[29][30] * mat_B[30][29] +
                  mat_A[29][31] * mat_B[31][29];
    mat_C[29][30] <= 
                  mat_A[29][0] * mat_B[0][30] +
                  mat_A[29][1] * mat_B[1][30] +
                  mat_A[29][2] * mat_B[2][30] +
                  mat_A[29][3] * mat_B[3][30] +
                  mat_A[29][4] * mat_B[4][30] +
                  mat_A[29][5] * mat_B[5][30] +
                  mat_A[29][6] * mat_B[6][30] +
                  mat_A[29][7] * mat_B[7][30] +
                  mat_A[29][8] * mat_B[8][30] +
                  mat_A[29][9] * mat_B[9][30] +
                  mat_A[29][10] * mat_B[10][30] +
                  mat_A[29][11] * mat_B[11][30] +
                  mat_A[29][12] * mat_B[12][30] +
                  mat_A[29][13] * mat_B[13][30] +
                  mat_A[29][14] * mat_B[14][30] +
                  mat_A[29][15] * mat_B[15][30] +
                  mat_A[29][16] * mat_B[16][30] +
                  mat_A[29][17] * mat_B[17][30] +
                  mat_A[29][18] * mat_B[18][30] +
                  mat_A[29][19] * mat_B[19][30] +
                  mat_A[29][20] * mat_B[20][30] +
                  mat_A[29][21] * mat_B[21][30] +
                  mat_A[29][22] * mat_B[22][30] +
                  mat_A[29][23] * mat_B[23][30] +
                  mat_A[29][24] * mat_B[24][30] +
                  mat_A[29][25] * mat_B[25][30] +
                  mat_A[29][26] * mat_B[26][30] +
                  mat_A[29][27] * mat_B[27][30] +
                  mat_A[29][28] * mat_B[28][30] +
                  mat_A[29][29] * mat_B[29][30] +
                  mat_A[29][30] * mat_B[30][30] +
                  mat_A[29][31] * mat_B[31][30];
    mat_C[29][31] <= 
                  mat_A[29][0] * mat_B[0][31] +
                  mat_A[29][1] * mat_B[1][31] +
                  mat_A[29][2] * mat_B[2][31] +
                  mat_A[29][3] * mat_B[3][31] +
                  mat_A[29][4] * mat_B[4][31] +
                  mat_A[29][5] * mat_B[5][31] +
                  mat_A[29][6] * mat_B[6][31] +
                  mat_A[29][7] * mat_B[7][31] +
                  mat_A[29][8] * mat_B[8][31] +
                  mat_A[29][9] * mat_B[9][31] +
                  mat_A[29][10] * mat_B[10][31] +
                  mat_A[29][11] * mat_B[11][31] +
                  mat_A[29][12] * mat_B[12][31] +
                  mat_A[29][13] * mat_B[13][31] +
                  mat_A[29][14] * mat_B[14][31] +
                  mat_A[29][15] * mat_B[15][31] +
                  mat_A[29][16] * mat_B[16][31] +
                  mat_A[29][17] * mat_B[17][31] +
                  mat_A[29][18] * mat_B[18][31] +
                  mat_A[29][19] * mat_B[19][31] +
                  mat_A[29][20] * mat_B[20][31] +
                  mat_A[29][21] * mat_B[21][31] +
                  mat_A[29][22] * mat_B[22][31] +
                  mat_A[29][23] * mat_B[23][31] +
                  mat_A[29][24] * mat_B[24][31] +
                  mat_A[29][25] * mat_B[25][31] +
                  mat_A[29][26] * mat_B[26][31] +
                  mat_A[29][27] * mat_B[27][31] +
                  mat_A[29][28] * mat_B[28][31] +
                  mat_A[29][29] * mat_B[29][31] +
                  mat_A[29][30] * mat_B[30][31] +
                  mat_A[29][31] * mat_B[31][31];
    mat_C[30][0] <= 
                  mat_A[30][0] * mat_B[0][0] +
                  mat_A[30][1] * mat_B[1][0] +
                  mat_A[30][2] * mat_B[2][0] +
                  mat_A[30][3] * mat_B[3][0] +
                  mat_A[30][4] * mat_B[4][0] +
                  mat_A[30][5] * mat_B[5][0] +
                  mat_A[30][6] * mat_B[6][0] +
                  mat_A[30][7] * mat_B[7][0] +
                  mat_A[30][8] * mat_B[8][0] +
                  mat_A[30][9] * mat_B[9][0] +
                  mat_A[30][10] * mat_B[10][0] +
                  mat_A[30][11] * mat_B[11][0] +
                  mat_A[30][12] * mat_B[12][0] +
                  mat_A[30][13] * mat_B[13][0] +
                  mat_A[30][14] * mat_B[14][0] +
                  mat_A[30][15] * mat_B[15][0] +
                  mat_A[30][16] * mat_B[16][0] +
                  mat_A[30][17] * mat_B[17][0] +
                  mat_A[30][18] * mat_B[18][0] +
                  mat_A[30][19] * mat_B[19][0] +
                  mat_A[30][20] * mat_B[20][0] +
                  mat_A[30][21] * mat_B[21][0] +
                  mat_A[30][22] * mat_B[22][0] +
                  mat_A[30][23] * mat_B[23][0] +
                  mat_A[30][24] * mat_B[24][0] +
                  mat_A[30][25] * mat_B[25][0] +
                  mat_A[30][26] * mat_B[26][0] +
                  mat_A[30][27] * mat_B[27][0] +
                  mat_A[30][28] * mat_B[28][0] +
                  mat_A[30][29] * mat_B[29][0] +
                  mat_A[30][30] * mat_B[30][0] +
                  mat_A[30][31] * mat_B[31][0];
    mat_C[30][1] <= 
                  mat_A[30][0] * mat_B[0][1] +
                  mat_A[30][1] * mat_B[1][1] +
                  mat_A[30][2] * mat_B[2][1] +
                  mat_A[30][3] * mat_B[3][1] +
                  mat_A[30][4] * mat_B[4][1] +
                  mat_A[30][5] * mat_B[5][1] +
                  mat_A[30][6] * mat_B[6][1] +
                  mat_A[30][7] * mat_B[7][1] +
                  mat_A[30][8] * mat_B[8][1] +
                  mat_A[30][9] * mat_B[9][1] +
                  mat_A[30][10] * mat_B[10][1] +
                  mat_A[30][11] * mat_B[11][1] +
                  mat_A[30][12] * mat_B[12][1] +
                  mat_A[30][13] * mat_B[13][1] +
                  mat_A[30][14] * mat_B[14][1] +
                  mat_A[30][15] * mat_B[15][1] +
                  mat_A[30][16] * mat_B[16][1] +
                  mat_A[30][17] * mat_B[17][1] +
                  mat_A[30][18] * mat_B[18][1] +
                  mat_A[30][19] * mat_B[19][1] +
                  mat_A[30][20] * mat_B[20][1] +
                  mat_A[30][21] * mat_B[21][1] +
                  mat_A[30][22] * mat_B[22][1] +
                  mat_A[30][23] * mat_B[23][1] +
                  mat_A[30][24] * mat_B[24][1] +
                  mat_A[30][25] * mat_B[25][1] +
                  mat_A[30][26] * mat_B[26][1] +
                  mat_A[30][27] * mat_B[27][1] +
                  mat_A[30][28] * mat_B[28][1] +
                  mat_A[30][29] * mat_B[29][1] +
                  mat_A[30][30] * mat_B[30][1] +
                  mat_A[30][31] * mat_B[31][1];
    mat_C[30][2] <= 
                  mat_A[30][0] * mat_B[0][2] +
                  mat_A[30][1] * mat_B[1][2] +
                  mat_A[30][2] * mat_B[2][2] +
                  mat_A[30][3] * mat_B[3][2] +
                  mat_A[30][4] * mat_B[4][2] +
                  mat_A[30][5] * mat_B[5][2] +
                  mat_A[30][6] * mat_B[6][2] +
                  mat_A[30][7] * mat_B[7][2] +
                  mat_A[30][8] * mat_B[8][2] +
                  mat_A[30][9] * mat_B[9][2] +
                  mat_A[30][10] * mat_B[10][2] +
                  mat_A[30][11] * mat_B[11][2] +
                  mat_A[30][12] * mat_B[12][2] +
                  mat_A[30][13] * mat_B[13][2] +
                  mat_A[30][14] * mat_B[14][2] +
                  mat_A[30][15] * mat_B[15][2] +
                  mat_A[30][16] * mat_B[16][2] +
                  mat_A[30][17] * mat_B[17][2] +
                  mat_A[30][18] * mat_B[18][2] +
                  mat_A[30][19] * mat_B[19][2] +
                  mat_A[30][20] * mat_B[20][2] +
                  mat_A[30][21] * mat_B[21][2] +
                  mat_A[30][22] * mat_B[22][2] +
                  mat_A[30][23] * mat_B[23][2] +
                  mat_A[30][24] * mat_B[24][2] +
                  mat_A[30][25] * mat_B[25][2] +
                  mat_A[30][26] * mat_B[26][2] +
                  mat_A[30][27] * mat_B[27][2] +
                  mat_A[30][28] * mat_B[28][2] +
                  mat_A[30][29] * mat_B[29][2] +
                  mat_A[30][30] * mat_B[30][2] +
                  mat_A[30][31] * mat_B[31][2];
    mat_C[30][3] <= 
                  mat_A[30][0] * mat_B[0][3] +
                  mat_A[30][1] * mat_B[1][3] +
                  mat_A[30][2] * mat_B[2][3] +
                  mat_A[30][3] * mat_B[3][3] +
                  mat_A[30][4] * mat_B[4][3] +
                  mat_A[30][5] * mat_B[5][3] +
                  mat_A[30][6] * mat_B[6][3] +
                  mat_A[30][7] * mat_B[7][3] +
                  mat_A[30][8] * mat_B[8][3] +
                  mat_A[30][9] * mat_B[9][3] +
                  mat_A[30][10] * mat_B[10][3] +
                  mat_A[30][11] * mat_B[11][3] +
                  mat_A[30][12] * mat_B[12][3] +
                  mat_A[30][13] * mat_B[13][3] +
                  mat_A[30][14] * mat_B[14][3] +
                  mat_A[30][15] * mat_B[15][3] +
                  mat_A[30][16] * mat_B[16][3] +
                  mat_A[30][17] * mat_B[17][3] +
                  mat_A[30][18] * mat_B[18][3] +
                  mat_A[30][19] * mat_B[19][3] +
                  mat_A[30][20] * mat_B[20][3] +
                  mat_A[30][21] * mat_B[21][3] +
                  mat_A[30][22] * mat_B[22][3] +
                  mat_A[30][23] * mat_B[23][3] +
                  mat_A[30][24] * mat_B[24][3] +
                  mat_A[30][25] * mat_B[25][3] +
                  mat_A[30][26] * mat_B[26][3] +
                  mat_A[30][27] * mat_B[27][3] +
                  mat_A[30][28] * mat_B[28][3] +
                  mat_A[30][29] * mat_B[29][3] +
                  mat_A[30][30] * mat_B[30][3] +
                  mat_A[30][31] * mat_B[31][3];
    mat_C[30][4] <= 
                  mat_A[30][0] * mat_B[0][4] +
                  mat_A[30][1] * mat_B[1][4] +
                  mat_A[30][2] * mat_B[2][4] +
                  mat_A[30][3] * mat_B[3][4] +
                  mat_A[30][4] * mat_B[4][4] +
                  mat_A[30][5] * mat_B[5][4] +
                  mat_A[30][6] * mat_B[6][4] +
                  mat_A[30][7] * mat_B[7][4] +
                  mat_A[30][8] * mat_B[8][4] +
                  mat_A[30][9] * mat_B[9][4] +
                  mat_A[30][10] * mat_B[10][4] +
                  mat_A[30][11] * mat_B[11][4] +
                  mat_A[30][12] * mat_B[12][4] +
                  mat_A[30][13] * mat_B[13][4] +
                  mat_A[30][14] * mat_B[14][4] +
                  mat_A[30][15] * mat_B[15][4] +
                  mat_A[30][16] * mat_B[16][4] +
                  mat_A[30][17] * mat_B[17][4] +
                  mat_A[30][18] * mat_B[18][4] +
                  mat_A[30][19] * mat_B[19][4] +
                  mat_A[30][20] * mat_B[20][4] +
                  mat_A[30][21] * mat_B[21][4] +
                  mat_A[30][22] * mat_B[22][4] +
                  mat_A[30][23] * mat_B[23][4] +
                  mat_A[30][24] * mat_B[24][4] +
                  mat_A[30][25] * mat_B[25][4] +
                  mat_A[30][26] * mat_B[26][4] +
                  mat_A[30][27] * mat_B[27][4] +
                  mat_A[30][28] * mat_B[28][4] +
                  mat_A[30][29] * mat_B[29][4] +
                  mat_A[30][30] * mat_B[30][4] +
                  mat_A[30][31] * mat_B[31][4];
    mat_C[30][5] <= 
                  mat_A[30][0] * mat_B[0][5] +
                  mat_A[30][1] * mat_B[1][5] +
                  mat_A[30][2] * mat_B[2][5] +
                  mat_A[30][3] * mat_B[3][5] +
                  mat_A[30][4] * mat_B[4][5] +
                  mat_A[30][5] * mat_B[5][5] +
                  mat_A[30][6] * mat_B[6][5] +
                  mat_A[30][7] * mat_B[7][5] +
                  mat_A[30][8] * mat_B[8][5] +
                  mat_A[30][9] * mat_B[9][5] +
                  mat_A[30][10] * mat_B[10][5] +
                  mat_A[30][11] * mat_B[11][5] +
                  mat_A[30][12] * mat_B[12][5] +
                  mat_A[30][13] * mat_B[13][5] +
                  mat_A[30][14] * mat_B[14][5] +
                  mat_A[30][15] * mat_B[15][5] +
                  mat_A[30][16] * mat_B[16][5] +
                  mat_A[30][17] * mat_B[17][5] +
                  mat_A[30][18] * mat_B[18][5] +
                  mat_A[30][19] * mat_B[19][5] +
                  mat_A[30][20] * mat_B[20][5] +
                  mat_A[30][21] * mat_B[21][5] +
                  mat_A[30][22] * mat_B[22][5] +
                  mat_A[30][23] * mat_B[23][5] +
                  mat_A[30][24] * mat_B[24][5] +
                  mat_A[30][25] * mat_B[25][5] +
                  mat_A[30][26] * mat_B[26][5] +
                  mat_A[30][27] * mat_B[27][5] +
                  mat_A[30][28] * mat_B[28][5] +
                  mat_A[30][29] * mat_B[29][5] +
                  mat_A[30][30] * mat_B[30][5] +
                  mat_A[30][31] * mat_B[31][5];
    mat_C[30][6] <= 
                  mat_A[30][0] * mat_B[0][6] +
                  mat_A[30][1] * mat_B[1][6] +
                  mat_A[30][2] * mat_B[2][6] +
                  mat_A[30][3] * mat_B[3][6] +
                  mat_A[30][4] * mat_B[4][6] +
                  mat_A[30][5] * mat_B[5][6] +
                  mat_A[30][6] * mat_B[6][6] +
                  mat_A[30][7] * mat_B[7][6] +
                  mat_A[30][8] * mat_B[8][6] +
                  mat_A[30][9] * mat_B[9][6] +
                  mat_A[30][10] * mat_B[10][6] +
                  mat_A[30][11] * mat_B[11][6] +
                  mat_A[30][12] * mat_B[12][6] +
                  mat_A[30][13] * mat_B[13][6] +
                  mat_A[30][14] * mat_B[14][6] +
                  mat_A[30][15] * mat_B[15][6] +
                  mat_A[30][16] * mat_B[16][6] +
                  mat_A[30][17] * mat_B[17][6] +
                  mat_A[30][18] * mat_B[18][6] +
                  mat_A[30][19] * mat_B[19][6] +
                  mat_A[30][20] * mat_B[20][6] +
                  mat_A[30][21] * mat_B[21][6] +
                  mat_A[30][22] * mat_B[22][6] +
                  mat_A[30][23] * mat_B[23][6] +
                  mat_A[30][24] * mat_B[24][6] +
                  mat_A[30][25] * mat_B[25][6] +
                  mat_A[30][26] * mat_B[26][6] +
                  mat_A[30][27] * mat_B[27][6] +
                  mat_A[30][28] * mat_B[28][6] +
                  mat_A[30][29] * mat_B[29][6] +
                  mat_A[30][30] * mat_B[30][6] +
                  mat_A[30][31] * mat_B[31][6];
    mat_C[30][7] <= 
                  mat_A[30][0] * mat_B[0][7] +
                  mat_A[30][1] * mat_B[1][7] +
                  mat_A[30][2] * mat_B[2][7] +
                  mat_A[30][3] * mat_B[3][7] +
                  mat_A[30][4] * mat_B[4][7] +
                  mat_A[30][5] * mat_B[5][7] +
                  mat_A[30][6] * mat_B[6][7] +
                  mat_A[30][7] * mat_B[7][7] +
                  mat_A[30][8] * mat_B[8][7] +
                  mat_A[30][9] * mat_B[9][7] +
                  mat_A[30][10] * mat_B[10][7] +
                  mat_A[30][11] * mat_B[11][7] +
                  mat_A[30][12] * mat_B[12][7] +
                  mat_A[30][13] * mat_B[13][7] +
                  mat_A[30][14] * mat_B[14][7] +
                  mat_A[30][15] * mat_B[15][7] +
                  mat_A[30][16] * mat_B[16][7] +
                  mat_A[30][17] * mat_B[17][7] +
                  mat_A[30][18] * mat_B[18][7] +
                  mat_A[30][19] * mat_B[19][7] +
                  mat_A[30][20] * mat_B[20][7] +
                  mat_A[30][21] * mat_B[21][7] +
                  mat_A[30][22] * mat_B[22][7] +
                  mat_A[30][23] * mat_B[23][7] +
                  mat_A[30][24] * mat_B[24][7] +
                  mat_A[30][25] * mat_B[25][7] +
                  mat_A[30][26] * mat_B[26][7] +
                  mat_A[30][27] * mat_B[27][7] +
                  mat_A[30][28] * mat_B[28][7] +
                  mat_A[30][29] * mat_B[29][7] +
                  mat_A[30][30] * mat_B[30][7] +
                  mat_A[30][31] * mat_B[31][7];
    mat_C[30][8] <= 
                  mat_A[30][0] * mat_B[0][8] +
                  mat_A[30][1] * mat_B[1][8] +
                  mat_A[30][2] * mat_B[2][8] +
                  mat_A[30][3] * mat_B[3][8] +
                  mat_A[30][4] * mat_B[4][8] +
                  mat_A[30][5] * mat_B[5][8] +
                  mat_A[30][6] * mat_B[6][8] +
                  mat_A[30][7] * mat_B[7][8] +
                  mat_A[30][8] * mat_B[8][8] +
                  mat_A[30][9] * mat_B[9][8] +
                  mat_A[30][10] * mat_B[10][8] +
                  mat_A[30][11] * mat_B[11][8] +
                  mat_A[30][12] * mat_B[12][8] +
                  mat_A[30][13] * mat_B[13][8] +
                  mat_A[30][14] * mat_B[14][8] +
                  mat_A[30][15] * mat_B[15][8] +
                  mat_A[30][16] * mat_B[16][8] +
                  mat_A[30][17] * mat_B[17][8] +
                  mat_A[30][18] * mat_B[18][8] +
                  mat_A[30][19] * mat_B[19][8] +
                  mat_A[30][20] * mat_B[20][8] +
                  mat_A[30][21] * mat_B[21][8] +
                  mat_A[30][22] * mat_B[22][8] +
                  mat_A[30][23] * mat_B[23][8] +
                  mat_A[30][24] * mat_B[24][8] +
                  mat_A[30][25] * mat_B[25][8] +
                  mat_A[30][26] * mat_B[26][8] +
                  mat_A[30][27] * mat_B[27][8] +
                  mat_A[30][28] * mat_B[28][8] +
                  mat_A[30][29] * mat_B[29][8] +
                  mat_A[30][30] * mat_B[30][8] +
                  mat_A[30][31] * mat_B[31][8];
    mat_C[30][9] <= 
                  mat_A[30][0] * mat_B[0][9] +
                  mat_A[30][1] * mat_B[1][9] +
                  mat_A[30][2] * mat_B[2][9] +
                  mat_A[30][3] * mat_B[3][9] +
                  mat_A[30][4] * mat_B[4][9] +
                  mat_A[30][5] * mat_B[5][9] +
                  mat_A[30][6] * mat_B[6][9] +
                  mat_A[30][7] * mat_B[7][9] +
                  mat_A[30][8] * mat_B[8][9] +
                  mat_A[30][9] * mat_B[9][9] +
                  mat_A[30][10] * mat_B[10][9] +
                  mat_A[30][11] * mat_B[11][9] +
                  mat_A[30][12] * mat_B[12][9] +
                  mat_A[30][13] * mat_B[13][9] +
                  mat_A[30][14] * mat_B[14][9] +
                  mat_A[30][15] * mat_B[15][9] +
                  mat_A[30][16] * mat_B[16][9] +
                  mat_A[30][17] * mat_B[17][9] +
                  mat_A[30][18] * mat_B[18][9] +
                  mat_A[30][19] * mat_B[19][9] +
                  mat_A[30][20] * mat_B[20][9] +
                  mat_A[30][21] * mat_B[21][9] +
                  mat_A[30][22] * mat_B[22][9] +
                  mat_A[30][23] * mat_B[23][9] +
                  mat_A[30][24] * mat_B[24][9] +
                  mat_A[30][25] * mat_B[25][9] +
                  mat_A[30][26] * mat_B[26][9] +
                  mat_A[30][27] * mat_B[27][9] +
                  mat_A[30][28] * mat_B[28][9] +
                  mat_A[30][29] * mat_B[29][9] +
                  mat_A[30][30] * mat_B[30][9] +
                  mat_A[30][31] * mat_B[31][9];
    mat_C[30][10] <= 
                  mat_A[30][0] * mat_B[0][10] +
                  mat_A[30][1] * mat_B[1][10] +
                  mat_A[30][2] * mat_B[2][10] +
                  mat_A[30][3] * mat_B[3][10] +
                  mat_A[30][4] * mat_B[4][10] +
                  mat_A[30][5] * mat_B[5][10] +
                  mat_A[30][6] * mat_B[6][10] +
                  mat_A[30][7] * mat_B[7][10] +
                  mat_A[30][8] * mat_B[8][10] +
                  mat_A[30][9] * mat_B[9][10] +
                  mat_A[30][10] * mat_B[10][10] +
                  mat_A[30][11] * mat_B[11][10] +
                  mat_A[30][12] * mat_B[12][10] +
                  mat_A[30][13] * mat_B[13][10] +
                  mat_A[30][14] * mat_B[14][10] +
                  mat_A[30][15] * mat_B[15][10] +
                  mat_A[30][16] * mat_B[16][10] +
                  mat_A[30][17] * mat_B[17][10] +
                  mat_A[30][18] * mat_B[18][10] +
                  mat_A[30][19] * mat_B[19][10] +
                  mat_A[30][20] * mat_B[20][10] +
                  mat_A[30][21] * mat_B[21][10] +
                  mat_A[30][22] * mat_B[22][10] +
                  mat_A[30][23] * mat_B[23][10] +
                  mat_A[30][24] * mat_B[24][10] +
                  mat_A[30][25] * mat_B[25][10] +
                  mat_A[30][26] * mat_B[26][10] +
                  mat_A[30][27] * mat_B[27][10] +
                  mat_A[30][28] * mat_B[28][10] +
                  mat_A[30][29] * mat_B[29][10] +
                  mat_A[30][30] * mat_B[30][10] +
                  mat_A[30][31] * mat_B[31][10];
    mat_C[30][11] <= 
                  mat_A[30][0] * mat_B[0][11] +
                  mat_A[30][1] * mat_B[1][11] +
                  mat_A[30][2] * mat_B[2][11] +
                  mat_A[30][3] * mat_B[3][11] +
                  mat_A[30][4] * mat_B[4][11] +
                  mat_A[30][5] * mat_B[5][11] +
                  mat_A[30][6] * mat_B[6][11] +
                  mat_A[30][7] * mat_B[7][11] +
                  mat_A[30][8] * mat_B[8][11] +
                  mat_A[30][9] * mat_B[9][11] +
                  mat_A[30][10] * mat_B[10][11] +
                  mat_A[30][11] * mat_B[11][11] +
                  mat_A[30][12] * mat_B[12][11] +
                  mat_A[30][13] * mat_B[13][11] +
                  mat_A[30][14] * mat_B[14][11] +
                  mat_A[30][15] * mat_B[15][11] +
                  mat_A[30][16] * mat_B[16][11] +
                  mat_A[30][17] * mat_B[17][11] +
                  mat_A[30][18] * mat_B[18][11] +
                  mat_A[30][19] * mat_B[19][11] +
                  mat_A[30][20] * mat_B[20][11] +
                  mat_A[30][21] * mat_B[21][11] +
                  mat_A[30][22] * mat_B[22][11] +
                  mat_A[30][23] * mat_B[23][11] +
                  mat_A[30][24] * mat_B[24][11] +
                  mat_A[30][25] * mat_B[25][11] +
                  mat_A[30][26] * mat_B[26][11] +
                  mat_A[30][27] * mat_B[27][11] +
                  mat_A[30][28] * mat_B[28][11] +
                  mat_A[30][29] * mat_B[29][11] +
                  mat_A[30][30] * mat_B[30][11] +
                  mat_A[30][31] * mat_B[31][11];
    mat_C[30][12] <= 
                  mat_A[30][0] * mat_B[0][12] +
                  mat_A[30][1] * mat_B[1][12] +
                  mat_A[30][2] * mat_B[2][12] +
                  mat_A[30][3] * mat_B[3][12] +
                  mat_A[30][4] * mat_B[4][12] +
                  mat_A[30][5] * mat_B[5][12] +
                  mat_A[30][6] * mat_B[6][12] +
                  mat_A[30][7] * mat_B[7][12] +
                  mat_A[30][8] * mat_B[8][12] +
                  mat_A[30][9] * mat_B[9][12] +
                  mat_A[30][10] * mat_B[10][12] +
                  mat_A[30][11] * mat_B[11][12] +
                  mat_A[30][12] * mat_B[12][12] +
                  mat_A[30][13] * mat_B[13][12] +
                  mat_A[30][14] * mat_B[14][12] +
                  mat_A[30][15] * mat_B[15][12] +
                  mat_A[30][16] * mat_B[16][12] +
                  mat_A[30][17] * mat_B[17][12] +
                  mat_A[30][18] * mat_B[18][12] +
                  mat_A[30][19] * mat_B[19][12] +
                  mat_A[30][20] * mat_B[20][12] +
                  mat_A[30][21] * mat_B[21][12] +
                  mat_A[30][22] * mat_B[22][12] +
                  mat_A[30][23] * mat_B[23][12] +
                  mat_A[30][24] * mat_B[24][12] +
                  mat_A[30][25] * mat_B[25][12] +
                  mat_A[30][26] * mat_B[26][12] +
                  mat_A[30][27] * mat_B[27][12] +
                  mat_A[30][28] * mat_B[28][12] +
                  mat_A[30][29] * mat_B[29][12] +
                  mat_A[30][30] * mat_B[30][12] +
                  mat_A[30][31] * mat_B[31][12];
    mat_C[30][13] <= 
                  mat_A[30][0] * mat_B[0][13] +
                  mat_A[30][1] * mat_B[1][13] +
                  mat_A[30][2] * mat_B[2][13] +
                  mat_A[30][3] * mat_B[3][13] +
                  mat_A[30][4] * mat_B[4][13] +
                  mat_A[30][5] * mat_B[5][13] +
                  mat_A[30][6] * mat_B[6][13] +
                  mat_A[30][7] * mat_B[7][13] +
                  mat_A[30][8] * mat_B[8][13] +
                  mat_A[30][9] * mat_B[9][13] +
                  mat_A[30][10] * mat_B[10][13] +
                  mat_A[30][11] * mat_B[11][13] +
                  mat_A[30][12] * mat_B[12][13] +
                  mat_A[30][13] * mat_B[13][13] +
                  mat_A[30][14] * mat_B[14][13] +
                  mat_A[30][15] * mat_B[15][13] +
                  mat_A[30][16] * mat_B[16][13] +
                  mat_A[30][17] * mat_B[17][13] +
                  mat_A[30][18] * mat_B[18][13] +
                  mat_A[30][19] * mat_B[19][13] +
                  mat_A[30][20] * mat_B[20][13] +
                  mat_A[30][21] * mat_B[21][13] +
                  mat_A[30][22] * mat_B[22][13] +
                  mat_A[30][23] * mat_B[23][13] +
                  mat_A[30][24] * mat_B[24][13] +
                  mat_A[30][25] * mat_B[25][13] +
                  mat_A[30][26] * mat_B[26][13] +
                  mat_A[30][27] * mat_B[27][13] +
                  mat_A[30][28] * mat_B[28][13] +
                  mat_A[30][29] * mat_B[29][13] +
                  mat_A[30][30] * mat_B[30][13] +
                  mat_A[30][31] * mat_B[31][13];
    mat_C[30][14] <= 
                  mat_A[30][0] * mat_B[0][14] +
                  mat_A[30][1] * mat_B[1][14] +
                  mat_A[30][2] * mat_B[2][14] +
                  mat_A[30][3] * mat_B[3][14] +
                  mat_A[30][4] * mat_B[4][14] +
                  mat_A[30][5] * mat_B[5][14] +
                  mat_A[30][6] * mat_B[6][14] +
                  mat_A[30][7] * mat_B[7][14] +
                  mat_A[30][8] * mat_B[8][14] +
                  mat_A[30][9] * mat_B[9][14] +
                  mat_A[30][10] * mat_B[10][14] +
                  mat_A[30][11] * mat_B[11][14] +
                  mat_A[30][12] * mat_B[12][14] +
                  mat_A[30][13] * mat_B[13][14] +
                  mat_A[30][14] * mat_B[14][14] +
                  mat_A[30][15] * mat_B[15][14] +
                  mat_A[30][16] * mat_B[16][14] +
                  mat_A[30][17] * mat_B[17][14] +
                  mat_A[30][18] * mat_B[18][14] +
                  mat_A[30][19] * mat_B[19][14] +
                  mat_A[30][20] * mat_B[20][14] +
                  mat_A[30][21] * mat_B[21][14] +
                  mat_A[30][22] * mat_B[22][14] +
                  mat_A[30][23] * mat_B[23][14] +
                  mat_A[30][24] * mat_B[24][14] +
                  mat_A[30][25] * mat_B[25][14] +
                  mat_A[30][26] * mat_B[26][14] +
                  mat_A[30][27] * mat_B[27][14] +
                  mat_A[30][28] * mat_B[28][14] +
                  mat_A[30][29] * mat_B[29][14] +
                  mat_A[30][30] * mat_B[30][14] +
                  mat_A[30][31] * mat_B[31][14];
    mat_C[30][15] <= 
                  mat_A[30][0] * mat_B[0][15] +
                  mat_A[30][1] * mat_B[1][15] +
                  mat_A[30][2] * mat_B[2][15] +
                  mat_A[30][3] * mat_B[3][15] +
                  mat_A[30][4] * mat_B[4][15] +
                  mat_A[30][5] * mat_B[5][15] +
                  mat_A[30][6] * mat_B[6][15] +
                  mat_A[30][7] * mat_B[7][15] +
                  mat_A[30][8] * mat_B[8][15] +
                  mat_A[30][9] * mat_B[9][15] +
                  mat_A[30][10] * mat_B[10][15] +
                  mat_A[30][11] * mat_B[11][15] +
                  mat_A[30][12] * mat_B[12][15] +
                  mat_A[30][13] * mat_B[13][15] +
                  mat_A[30][14] * mat_B[14][15] +
                  mat_A[30][15] * mat_B[15][15] +
                  mat_A[30][16] * mat_B[16][15] +
                  mat_A[30][17] * mat_B[17][15] +
                  mat_A[30][18] * mat_B[18][15] +
                  mat_A[30][19] * mat_B[19][15] +
                  mat_A[30][20] * mat_B[20][15] +
                  mat_A[30][21] * mat_B[21][15] +
                  mat_A[30][22] * mat_B[22][15] +
                  mat_A[30][23] * mat_B[23][15] +
                  mat_A[30][24] * mat_B[24][15] +
                  mat_A[30][25] * mat_B[25][15] +
                  mat_A[30][26] * mat_B[26][15] +
                  mat_A[30][27] * mat_B[27][15] +
                  mat_A[30][28] * mat_B[28][15] +
                  mat_A[30][29] * mat_B[29][15] +
                  mat_A[30][30] * mat_B[30][15] +
                  mat_A[30][31] * mat_B[31][15];
    mat_C[30][16] <= 
                  mat_A[30][0] * mat_B[0][16] +
                  mat_A[30][1] * mat_B[1][16] +
                  mat_A[30][2] * mat_B[2][16] +
                  mat_A[30][3] * mat_B[3][16] +
                  mat_A[30][4] * mat_B[4][16] +
                  mat_A[30][5] * mat_B[5][16] +
                  mat_A[30][6] * mat_B[6][16] +
                  mat_A[30][7] * mat_B[7][16] +
                  mat_A[30][8] * mat_B[8][16] +
                  mat_A[30][9] * mat_B[9][16] +
                  mat_A[30][10] * mat_B[10][16] +
                  mat_A[30][11] * mat_B[11][16] +
                  mat_A[30][12] * mat_B[12][16] +
                  mat_A[30][13] * mat_B[13][16] +
                  mat_A[30][14] * mat_B[14][16] +
                  mat_A[30][15] * mat_B[15][16] +
                  mat_A[30][16] * mat_B[16][16] +
                  mat_A[30][17] * mat_B[17][16] +
                  mat_A[30][18] * mat_B[18][16] +
                  mat_A[30][19] * mat_B[19][16] +
                  mat_A[30][20] * mat_B[20][16] +
                  mat_A[30][21] * mat_B[21][16] +
                  mat_A[30][22] * mat_B[22][16] +
                  mat_A[30][23] * mat_B[23][16] +
                  mat_A[30][24] * mat_B[24][16] +
                  mat_A[30][25] * mat_B[25][16] +
                  mat_A[30][26] * mat_B[26][16] +
                  mat_A[30][27] * mat_B[27][16] +
                  mat_A[30][28] * mat_B[28][16] +
                  mat_A[30][29] * mat_B[29][16] +
                  mat_A[30][30] * mat_B[30][16] +
                  mat_A[30][31] * mat_B[31][16];
    mat_C[30][17] <= 
                  mat_A[30][0] * mat_B[0][17] +
                  mat_A[30][1] * mat_B[1][17] +
                  mat_A[30][2] * mat_B[2][17] +
                  mat_A[30][3] * mat_B[3][17] +
                  mat_A[30][4] * mat_B[4][17] +
                  mat_A[30][5] * mat_B[5][17] +
                  mat_A[30][6] * mat_B[6][17] +
                  mat_A[30][7] * mat_B[7][17] +
                  mat_A[30][8] * mat_B[8][17] +
                  mat_A[30][9] * mat_B[9][17] +
                  mat_A[30][10] * mat_B[10][17] +
                  mat_A[30][11] * mat_B[11][17] +
                  mat_A[30][12] * mat_B[12][17] +
                  mat_A[30][13] * mat_B[13][17] +
                  mat_A[30][14] * mat_B[14][17] +
                  mat_A[30][15] * mat_B[15][17] +
                  mat_A[30][16] * mat_B[16][17] +
                  mat_A[30][17] * mat_B[17][17] +
                  mat_A[30][18] * mat_B[18][17] +
                  mat_A[30][19] * mat_B[19][17] +
                  mat_A[30][20] * mat_B[20][17] +
                  mat_A[30][21] * mat_B[21][17] +
                  mat_A[30][22] * mat_B[22][17] +
                  mat_A[30][23] * mat_B[23][17] +
                  mat_A[30][24] * mat_B[24][17] +
                  mat_A[30][25] * mat_B[25][17] +
                  mat_A[30][26] * mat_B[26][17] +
                  mat_A[30][27] * mat_B[27][17] +
                  mat_A[30][28] * mat_B[28][17] +
                  mat_A[30][29] * mat_B[29][17] +
                  mat_A[30][30] * mat_B[30][17] +
                  mat_A[30][31] * mat_B[31][17];
    mat_C[30][18] <= 
                  mat_A[30][0] * mat_B[0][18] +
                  mat_A[30][1] * mat_B[1][18] +
                  mat_A[30][2] * mat_B[2][18] +
                  mat_A[30][3] * mat_B[3][18] +
                  mat_A[30][4] * mat_B[4][18] +
                  mat_A[30][5] * mat_B[5][18] +
                  mat_A[30][6] * mat_B[6][18] +
                  mat_A[30][7] * mat_B[7][18] +
                  mat_A[30][8] * mat_B[8][18] +
                  mat_A[30][9] * mat_B[9][18] +
                  mat_A[30][10] * mat_B[10][18] +
                  mat_A[30][11] * mat_B[11][18] +
                  mat_A[30][12] * mat_B[12][18] +
                  mat_A[30][13] * mat_B[13][18] +
                  mat_A[30][14] * mat_B[14][18] +
                  mat_A[30][15] * mat_B[15][18] +
                  mat_A[30][16] * mat_B[16][18] +
                  mat_A[30][17] * mat_B[17][18] +
                  mat_A[30][18] * mat_B[18][18] +
                  mat_A[30][19] * mat_B[19][18] +
                  mat_A[30][20] * mat_B[20][18] +
                  mat_A[30][21] * mat_B[21][18] +
                  mat_A[30][22] * mat_B[22][18] +
                  mat_A[30][23] * mat_B[23][18] +
                  mat_A[30][24] * mat_B[24][18] +
                  mat_A[30][25] * mat_B[25][18] +
                  mat_A[30][26] * mat_B[26][18] +
                  mat_A[30][27] * mat_B[27][18] +
                  mat_A[30][28] * mat_B[28][18] +
                  mat_A[30][29] * mat_B[29][18] +
                  mat_A[30][30] * mat_B[30][18] +
                  mat_A[30][31] * mat_B[31][18];
    mat_C[30][19] <= 
                  mat_A[30][0] * mat_B[0][19] +
                  mat_A[30][1] * mat_B[1][19] +
                  mat_A[30][2] * mat_B[2][19] +
                  mat_A[30][3] * mat_B[3][19] +
                  mat_A[30][4] * mat_B[4][19] +
                  mat_A[30][5] * mat_B[5][19] +
                  mat_A[30][6] * mat_B[6][19] +
                  mat_A[30][7] * mat_B[7][19] +
                  mat_A[30][8] * mat_B[8][19] +
                  mat_A[30][9] * mat_B[9][19] +
                  mat_A[30][10] * mat_B[10][19] +
                  mat_A[30][11] * mat_B[11][19] +
                  mat_A[30][12] * mat_B[12][19] +
                  mat_A[30][13] * mat_B[13][19] +
                  mat_A[30][14] * mat_B[14][19] +
                  mat_A[30][15] * mat_B[15][19] +
                  mat_A[30][16] * mat_B[16][19] +
                  mat_A[30][17] * mat_B[17][19] +
                  mat_A[30][18] * mat_B[18][19] +
                  mat_A[30][19] * mat_B[19][19] +
                  mat_A[30][20] * mat_B[20][19] +
                  mat_A[30][21] * mat_B[21][19] +
                  mat_A[30][22] * mat_B[22][19] +
                  mat_A[30][23] * mat_B[23][19] +
                  mat_A[30][24] * mat_B[24][19] +
                  mat_A[30][25] * mat_B[25][19] +
                  mat_A[30][26] * mat_B[26][19] +
                  mat_A[30][27] * mat_B[27][19] +
                  mat_A[30][28] * mat_B[28][19] +
                  mat_A[30][29] * mat_B[29][19] +
                  mat_A[30][30] * mat_B[30][19] +
                  mat_A[30][31] * mat_B[31][19];
    mat_C[30][20] <= 
                  mat_A[30][0] * mat_B[0][20] +
                  mat_A[30][1] * mat_B[1][20] +
                  mat_A[30][2] * mat_B[2][20] +
                  mat_A[30][3] * mat_B[3][20] +
                  mat_A[30][4] * mat_B[4][20] +
                  mat_A[30][5] * mat_B[5][20] +
                  mat_A[30][6] * mat_B[6][20] +
                  mat_A[30][7] * mat_B[7][20] +
                  mat_A[30][8] * mat_B[8][20] +
                  mat_A[30][9] * mat_B[9][20] +
                  mat_A[30][10] * mat_B[10][20] +
                  mat_A[30][11] * mat_B[11][20] +
                  mat_A[30][12] * mat_B[12][20] +
                  mat_A[30][13] * mat_B[13][20] +
                  mat_A[30][14] * mat_B[14][20] +
                  mat_A[30][15] * mat_B[15][20] +
                  mat_A[30][16] * mat_B[16][20] +
                  mat_A[30][17] * mat_B[17][20] +
                  mat_A[30][18] * mat_B[18][20] +
                  mat_A[30][19] * mat_B[19][20] +
                  mat_A[30][20] * mat_B[20][20] +
                  mat_A[30][21] * mat_B[21][20] +
                  mat_A[30][22] * mat_B[22][20] +
                  mat_A[30][23] * mat_B[23][20] +
                  mat_A[30][24] * mat_B[24][20] +
                  mat_A[30][25] * mat_B[25][20] +
                  mat_A[30][26] * mat_B[26][20] +
                  mat_A[30][27] * mat_B[27][20] +
                  mat_A[30][28] * mat_B[28][20] +
                  mat_A[30][29] * mat_B[29][20] +
                  mat_A[30][30] * mat_B[30][20] +
                  mat_A[30][31] * mat_B[31][20];
    mat_C[30][21] <= 
                  mat_A[30][0] * mat_B[0][21] +
                  mat_A[30][1] * mat_B[1][21] +
                  mat_A[30][2] * mat_B[2][21] +
                  mat_A[30][3] * mat_B[3][21] +
                  mat_A[30][4] * mat_B[4][21] +
                  mat_A[30][5] * mat_B[5][21] +
                  mat_A[30][6] * mat_B[6][21] +
                  mat_A[30][7] * mat_B[7][21] +
                  mat_A[30][8] * mat_B[8][21] +
                  mat_A[30][9] * mat_B[9][21] +
                  mat_A[30][10] * mat_B[10][21] +
                  mat_A[30][11] * mat_B[11][21] +
                  mat_A[30][12] * mat_B[12][21] +
                  mat_A[30][13] * mat_B[13][21] +
                  mat_A[30][14] * mat_B[14][21] +
                  mat_A[30][15] * mat_B[15][21] +
                  mat_A[30][16] * mat_B[16][21] +
                  mat_A[30][17] * mat_B[17][21] +
                  mat_A[30][18] * mat_B[18][21] +
                  mat_A[30][19] * mat_B[19][21] +
                  mat_A[30][20] * mat_B[20][21] +
                  mat_A[30][21] * mat_B[21][21] +
                  mat_A[30][22] * mat_B[22][21] +
                  mat_A[30][23] * mat_B[23][21] +
                  mat_A[30][24] * mat_B[24][21] +
                  mat_A[30][25] * mat_B[25][21] +
                  mat_A[30][26] * mat_B[26][21] +
                  mat_A[30][27] * mat_B[27][21] +
                  mat_A[30][28] * mat_B[28][21] +
                  mat_A[30][29] * mat_B[29][21] +
                  mat_A[30][30] * mat_B[30][21] +
                  mat_A[30][31] * mat_B[31][21];
    mat_C[30][22] <= 
                  mat_A[30][0] * mat_B[0][22] +
                  mat_A[30][1] * mat_B[1][22] +
                  mat_A[30][2] * mat_B[2][22] +
                  mat_A[30][3] * mat_B[3][22] +
                  mat_A[30][4] * mat_B[4][22] +
                  mat_A[30][5] * mat_B[5][22] +
                  mat_A[30][6] * mat_B[6][22] +
                  mat_A[30][7] * mat_B[7][22] +
                  mat_A[30][8] * mat_B[8][22] +
                  mat_A[30][9] * mat_B[9][22] +
                  mat_A[30][10] * mat_B[10][22] +
                  mat_A[30][11] * mat_B[11][22] +
                  mat_A[30][12] * mat_B[12][22] +
                  mat_A[30][13] * mat_B[13][22] +
                  mat_A[30][14] * mat_B[14][22] +
                  mat_A[30][15] * mat_B[15][22] +
                  mat_A[30][16] * mat_B[16][22] +
                  mat_A[30][17] * mat_B[17][22] +
                  mat_A[30][18] * mat_B[18][22] +
                  mat_A[30][19] * mat_B[19][22] +
                  mat_A[30][20] * mat_B[20][22] +
                  mat_A[30][21] * mat_B[21][22] +
                  mat_A[30][22] * mat_B[22][22] +
                  mat_A[30][23] * mat_B[23][22] +
                  mat_A[30][24] * mat_B[24][22] +
                  mat_A[30][25] * mat_B[25][22] +
                  mat_A[30][26] * mat_B[26][22] +
                  mat_A[30][27] * mat_B[27][22] +
                  mat_A[30][28] * mat_B[28][22] +
                  mat_A[30][29] * mat_B[29][22] +
                  mat_A[30][30] * mat_B[30][22] +
                  mat_A[30][31] * mat_B[31][22];
    mat_C[30][23] <= 
                  mat_A[30][0] * mat_B[0][23] +
                  mat_A[30][1] * mat_B[1][23] +
                  mat_A[30][2] * mat_B[2][23] +
                  mat_A[30][3] * mat_B[3][23] +
                  mat_A[30][4] * mat_B[4][23] +
                  mat_A[30][5] * mat_B[5][23] +
                  mat_A[30][6] * mat_B[6][23] +
                  mat_A[30][7] * mat_B[7][23] +
                  mat_A[30][8] * mat_B[8][23] +
                  mat_A[30][9] * mat_B[9][23] +
                  mat_A[30][10] * mat_B[10][23] +
                  mat_A[30][11] * mat_B[11][23] +
                  mat_A[30][12] * mat_B[12][23] +
                  mat_A[30][13] * mat_B[13][23] +
                  mat_A[30][14] * mat_B[14][23] +
                  mat_A[30][15] * mat_B[15][23] +
                  mat_A[30][16] * mat_B[16][23] +
                  mat_A[30][17] * mat_B[17][23] +
                  mat_A[30][18] * mat_B[18][23] +
                  mat_A[30][19] * mat_B[19][23] +
                  mat_A[30][20] * mat_B[20][23] +
                  mat_A[30][21] * mat_B[21][23] +
                  mat_A[30][22] * mat_B[22][23] +
                  mat_A[30][23] * mat_B[23][23] +
                  mat_A[30][24] * mat_B[24][23] +
                  mat_A[30][25] * mat_B[25][23] +
                  mat_A[30][26] * mat_B[26][23] +
                  mat_A[30][27] * mat_B[27][23] +
                  mat_A[30][28] * mat_B[28][23] +
                  mat_A[30][29] * mat_B[29][23] +
                  mat_A[30][30] * mat_B[30][23] +
                  mat_A[30][31] * mat_B[31][23];
    mat_C[30][24] <= 
                  mat_A[30][0] * mat_B[0][24] +
                  mat_A[30][1] * mat_B[1][24] +
                  mat_A[30][2] * mat_B[2][24] +
                  mat_A[30][3] * mat_B[3][24] +
                  mat_A[30][4] * mat_B[4][24] +
                  mat_A[30][5] * mat_B[5][24] +
                  mat_A[30][6] * mat_B[6][24] +
                  mat_A[30][7] * mat_B[7][24] +
                  mat_A[30][8] * mat_B[8][24] +
                  mat_A[30][9] * mat_B[9][24] +
                  mat_A[30][10] * mat_B[10][24] +
                  mat_A[30][11] * mat_B[11][24] +
                  mat_A[30][12] * mat_B[12][24] +
                  mat_A[30][13] * mat_B[13][24] +
                  mat_A[30][14] * mat_B[14][24] +
                  mat_A[30][15] * mat_B[15][24] +
                  mat_A[30][16] * mat_B[16][24] +
                  mat_A[30][17] * mat_B[17][24] +
                  mat_A[30][18] * mat_B[18][24] +
                  mat_A[30][19] * mat_B[19][24] +
                  mat_A[30][20] * mat_B[20][24] +
                  mat_A[30][21] * mat_B[21][24] +
                  mat_A[30][22] * mat_B[22][24] +
                  mat_A[30][23] * mat_B[23][24] +
                  mat_A[30][24] * mat_B[24][24] +
                  mat_A[30][25] * mat_B[25][24] +
                  mat_A[30][26] * mat_B[26][24] +
                  mat_A[30][27] * mat_B[27][24] +
                  mat_A[30][28] * mat_B[28][24] +
                  mat_A[30][29] * mat_B[29][24] +
                  mat_A[30][30] * mat_B[30][24] +
                  mat_A[30][31] * mat_B[31][24];
    mat_C[30][25] <= 
                  mat_A[30][0] * mat_B[0][25] +
                  mat_A[30][1] * mat_B[1][25] +
                  mat_A[30][2] * mat_B[2][25] +
                  mat_A[30][3] * mat_B[3][25] +
                  mat_A[30][4] * mat_B[4][25] +
                  mat_A[30][5] * mat_B[5][25] +
                  mat_A[30][6] * mat_B[6][25] +
                  mat_A[30][7] * mat_B[7][25] +
                  mat_A[30][8] * mat_B[8][25] +
                  mat_A[30][9] * mat_B[9][25] +
                  mat_A[30][10] * mat_B[10][25] +
                  mat_A[30][11] * mat_B[11][25] +
                  mat_A[30][12] * mat_B[12][25] +
                  mat_A[30][13] * mat_B[13][25] +
                  mat_A[30][14] * mat_B[14][25] +
                  mat_A[30][15] * mat_B[15][25] +
                  mat_A[30][16] * mat_B[16][25] +
                  mat_A[30][17] * mat_B[17][25] +
                  mat_A[30][18] * mat_B[18][25] +
                  mat_A[30][19] * mat_B[19][25] +
                  mat_A[30][20] * mat_B[20][25] +
                  mat_A[30][21] * mat_B[21][25] +
                  mat_A[30][22] * mat_B[22][25] +
                  mat_A[30][23] * mat_B[23][25] +
                  mat_A[30][24] * mat_B[24][25] +
                  mat_A[30][25] * mat_B[25][25] +
                  mat_A[30][26] * mat_B[26][25] +
                  mat_A[30][27] * mat_B[27][25] +
                  mat_A[30][28] * mat_B[28][25] +
                  mat_A[30][29] * mat_B[29][25] +
                  mat_A[30][30] * mat_B[30][25] +
                  mat_A[30][31] * mat_B[31][25];
    mat_C[30][26] <= 
                  mat_A[30][0] * mat_B[0][26] +
                  mat_A[30][1] * mat_B[1][26] +
                  mat_A[30][2] * mat_B[2][26] +
                  mat_A[30][3] * mat_B[3][26] +
                  mat_A[30][4] * mat_B[4][26] +
                  mat_A[30][5] * mat_B[5][26] +
                  mat_A[30][6] * mat_B[6][26] +
                  mat_A[30][7] * mat_B[7][26] +
                  mat_A[30][8] * mat_B[8][26] +
                  mat_A[30][9] * mat_B[9][26] +
                  mat_A[30][10] * mat_B[10][26] +
                  mat_A[30][11] * mat_B[11][26] +
                  mat_A[30][12] * mat_B[12][26] +
                  mat_A[30][13] * mat_B[13][26] +
                  mat_A[30][14] * mat_B[14][26] +
                  mat_A[30][15] * mat_B[15][26] +
                  mat_A[30][16] * mat_B[16][26] +
                  mat_A[30][17] * mat_B[17][26] +
                  mat_A[30][18] * mat_B[18][26] +
                  mat_A[30][19] * mat_B[19][26] +
                  mat_A[30][20] * mat_B[20][26] +
                  mat_A[30][21] * mat_B[21][26] +
                  mat_A[30][22] * mat_B[22][26] +
                  mat_A[30][23] * mat_B[23][26] +
                  mat_A[30][24] * mat_B[24][26] +
                  mat_A[30][25] * mat_B[25][26] +
                  mat_A[30][26] * mat_B[26][26] +
                  mat_A[30][27] * mat_B[27][26] +
                  mat_A[30][28] * mat_B[28][26] +
                  mat_A[30][29] * mat_B[29][26] +
                  mat_A[30][30] * mat_B[30][26] +
                  mat_A[30][31] * mat_B[31][26];
    mat_C[30][27] <= 
                  mat_A[30][0] * mat_B[0][27] +
                  mat_A[30][1] * mat_B[1][27] +
                  mat_A[30][2] * mat_B[2][27] +
                  mat_A[30][3] * mat_B[3][27] +
                  mat_A[30][4] * mat_B[4][27] +
                  mat_A[30][5] * mat_B[5][27] +
                  mat_A[30][6] * mat_B[6][27] +
                  mat_A[30][7] * mat_B[7][27] +
                  mat_A[30][8] * mat_B[8][27] +
                  mat_A[30][9] * mat_B[9][27] +
                  mat_A[30][10] * mat_B[10][27] +
                  mat_A[30][11] * mat_B[11][27] +
                  mat_A[30][12] * mat_B[12][27] +
                  mat_A[30][13] * mat_B[13][27] +
                  mat_A[30][14] * mat_B[14][27] +
                  mat_A[30][15] * mat_B[15][27] +
                  mat_A[30][16] * mat_B[16][27] +
                  mat_A[30][17] * mat_B[17][27] +
                  mat_A[30][18] * mat_B[18][27] +
                  mat_A[30][19] * mat_B[19][27] +
                  mat_A[30][20] * mat_B[20][27] +
                  mat_A[30][21] * mat_B[21][27] +
                  mat_A[30][22] * mat_B[22][27] +
                  mat_A[30][23] * mat_B[23][27] +
                  mat_A[30][24] * mat_B[24][27] +
                  mat_A[30][25] * mat_B[25][27] +
                  mat_A[30][26] * mat_B[26][27] +
                  mat_A[30][27] * mat_B[27][27] +
                  mat_A[30][28] * mat_B[28][27] +
                  mat_A[30][29] * mat_B[29][27] +
                  mat_A[30][30] * mat_B[30][27] +
                  mat_A[30][31] * mat_B[31][27];
    mat_C[30][28] <= 
                  mat_A[30][0] * mat_B[0][28] +
                  mat_A[30][1] * mat_B[1][28] +
                  mat_A[30][2] * mat_B[2][28] +
                  mat_A[30][3] * mat_B[3][28] +
                  mat_A[30][4] * mat_B[4][28] +
                  mat_A[30][5] * mat_B[5][28] +
                  mat_A[30][6] * mat_B[6][28] +
                  mat_A[30][7] * mat_B[7][28] +
                  mat_A[30][8] * mat_B[8][28] +
                  mat_A[30][9] * mat_B[9][28] +
                  mat_A[30][10] * mat_B[10][28] +
                  mat_A[30][11] * mat_B[11][28] +
                  mat_A[30][12] * mat_B[12][28] +
                  mat_A[30][13] * mat_B[13][28] +
                  mat_A[30][14] * mat_B[14][28] +
                  mat_A[30][15] * mat_B[15][28] +
                  mat_A[30][16] * mat_B[16][28] +
                  mat_A[30][17] * mat_B[17][28] +
                  mat_A[30][18] * mat_B[18][28] +
                  mat_A[30][19] * mat_B[19][28] +
                  mat_A[30][20] * mat_B[20][28] +
                  mat_A[30][21] * mat_B[21][28] +
                  mat_A[30][22] * mat_B[22][28] +
                  mat_A[30][23] * mat_B[23][28] +
                  mat_A[30][24] * mat_B[24][28] +
                  mat_A[30][25] * mat_B[25][28] +
                  mat_A[30][26] * mat_B[26][28] +
                  mat_A[30][27] * mat_B[27][28] +
                  mat_A[30][28] * mat_B[28][28] +
                  mat_A[30][29] * mat_B[29][28] +
                  mat_A[30][30] * mat_B[30][28] +
                  mat_A[30][31] * mat_B[31][28];
    mat_C[30][29] <= 
                  mat_A[30][0] * mat_B[0][29] +
                  mat_A[30][1] * mat_B[1][29] +
                  mat_A[30][2] * mat_B[2][29] +
                  mat_A[30][3] * mat_B[3][29] +
                  mat_A[30][4] * mat_B[4][29] +
                  mat_A[30][5] * mat_B[5][29] +
                  mat_A[30][6] * mat_B[6][29] +
                  mat_A[30][7] * mat_B[7][29] +
                  mat_A[30][8] * mat_B[8][29] +
                  mat_A[30][9] * mat_B[9][29] +
                  mat_A[30][10] * mat_B[10][29] +
                  mat_A[30][11] * mat_B[11][29] +
                  mat_A[30][12] * mat_B[12][29] +
                  mat_A[30][13] * mat_B[13][29] +
                  mat_A[30][14] * mat_B[14][29] +
                  mat_A[30][15] * mat_B[15][29] +
                  mat_A[30][16] * mat_B[16][29] +
                  mat_A[30][17] * mat_B[17][29] +
                  mat_A[30][18] * mat_B[18][29] +
                  mat_A[30][19] * mat_B[19][29] +
                  mat_A[30][20] * mat_B[20][29] +
                  mat_A[30][21] * mat_B[21][29] +
                  mat_A[30][22] * mat_B[22][29] +
                  mat_A[30][23] * mat_B[23][29] +
                  mat_A[30][24] * mat_B[24][29] +
                  mat_A[30][25] * mat_B[25][29] +
                  mat_A[30][26] * mat_B[26][29] +
                  mat_A[30][27] * mat_B[27][29] +
                  mat_A[30][28] * mat_B[28][29] +
                  mat_A[30][29] * mat_B[29][29] +
                  mat_A[30][30] * mat_B[30][29] +
                  mat_A[30][31] * mat_B[31][29];
    mat_C[30][30] <= 
                  mat_A[30][0] * mat_B[0][30] +
                  mat_A[30][1] * mat_B[1][30] +
                  mat_A[30][2] * mat_B[2][30] +
                  mat_A[30][3] * mat_B[3][30] +
                  mat_A[30][4] * mat_B[4][30] +
                  mat_A[30][5] * mat_B[5][30] +
                  mat_A[30][6] * mat_B[6][30] +
                  mat_A[30][7] * mat_B[7][30] +
                  mat_A[30][8] * mat_B[8][30] +
                  mat_A[30][9] * mat_B[9][30] +
                  mat_A[30][10] * mat_B[10][30] +
                  mat_A[30][11] * mat_B[11][30] +
                  mat_A[30][12] * mat_B[12][30] +
                  mat_A[30][13] * mat_B[13][30] +
                  mat_A[30][14] * mat_B[14][30] +
                  mat_A[30][15] * mat_B[15][30] +
                  mat_A[30][16] * mat_B[16][30] +
                  mat_A[30][17] * mat_B[17][30] +
                  mat_A[30][18] * mat_B[18][30] +
                  mat_A[30][19] * mat_B[19][30] +
                  mat_A[30][20] * mat_B[20][30] +
                  mat_A[30][21] * mat_B[21][30] +
                  mat_A[30][22] * mat_B[22][30] +
                  mat_A[30][23] * mat_B[23][30] +
                  mat_A[30][24] * mat_B[24][30] +
                  mat_A[30][25] * mat_B[25][30] +
                  mat_A[30][26] * mat_B[26][30] +
                  mat_A[30][27] * mat_B[27][30] +
                  mat_A[30][28] * mat_B[28][30] +
                  mat_A[30][29] * mat_B[29][30] +
                  mat_A[30][30] * mat_B[30][30] +
                  mat_A[30][31] * mat_B[31][30];
    mat_C[30][31] <= 
                  mat_A[30][0] * mat_B[0][31] +
                  mat_A[30][1] * mat_B[1][31] +
                  mat_A[30][2] * mat_B[2][31] +
                  mat_A[30][3] * mat_B[3][31] +
                  mat_A[30][4] * mat_B[4][31] +
                  mat_A[30][5] * mat_B[5][31] +
                  mat_A[30][6] * mat_B[6][31] +
                  mat_A[30][7] * mat_B[7][31] +
                  mat_A[30][8] * mat_B[8][31] +
                  mat_A[30][9] * mat_B[9][31] +
                  mat_A[30][10] * mat_B[10][31] +
                  mat_A[30][11] * mat_B[11][31] +
                  mat_A[30][12] * mat_B[12][31] +
                  mat_A[30][13] * mat_B[13][31] +
                  mat_A[30][14] * mat_B[14][31] +
                  mat_A[30][15] * mat_B[15][31] +
                  mat_A[30][16] * mat_B[16][31] +
                  mat_A[30][17] * mat_B[17][31] +
                  mat_A[30][18] * mat_B[18][31] +
                  mat_A[30][19] * mat_B[19][31] +
                  mat_A[30][20] * mat_B[20][31] +
                  mat_A[30][21] * mat_B[21][31] +
                  mat_A[30][22] * mat_B[22][31] +
                  mat_A[30][23] * mat_B[23][31] +
                  mat_A[30][24] * mat_B[24][31] +
                  mat_A[30][25] * mat_B[25][31] +
                  mat_A[30][26] * mat_B[26][31] +
                  mat_A[30][27] * mat_B[27][31] +
                  mat_A[30][28] * mat_B[28][31] +
                  mat_A[30][29] * mat_B[29][31] +
                  mat_A[30][30] * mat_B[30][31] +
                  mat_A[30][31] * mat_B[31][31];
    mat_C[31][0] <= 
                  mat_A[31][0] * mat_B[0][0] +
                  mat_A[31][1] * mat_B[1][0] +
                  mat_A[31][2] * mat_B[2][0] +
                  mat_A[31][3] * mat_B[3][0] +
                  mat_A[31][4] * mat_B[4][0] +
                  mat_A[31][5] * mat_B[5][0] +
                  mat_A[31][6] * mat_B[6][0] +
                  mat_A[31][7] * mat_B[7][0] +
                  mat_A[31][8] * mat_B[8][0] +
                  mat_A[31][9] * mat_B[9][0] +
                  mat_A[31][10] * mat_B[10][0] +
                  mat_A[31][11] * mat_B[11][0] +
                  mat_A[31][12] * mat_B[12][0] +
                  mat_A[31][13] * mat_B[13][0] +
                  mat_A[31][14] * mat_B[14][0] +
                  mat_A[31][15] * mat_B[15][0] +
                  mat_A[31][16] * mat_B[16][0] +
                  mat_A[31][17] * mat_B[17][0] +
                  mat_A[31][18] * mat_B[18][0] +
                  mat_A[31][19] * mat_B[19][0] +
                  mat_A[31][20] * mat_B[20][0] +
                  mat_A[31][21] * mat_B[21][0] +
                  mat_A[31][22] * mat_B[22][0] +
                  mat_A[31][23] * mat_B[23][0] +
                  mat_A[31][24] * mat_B[24][0] +
                  mat_A[31][25] * mat_B[25][0] +
                  mat_A[31][26] * mat_B[26][0] +
                  mat_A[31][27] * mat_B[27][0] +
                  mat_A[31][28] * mat_B[28][0] +
                  mat_A[31][29] * mat_B[29][0] +
                  mat_A[31][30] * mat_B[30][0] +
                  mat_A[31][31] * mat_B[31][0];
    mat_C[31][1] <= 
                  mat_A[31][0] * mat_B[0][1] +
                  mat_A[31][1] * mat_B[1][1] +
                  mat_A[31][2] * mat_B[2][1] +
                  mat_A[31][3] * mat_B[3][1] +
                  mat_A[31][4] * mat_B[4][1] +
                  mat_A[31][5] * mat_B[5][1] +
                  mat_A[31][6] * mat_B[6][1] +
                  mat_A[31][7] * mat_B[7][1] +
                  mat_A[31][8] * mat_B[8][1] +
                  mat_A[31][9] * mat_B[9][1] +
                  mat_A[31][10] * mat_B[10][1] +
                  mat_A[31][11] * mat_B[11][1] +
                  mat_A[31][12] * mat_B[12][1] +
                  mat_A[31][13] * mat_B[13][1] +
                  mat_A[31][14] * mat_B[14][1] +
                  mat_A[31][15] * mat_B[15][1] +
                  mat_A[31][16] * mat_B[16][1] +
                  mat_A[31][17] * mat_B[17][1] +
                  mat_A[31][18] * mat_B[18][1] +
                  mat_A[31][19] * mat_B[19][1] +
                  mat_A[31][20] * mat_B[20][1] +
                  mat_A[31][21] * mat_B[21][1] +
                  mat_A[31][22] * mat_B[22][1] +
                  mat_A[31][23] * mat_B[23][1] +
                  mat_A[31][24] * mat_B[24][1] +
                  mat_A[31][25] * mat_B[25][1] +
                  mat_A[31][26] * mat_B[26][1] +
                  mat_A[31][27] * mat_B[27][1] +
                  mat_A[31][28] * mat_B[28][1] +
                  mat_A[31][29] * mat_B[29][1] +
                  mat_A[31][30] * mat_B[30][1] +
                  mat_A[31][31] * mat_B[31][1];
    mat_C[31][2] <= 
                  mat_A[31][0] * mat_B[0][2] +
                  mat_A[31][1] * mat_B[1][2] +
                  mat_A[31][2] * mat_B[2][2] +
                  mat_A[31][3] * mat_B[3][2] +
                  mat_A[31][4] * mat_B[4][2] +
                  mat_A[31][5] * mat_B[5][2] +
                  mat_A[31][6] * mat_B[6][2] +
                  mat_A[31][7] * mat_B[7][2] +
                  mat_A[31][8] * mat_B[8][2] +
                  mat_A[31][9] * mat_B[9][2] +
                  mat_A[31][10] * mat_B[10][2] +
                  mat_A[31][11] * mat_B[11][2] +
                  mat_A[31][12] * mat_B[12][2] +
                  mat_A[31][13] * mat_B[13][2] +
                  mat_A[31][14] * mat_B[14][2] +
                  mat_A[31][15] * mat_B[15][2] +
                  mat_A[31][16] * mat_B[16][2] +
                  mat_A[31][17] * mat_B[17][2] +
                  mat_A[31][18] * mat_B[18][2] +
                  mat_A[31][19] * mat_B[19][2] +
                  mat_A[31][20] * mat_B[20][2] +
                  mat_A[31][21] * mat_B[21][2] +
                  mat_A[31][22] * mat_B[22][2] +
                  mat_A[31][23] * mat_B[23][2] +
                  mat_A[31][24] * mat_B[24][2] +
                  mat_A[31][25] * mat_B[25][2] +
                  mat_A[31][26] * mat_B[26][2] +
                  mat_A[31][27] * mat_B[27][2] +
                  mat_A[31][28] * mat_B[28][2] +
                  mat_A[31][29] * mat_B[29][2] +
                  mat_A[31][30] * mat_B[30][2] +
                  mat_A[31][31] * mat_B[31][2];
    mat_C[31][3] <= 
                  mat_A[31][0] * mat_B[0][3] +
                  mat_A[31][1] * mat_B[1][3] +
                  mat_A[31][2] * mat_B[2][3] +
                  mat_A[31][3] * mat_B[3][3] +
                  mat_A[31][4] * mat_B[4][3] +
                  mat_A[31][5] * mat_B[5][3] +
                  mat_A[31][6] * mat_B[6][3] +
                  mat_A[31][7] * mat_B[7][3] +
                  mat_A[31][8] * mat_B[8][3] +
                  mat_A[31][9] * mat_B[9][3] +
                  mat_A[31][10] * mat_B[10][3] +
                  mat_A[31][11] * mat_B[11][3] +
                  mat_A[31][12] * mat_B[12][3] +
                  mat_A[31][13] * mat_B[13][3] +
                  mat_A[31][14] * mat_B[14][3] +
                  mat_A[31][15] * mat_B[15][3] +
                  mat_A[31][16] * mat_B[16][3] +
                  mat_A[31][17] * mat_B[17][3] +
                  mat_A[31][18] * mat_B[18][3] +
                  mat_A[31][19] * mat_B[19][3] +
                  mat_A[31][20] * mat_B[20][3] +
                  mat_A[31][21] * mat_B[21][3] +
                  mat_A[31][22] * mat_B[22][3] +
                  mat_A[31][23] * mat_B[23][3] +
                  mat_A[31][24] * mat_B[24][3] +
                  mat_A[31][25] * mat_B[25][3] +
                  mat_A[31][26] * mat_B[26][3] +
                  mat_A[31][27] * mat_B[27][3] +
                  mat_A[31][28] * mat_B[28][3] +
                  mat_A[31][29] * mat_B[29][3] +
                  mat_A[31][30] * mat_B[30][3] +
                  mat_A[31][31] * mat_B[31][3];
    mat_C[31][4] <= 
                  mat_A[31][0] * mat_B[0][4] +
                  mat_A[31][1] * mat_B[1][4] +
                  mat_A[31][2] * mat_B[2][4] +
                  mat_A[31][3] * mat_B[3][4] +
                  mat_A[31][4] * mat_B[4][4] +
                  mat_A[31][5] * mat_B[5][4] +
                  mat_A[31][6] * mat_B[6][4] +
                  mat_A[31][7] * mat_B[7][4] +
                  mat_A[31][8] * mat_B[8][4] +
                  mat_A[31][9] * mat_B[9][4] +
                  mat_A[31][10] * mat_B[10][4] +
                  mat_A[31][11] * mat_B[11][4] +
                  mat_A[31][12] * mat_B[12][4] +
                  mat_A[31][13] * mat_B[13][4] +
                  mat_A[31][14] * mat_B[14][4] +
                  mat_A[31][15] * mat_B[15][4] +
                  mat_A[31][16] * mat_B[16][4] +
                  mat_A[31][17] * mat_B[17][4] +
                  mat_A[31][18] * mat_B[18][4] +
                  mat_A[31][19] * mat_B[19][4] +
                  mat_A[31][20] * mat_B[20][4] +
                  mat_A[31][21] * mat_B[21][4] +
                  mat_A[31][22] * mat_B[22][4] +
                  mat_A[31][23] * mat_B[23][4] +
                  mat_A[31][24] * mat_B[24][4] +
                  mat_A[31][25] * mat_B[25][4] +
                  mat_A[31][26] * mat_B[26][4] +
                  mat_A[31][27] * mat_B[27][4] +
                  mat_A[31][28] * mat_B[28][4] +
                  mat_A[31][29] * mat_B[29][4] +
                  mat_A[31][30] * mat_B[30][4] +
                  mat_A[31][31] * mat_B[31][4];
    mat_C[31][5] <= 
                  mat_A[31][0] * mat_B[0][5] +
                  mat_A[31][1] * mat_B[1][5] +
                  mat_A[31][2] * mat_B[2][5] +
                  mat_A[31][3] * mat_B[3][5] +
                  mat_A[31][4] * mat_B[4][5] +
                  mat_A[31][5] * mat_B[5][5] +
                  mat_A[31][6] * mat_B[6][5] +
                  mat_A[31][7] * mat_B[7][5] +
                  mat_A[31][8] * mat_B[8][5] +
                  mat_A[31][9] * mat_B[9][5] +
                  mat_A[31][10] * mat_B[10][5] +
                  mat_A[31][11] * mat_B[11][5] +
                  mat_A[31][12] * mat_B[12][5] +
                  mat_A[31][13] * mat_B[13][5] +
                  mat_A[31][14] * mat_B[14][5] +
                  mat_A[31][15] * mat_B[15][5] +
                  mat_A[31][16] * mat_B[16][5] +
                  mat_A[31][17] * mat_B[17][5] +
                  mat_A[31][18] * mat_B[18][5] +
                  mat_A[31][19] * mat_B[19][5] +
                  mat_A[31][20] * mat_B[20][5] +
                  mat_A[31][21] * mat_B[21][5] +
                  mat_A[31][22] * mat_B[22][5] +
                  mat_A[31][23] * mat_B[23][5] +
                  mat_A[31][24] * mat_B[24][5] +
                  mat_A[31][25] * mat_B[25][5] +
                  mat_A[31][26] * mat_B[26][5] +
                  mat_A[31][27] * mat_B[27][5] +
                  mat_A[31][28] * mat_B[28][5] +
                  mat_A[31][29] * mat_B[29][5] +
                  mat_A[31][30] * mat_B[30][5] +
                  mat_A[31][31] * mat_B[31][5];
    mat_C[31][6] <= 
                  mat_A[31][0] * mat_B[0][6] +
                  mat_A[31][1] * mat_B[1][6] +
                  mat_A[31][2] * mat_B[2][6] +
                  mat_A[31][3] * mat_B[3][6] +
                  mat_A[31][4] * mat_B[4][6] +
                  mat_A[31][5] * mat_B[5][6] +
                  mat_A[31][6] * mat_B[6][6] +
                  mat_A[31][7] * mat_B[7][6] +
                  mat_A[31][8] * mat_B[8][6] +
                  mat_A[31][9] * mat_B[9][6] +
                  mat_A[31][10] * mat_B[10][6] +
                  mat_A[31][11] * mat_B[11][6] +
                  mat_A[31][12] * mat_B[12][6] +
                  mat_A[31][13] * mat_B[13][6] +
                  mat_A[31][14] * mat_B[14][6] +
                  mat_A[31][15] * mat_B[15][6] +
                  mat_A[31][16] * mat_B[16][6] +
                  mat_A[31][17] * mat_B[17][6] +
                  mat_A[31][18] * mat_B[18][6] +
                  mat_A[31][19] * mat_B[19][6] +
                  mat_A[31][20] * mat_B[20][6] +
                  mat_A[31][21] * mat_B[21][6] +
                  mat_A[31][22] * mat_B[22][6] +
                  mat_A[31][23] * mat_B[23][6] +
                  mat_A[31][24] * mat_B[24][6] +
                  mat_A[31][25] * mat_B[25][6] +
                  mat_A[31][26] * mat_B[26][6] +
                  mat_A[31][27] * mat_B[27][6] +
                  mat_A[31][28] * mat_B[28][6] +
                  mat_A[31][29] * mat_B[29][6] +
                  mat_A[31][30] * mat_B[30][6] +
                  mat_A[31][31] * mat_B[31][6];
    mat_C[31][7] <= 
                  mat_A[31][0] * mat_B[0][7] +
                  mat_A[31][1] * mat_B[1][7] +
                  mat_A[31][2] * mat_B[2][7] +
                  mat_A[31][3] * mat_B[3][7] +
                  mat_A[31][4] * mat_B[4][7] +
                  mat_A[31][5] * mat_B[5][7] +
                  mat_A[31][6] * mat_B[6][7] +
                  mat_A[31][7] * mat_B[7][7] +
                  mat_A[31][8] * mat_B[8][7] +
                  mat_A[31][9] * mat_B[9][7] +
                  mat_A[31][10] * mat_B[10][7] +
                  mat_A[31][11] * mat_B[11][7] +
                  mat_A[31][12] * mat_B[12][7] +
                  mat_A[31][13] * mat_B[13][7] +
                  mat_A[31][14] * mat_B[14][7] +
                  mat_A[31][15] * mat_B[15][7] +
                  mat_A[31][16] * mat_B[16][7] +
                  mat_A[31][17] * mat_B[17][7] +
                  mat_A[31][18] * mat_B[18][7] +
                  mat_A[31][19] * mat_B[19][7] +
                  mat_A[31][20] * mat_B[20][7] +
                  mat_A[31][21] * mat_B[21][7] +
                  mat_A[31][22] * mat_B[22][7] +
                  mat_A[31][23] * mat_B[23][7] +
                  mat_A[31][24] * mat_B[24][7] +
                  mat_A[31][25] * mat_B[25][7] +
                  mat_A[31][26] * mat_B[26][7] +
                  mat_A[31][27] * mat_B[27][7] +
                  mat_A[31][28] * mat_B[28][7] +
                  mat_A[31][29] * mat_B[29][7] +
                  mat_A[31][30] * mat_B[30][7] +
                  mat_A[31][31] * mat_B[31][7];
    mat_C[31][8] <= 
                  mat_A[31][0] * mat_B[0][8] +
                  mat_A[31][1] * mat_B[1][8] +
                  mat_A[31][2] * mat_B[2][8] +
                  mat_A[31][3] * mat_B[3][8] +
                  mat_A[31][4] * mat_B[4][8] +
                  mat_A[31][5] * mat_B[5][8] +
                  mat_A[31][6] * mat_B[6][8] +
                  mat_A[31][7] * mat_B[7][8] +
                  mat_A[31][8] * mat_B[8][8] +
                  mat_A[31][9] * mat_B[9][8] +
                  mat_A[31][10] * mat_B[10][8] +
                  mat_A[31][11] * mat_B[11][8] +
                  mat_A[31][12] * mat_B[12][8] +
                  mat_A[31][13] * mat_B[13][8] +
                  mat_A[31][14] * mat_B[14][8] +
                  mat_A[31][15] * mat_B[15][8] +
                  mat_A[31][16] * mat_B[16][8] +
                  mat_A[31][17] * mat_B[17][8] +
                  mat_A[31][18] * mat_B[18][8] +
                  mat_A[31][19] * mat_B[19][8] +
                  mat_A[31][20] * mat_B[20][8] +
                  mat_A[31][21] * mat_B[21][8] +
                  mat_A[31][22] * mat_B[22][8] +
                  mat_A[31][23] * mat_B[23][8] +
                  mat_A[31][24] * mat_B[24][8] +
                  mat_A[31][25] * mat_B[25][8] +
                  mat_A[31][26] * mat_B[26][8] +
                  mat_A[31][27] * mat_B[27][8] +
                  mat_A[31][28] * mat_B[28][8] +
                  mat_A[31][29] * mat_B[29][8] +
                  mat_A[31][30] * mat_B[30][8] +
                  mat_A[31][31] * mat_B[31][8];
    mat_C[31][9] <= 
                  mat_A[31][0] * mat_B[0][9] +
                  mat_A[31][1] * mat_B[1][9] +
                  mat_A[31][2] * mat_B[2][9] +
                  mat_A[31][3] * mat_B[3][9] +
                  mat_A[31][4] * mat_B[4][9] +
                  mat_A[31][5] * mat_B[5][9] +
                  mat_A[31][6] * mat_B[6][9] +
                  mat_A[31][7] * mat_B[7][9] +
                  mat_A[31][8] * mat_B[8][9] +
                  mat_A[31][9] * mat_B[9][9] +
                  mat_A[31][10] * mat_B[10][9] +
                  mat_A[31][11] * mat_B[11][9] +
                  mat_A[31][12] * mat_B[12][9] +
                  mat_A[31][13] * mat_B[13][9] +
                  mat_A[31][14] * mat_B[14][9] +
                  mat_A[31][15] * mat_B[15][9] +
                  mat_A[31][16] * mat_B[16][9] +
                  mat_A[31][17] * mat_B[17][9] +
                  mat_A[31][18] * mat_B[18][9] +
                  mat_A[31][19] * mat_B[19][9] +
                  mat_A[31][20] * mat_B[20][9] +
                  mat_A[31][21] * mat_B[21][9] +
                  mat_A[31][22] * mat_B[22][9] +
                  mat_A[31][23] * mat_B[23][9] +
                  mat_A[31][24] * mat_B[24][9] +
                  mat_A[31][25] * mat_B[25][9] +
                  mat_A[31][26] * mat_B[26][9] +
                  mat_A[31][27] * mat_B[27][9] +
                  mat_A[31][28] * mat_B[28][9] +
                  mat_A[31][29] * mat_B[29][9] +
                  mat_A[31][30] * mat_B[30][9] +
                  mat_A[31][31] * mat_B[31][9];
    mat_C[31][10] <= 
                  mat_A[31][0] * mat_B[0][10] +
                  mat_A[31][1] * mat_B[1][10] +
                  mat_A[31][2] * mat_B[2][10] +
                  mat_A[31][3] * mat_B[3][10] +
                  mat_A[31][4] * mat_B[4][10] +
                  mat_A[31][5] * mat_B[5][10] +
                  mat_A[31][6] * mat_B[6][10] +
                  mat_A[31][7] * mat_B[7][10] +
                  mat_A[31][8] * mat_B[8][10] +
                  mat_A[31][9] * mat_B[9][10] +
                  mat_A[31][10] * mat_B[10][10] +
                  mat_A[31][11] * mat_B[11][10] +
                  mat_A[31][12] * mat_B[12][10] +
                  mat_A[31][13] * mat_B[13][10] +
                  mat_A[31][14] * mat_B[14][10] +
                  mat_A[31][15] * mat_B[15][10] +
                  mat_A[31][16] * mat_B[16][10] +
                  mat_A[31][17] * mat_B[17][10] +
                  mat_A[31][18] * mat_B[18][10] +
                  mat_A[31][19] * mat_B[19][10] +
                  mat_A[31][20] * mat_B[20][10] +
                  mat_A[31][21] * mat_B[21][10] +
                  mat_A[31][22] * mat_B[22][10] +
                  mat_A[31][23] * mat_B[23][10] +
                  mat_A[31][24] * mat_B[24][10] +
                  mat_A[31][25] * mat_B[25][10] +
                  mat_A[31][26] * mat_B[26][10] +
                  mat_A[31][27] * mat_B[27][10] +
                  mat_A[31][28] * mat_B[28][10] +
                  mat_A[31][29] * mat_B[29][10] +
                  mat_A[31][30] * mat_B[30][10] +
                  mat_A[31][31] * mat_B[31][10];
    mat_C[31][11] <= 
                  mat_A[31][0] * mat_B[0][11] +
                  mat_A[31][1] * mat_B[1][11] +
                  mat_A[31][2] * mat_B[2][11] +
                  mat_A[31][3] * mat_B[3][11] +
                  mat_A[31][4] * mat_B[4][11] +
                  mat_A[31][5] * mat_B[5][11] +
                  mat_A[31][6] * mat_B[6][11] +
                  mat_A[31][7] * mat_B[7][11] +
                  mat_A[31][8] * mat_B[8][11] +
                  mat_A[31][9] * mat_B[9][11] +
                  mat_A[31][10] * mat_B[10][11] +
                  mat_A[31][11] * mat_B[11][11] +
                  mat_A[31][12] * mat_B[12][11] +
                  mat_A[31][13] * mat_B[13][11] +
                  mat_A[31][14] * mat_B[14][11] +
                  mat_A[31][15] * mat_B[15][11] +
                  mat_A[31][16] * mat_B[16][11] +
                  mat_A[31][17] * mat_B[17][11] +
                  mat_A[31][18] * mat_B[18][11] +
                  mat_A[31][19] * mat_B[19][11] +
                  mat_A[31][20] * mat_B[20][11] +
                  mat_A[31][21] * mat_B[21][11] +
                  mat_A[31][22] * mat_B[22][11] +
                  mat_A[31][23] * mat_B[23][11] +
                  mat_A[31][24] * mat_B[24][11] +
                  mat_A[31][25] * mat_B[25][11] +
                  mat_A[31][26] * mat_B[26][11] +
                  mat_A[31][27] * mat_B[27][11] +
                  mat_A[31][28] * mat_B[28][11] +
                  mat_A[31][29] * mat_B[29][11] +
                  mat_A[31][30] * mat_B[30][11] +
                  mat_A[31][31] * mat_B[31][11];
    mat_C[31][12] <= 
                  mat_A[31][0] * mat_B[0][12] +
                  mat_A[31][1] * mat_B[1][12] +
                  mat_A[31][2] * mat_B[2][12] +
                  mat_A[31][3] * mat_B[3][12] +
                  mat_A[31][4] * mat_B[4][12] +
                  mat_A[31][5] * mat_B[5][12] +
                  mat_A[31][6] * mat_B[6][12] +
                  mat_A[31][7] * mat_B[7][12] +
                  mat_A[31][8] * mat_B[8][12] +
                  mat_A[31][9] * mat_B[9][12] +
                  mat_A[31][10] * mat_B[10][12] +
                  mat_A[31][11] * mat_B[11][12] +
                  mat_A[31][12] * mat_B[12][12] +
                  mat_A[31][13] * mat_B[13][12] +
                  mat_A[31][14] * mat_B[14][12] +
                  mat_A[31][15] * mat_B[15][12] +
                  mat_A[31][16] * mat_B[16][12] +
                  mat_A[31][17] * mat_B[17][12] +
                  mat_A[31][18] * mat_B[18][12] +
                  mat_A[31][19] * mat_B[19][12] +
                  mat_A[31][20] * mat_B[20][12] +
                  mat_A[31][21] * mat_B[21][12] +
                  mat_A[31][22] * mat_B[22][12] +
                  mat_A[31][23] * mat_B[23][12] +
                  mat_A[31][24] * mat_B[24][12] +
                  mat_A[31][25] * mat_B[25][12] +
                  mat_A[31][26] * mat_B[26][12] +
                  mat_A[31][27] * mat_B[27][12] +
                  mat_A[31][28] * mat_B[28][12] +
                  mat_A[31][29] * mat_B[29][12] +
                  mat_A[31][30] * mat_B[30][12] +
                  mat_A[31][31] * mat_B[31][12];
    mat_C[31][13] <= 
                  mat_A[31][0] * mat_B[0][13] +
                  mat_A[31][1] * mat_B[1][13] +
                  mat_A[31][2] * mat_B[2][13] +
                  mat_A[31][3] * mat_B[3][13] +
                  mat_A[31][4] * mat_B[4][13] +
                  mat_A[31][5] * mat_B[5][13] +
                  mat_A[31][6] * mat_B[6][13] +
                  mat_A[31][7] * mat_B[7][13] +
                  mat_A[31][8] * mat_B[8][13] +
                  mat_A[31][9] * mat_B[9][13] +
                  mat_A[31][10] * mat_B[10][13] +
                  mat_A[31][11] * mat_B[11][13] +
                  mat_A[31][12] * mat_B[12][13] +
                  mat_A[31][13] * mat_B[13][13] +
                  mat_A[31][14] * mat_B[14][13] +
                  mat_A[31][15] * mat_B[15][13] +
                  mat_A[31][16] * mat_B[16][13] +
                  mat_A[31][17] * mat_B[17][13] +
                  mat_A[31][18] * mat_B[18][13] +
                  mat_A[31][19] * mat_B[19][13] +
                  mat_A[31][20] * mat_B[20][13] +
                  mat_A[31][21] * mat_B[21][13] +
                  mat_A[31][22] * mat_B[22][13] +
                  mat_A[31][23] * mat_B[23][13] +
                  mat_A[31][24] * mat_B[24][13] +
                  mat_A[31][25] * mat_B[25][13] +
                  mat_A[31][26] * mat_B[26][13] +
                  mat_A[31][27] * mat_B[27][13] +
                  mat_A[31][28] * mat_B[28][13] +
                  mat_A[31][29] * mat_B[29][13] +
                  mat_A[31][30] * mat_B[30][13] +
                  mat_A[31][31] * mat_B[31][13];
    mat_C[31][14] <= 
                  mat_A[31][0] * mat_B[0][14] +
                  mat_A[31][1] * mat_B[1][14] +
                  mat_A[31][2] * mat_B[2][14] +
                  mat_A[31][3] * mat_B[3][14] +
                  mat_A[31][4] * mat_B[4][14] +
                  mat_A[31][5] * mat_B[5][14] +
                  mat_A[31][6] * mat_B[6][14] +
                  mat_A[31][7] * mat_B[7][14] +
                  mat_A[31][8] * mat_B[8][14] +
                  mat_A[31][9] * mat_B[9][14] +
                  mat_A[31][10] * mat_B[10][14] +
                  mat_A[31][11] * mat_B[11][14] +
                  mat_A[31][12] * mat_B[12][14] +
                  mat_A[31][13] * mat_B[13][14] +
                  mat_A[31][14] * mat_B[14][14] +
                  mat_A[31][15] * mat_B[15][14] +
                  mat_A[31][16] * mat_B[16][14] +
                  mat_A[31][17] * mat_B[17][14] +
                  mat_A[31][18] * mat_B[18][14] +
                  mat_A[31][19] * mat_B[19][14] +
                  mat_A[31][20] * mat_B[20][14] +
                  mat_A[31][21] * mat_B[21][14] +
                  mat_A[31][22] * mat_B[22][14] +
                  mat_A[31][23] * mat_B[23][14] +
                  mat_A[31][24] * mat_B[24][14] +
                  mat_A[31][25] * mat_B[25][14] +
                  mat_A[31][26] * mat_B[26][14] +
                  mat_A[31][27] * mat_B[27][14] +
                  mat_A[31][28] * mat_B[28][14] +
                  mat_A[31][29] * mat_B[29][14] +
                  mat_A[31][30] * mat_B[30][14] +
                  mat_A[31][31] * mat_B[31][14];
    mat_C[31][15] <= 
                  mat_A[31][0] * mat_B[0][15] +
                  mat_A[31][1] * mat_B[1][15] +
                  mat_A[31][2] * mat_B[2][15] +
                  mat_A[31][3] * mat_B[3][15] +
                  mat_A[31][4] * mat_B[4][15] +
                  mat_A[31][5] * mat_B[5][15] +
                  mat_A[31][6] * mat_B[6][15] +
                  mat_A[31][7] * mat_B[7][15] +
                  mat_A[31][8] * mat_B[8][15] +
                  mat_A[31][9] * mat_B[9][15] +
                  mat_A[31][10] * mat_B[10][15] +
                  mat_A[31][11] * mat_B[11][15] +
                  mat_A[31][12] * mat_B[12][15] +
                  mat_A[31][13] * mat_B[13][15] +
                  mat_A[31][14] * mat_B[14][15] +
                  mat_A[31][15] * mat_B[15][15] +
                  mat_A[31][16] * mat_B[16][15] +
                  mat_A[31][17] * mat_B[17][15] +
                  mat_A[31][18] * mat_B[18][15] +
                  mat_A[31][19] * mat_B[19][15] +
                  mat_A[31][20] * mat_B[20][15] +
                  mat_A[31][21] * mat_B[21][15] +
                  mat_A[31][22] * mat_B[22][15] +
                  mat_A[31][23] * mat_B[23][15] +
                  mat_A[31][24] * mat_B[24][15] +
                  mat_A[31][25] * mat_B[25][15] +
                  mat_A[31][26] * mat_B[26][15] +
                  mat_A[31][27] * mat_B[27][15] +
                  mat_A[31][28] * mat_B[28][15] +
                  mat_A[31][29] * mat_B[29][15] +
                  mat_A[31][30] * mat_B[30][15] +
                  mat_A[31][31] * mat_B[31][15];
    mat_C[31][16] <= 
                  mat_A[31][0] * mat_B[0][16] +
                  mat_A[31][1] * mat_B[1][16] +
                  mat_A[31][2] * mat_B[2][16] +
                  mat_A[31][3] * mat_B[3][16] +
                  mat_A[31][4] * mat_B[4][16] +
                  mat_A[31][5] * mat_B[5][16] +
                  mat_A[31][6] * mat_B[6][16] +
                  mat_A[31][7] * mat_B[7][16] +
                  mat_A[31][8] * mat_B[8][16] +
                  mat_A[31][9] * mat_B[9][16] +
                  mat_A[31][10] * mat_B[10][16] +
                  mat_A[31][11] * mat_B[11][16] +
                  mat_A[31][12] * mat_B[12][16] +
                  mat_A[31][13] * mat_B[13][16] +
                  mat_A[31][14] * mat_B[14][16] +
                  mat_A[31][15] * mat_B[15][16] +
                  mat_A[31][16] * mat_B[16][16] +
                  mat_A[31][17] * mat_B[17][16] +
                  mat_A[31][18] * mat_B[18][16] +
                  mat_A[31][19] * mat_B[19][16] +
                  mat_A[31][20] * mat_B[20][16] +
                  mat_A[31][21] * mat_B[21][16] +
                  mat_A[31][22] * mat_B[22][16] +
                  mat_A[31][23] * mat_B[23][16] +
                  mat_A[31][24] * mat_B[24][16] +
                  mat_A[31][25] * mat_B[25][16] +
                  mat_A[31][26] * mat_B[26][16] +
                  mat_A[31][27] * mat_B[27][16] +
                  mat_A[31][28] * mat_B[28][16] +
                  mat_A[31][29] * mat_B[29][16] +
                  mat_A[31][30] * mat_B[30][16] +
                  mat_A[31][31] * mat_B[31][16];
    mat_C[31][17] <= 
                  mat_A[31][0] * mat_B[0][17] +
                  mat_A[31][1] * mat_B[1][17] +
                  mat_A[31][2] * mat_B[2][17] +
                  mat_A[31][3] * mat_B[3][17] +
                  mat_A[31][4] * mat_B[4][17] +
                  mat_A[31][5] * mat_B[5][17] +
                  mat_A[31][6] * mat_B[6][17] +
                  mat_A[31][7] * mat_B[7][17] +
                  mat_A[31][8] * mat_B[8][17] +
                  mat_A[31][9] * mat_B[9][17] +
                  mat_A[31][10] * mat_B[10][17] +
                  mat_A[31][11] * mat_B[11][17] +
                  mat_A[31][12] * mat_B[12][17] +
                  mat_A[31][13] * mat_B[13][17] +
                  mat_A[31][14] * mat_B[14][17] +
                  mat_A[31][15] * mat_B[15][17] +
                  mat_A[31][16] * mat_B[16][17] +
                  mat_A[31][17] * mat_B[17][17] +
                  mat_A[31][18] * mat_B[18][17] +
                  mat_A[31][19] * mat_B[19][17] +
                  mat_A[31][20] * mat_B[20][17] +
                  mat_A[31][21] * mat_B[21][17] +
                  mat_A[31][22] * mat_B[22][17] +
                  mat_A[31][23] * mat_B[23][17] +
                  mat_A[31][24] * mat_B[24][17] +
                  mat_A[31][25] * mat_B[25][17] +
                  mat_A[31][26] * mat_B[26][17] +
                  mat_A[31][27] * mat_B[27][17] +
                  mat_A[31][28] * mat_B[28][17] +
                  mat_A[31][29] * mat_B[29][17] +
                  mat_A[31][30] * mat_B[30][17] +
                  mat_A[31][31] * mat_B[31][17];
    mat_C[31][18] <= 
                  mat_A[31][0] * mat_B[0][18] +
                  mat_A[31][1] * mat_B[1][18] +
                  mat_A[31][2] * mat_B[2][18] +
                  mat_A[31][3] * mat_B[3][18] +
                  mat_A[31][4] * mat_B[4][18] +
                  mat_A[31][5] * mat_B[5][18] +
                  mat_A[31][6] * mat_B[6][18] +
                  mat_A[31][7] * mat_B[7][18] +
                  mat_A[31][8] * mat_B[8][18] +
                  mat_A[31][9] * mat_B[9][18] +
                  mat_A[31][10] * mat_B[10][18] +
                  mat_A[31][11] * mat_B[11][18] +
                  mat_A[31][12] * mat_B[12][18] +
                  mat_A[31][13] * mat_B[13][18] +
                  mat_A[31][14] * mat_B[14][18] +
                  mat_A[31][15] * mat_B[15][18] +
                  mat_A[31][16] * mat_B[16][18] +
                  mat_A[31][17] * mat_B[17][18] +
                  mat_A[31][18] * mat_B[18][18] +
                  mat_A[31][19] * mat_B[19][18] +
                  mat_A[31][20] * mat_B[20][18] +
                  mat_A[31][21] * mat_B[21][18] +
                  mat_A[31][22] * mat_B[22][18] +
                  mat_A[31][23] * mat_B[23][18] +
                  mat_A[31][24] * mat_B[24][18] +
                  mat_A[31][25] * mat_B[25][18] +
                  mat_A[31][26] * mat_B[26][18] +
                  mat_A[31][27] * mat_B[27][18] +
                  mat_A[31][28] * mat_B[28][18] +
                  mat_A[31][29] * mat_B[29][18] +
                  mat_A[31][30] * mat_B[30][18] +
                  mat_A[31][31] * mat_B[31][18];
    mat_C[31][19] <= 
                  mat_A[31][0] * mat_B[0][19] +
                  mat_A[31][1] * mat_B[1][19] +
                  mat_A[31][2] * mat_B[2][19] +
                  mat_A[31][3] * mat_B[3][19] +
                  mat_A[31][4] * mat_B[4][19] +
                  mat_A[31][5] * mat_B[5][19] +
                  mat_A[31][6] * mat_B[6][19] +
                  mat_A[31][7] * mat_B[7][19] +
                  mat_A[31][8] * mat_B[8][19] +
                  mat_A[31][9] * mat_B[9][19] +
                  mat_A[31][10] * mat_B[10][19] +
                  mat_A[31][11] * mat_B[11][19] +
                  mat_A[31][12] * mat_B[12][19] +
                  mat_A[31][13] * mat_B[13][19] +
                  mat_A[31][14] * mat_B[14][19] +
                  mat_A[31][15] * mat_B[15][19] +
                  mat_A[31][16] * mat_B[16][19] +
                  mat_A[31][17] * mat_B[17][19] +
                  mat_A[31][18] * mat_B[18][19] +
                  mat_A[31][19] * mat_B[19][19] +
                  mat_A[31][20] * mat_B[20][19] +
                  mat_A[31][21] * mat_B[21][19] +
                  mat_A[31][22] * mat_B[22][19] +
                  mat_A[31][23] * mat_B[23][19] +
                  mat_A[31][24] * mat_B[24][19] +
                  mat_A[31][25] * mat_B[25][19] +
                  mat_A[31][26] * mat_B[26][19] +
                  mat_A[31][27] * mat_B[27][19] +
                  mat_A[31][28] * mat_B[28][19] +
                  mat_A[31][29] * mat_B[29][19] +
                  mat_A[31][30] * mat_B[30][19] +
                  mat_A[31][31] * mat_B[31][19];
    mat_C[31][20] <= 
                  mat_A[31][0] * mat_B[0][20] +
                  mat_A[31][1] * mat_B[1][20] +
                  mat_A[31][2] * mat_B[2][20] +
                  mat_A[31][3] * mat_B[3][20] +
                  mat_A[31][4] * mat_B[4][20] +
                  mat_A[31][5] * mat_B[5][20] +
                  mat_A[31][6] * mat_B[6][20] +
                  mat_A[31][7] * mat_B[7][20] +
                  mat_A[31][8] * mat_B[8][20] +
                  mat_A[31][9] * mat_B[9][20] +
                  mat_A[31][10] * mat_B[10][20] +
                  mat_A[31][11] * mat_B[11][20] +
                  mat_A[31][12] * mat_B[12][20] +
                  mat_A[31][13] * mat_B[13][20] +
                  mat_A[31][14] * mat_B[14][20] +
                  mat_A[31][15] * mat_B[15][20] +
                  mat_A[31][16] * mat_B[16][20] +
                  mat_A[31][17] * mat_B[17][20] +
                  mat_A[31][18] * mat_B[18][20] +
                  mat_A[31][19] * mat_B[19][20] +
                  mat_A[31][20] * mat_B[20][20] +
                  mat_A[31][21] * mat_B[21][20] +
                  mat_A[31][22] * mat_B[22][20] +
                  mat_A[31][23] * mat_B[23][20] +
                  mat_A[31][24] * mat_B[24][20] +
                  mat_A[31][25] * mat_B[25][20] +
                  mat_A[31][26] * mat_B[26][20] +
                  mat_A[31][27] * mat_B[27][20] +
                  mat_A[31][28] * mat_B[28][20] +
                  mat_A[31][29] * mat_B[29][20] +
                  mat_A[31][30] * mat_B[30][20] +
                  mat_A[31][31] * mat_B[31][20];
    mat_C[31][21] <= 
                  mat_A[31][0] * mat_B[0][21] +
                  mat_A[31][1] * mat_B[1][21] +
                  mat_A[31][2] * mat_B[2][21] +
                  mat_A[31][3] * mat_B[3][21] +
                  mat_A[31][4] * mat_B[4][21] +
                  mat_A[31][5] * mat_B[5][21] +
                  mat_A[31][6] * mat_B[6][21] +
                  mat_A[31][7] * mat_B[7][21] +
                  mat_A[31][8] * mat_B[8][21] +
                  mat_A[31][9] * mat_B[9][21] +
                  mat_A[31][10] * mat_B[10][21] +
                  mat_A[31][11] * mat_B[11][21] +
                  mat_A[31][12] * mat_B[12][21] +
                  mat_A[31][13] * mat_B[13][21] +
                  mat_A[31][14] * mat_B[14][21] +
                  mat_A[31][15] * mat_B[15][21] +
                  mat_A[31][16] * mat_B[16][21] +
                  mat_A[31][17] * mat_B[17][21] +
                  mat_A[31][18] * mat_B[18][21] +
                  mat_A[31][19] * mat_B[19][21] +
                  mat_A[31][20] * mat_B[20][21] +
                  mat_A[31][21] * mat_B[21][21] +
                  mat_A[31][22] * mat_B[22][21] +
                  mat_A[31][23] * mat_B[23][21] +
                  mat_A[31][24] * mat_B[24][21] +
                  mat_A[31][25] * mat_B[25][21] +
                  mat_A[31][26] * mat_B[26][21] +
                  mat_A[31][27] * mat_B[27][21] +
                  mat_A[31][28] * mat_B[28][21] +
                  mat_A[31][29] * mat_B[29][21] +
                  mat_A[31][30] * mat_B[30][21] +
                  mat_A[31][31] * mat_B[31][21];
    mat_C[31][22] <= 
                  mat_A[31][0] * mat_B[0][22] +
                  mat_A[31][1] * mat_B[1][22] +
                  mat_A[31][2] * mat_B[2][22] +
                  mat_A[31][3] * mat_B[3][22] +
                  mat_A[31][4] * mat_B[4][22] +
                  mat_A[31][5] * mat_B[5][22] +
                  mat_A[31][6] * mat_B[6][22] +
                  mat_A[31][7] * mat_B[7][22] +
                  mat_A[31][8] * mat_B[8][22] +
                  mat_A[31][9] * mat_B[9][22] +
                  mat_A[31][10] * mat_B[10][22] +
                  mat_A[31][11] * mat_B[11][22] +
                  mat_A[31][12] * mat_B[12][22] +
                  mat_A[31][13] * mat_B[13][22] +
                  mat_A[31][14] * mat_B[14][22] +
                  mat_A[31][15] * mat_B[15][22] +
                  mat_A[31][16] * mat_B[16][22] +
                  mat_A[31][17] * mat_B[17][22] +
                  mat_A[31][18] * mat_B[18][22] +
                  mat_A[31][19] * mat_B[19][22] +
                  mat_A[31][20] * mat_B[20][22] +
                  mat_A[31][21] * mat_B[21][22] +
                  mat_A[31][22] * mat_B[22][22] +
                  mat_A[31][23] * mat_B[23][22] +
                  mat_A[31][24] * mat_B[24][22] +
                  mat_A[31][25] * mat_B[25][22] +
                  mat_A[31][26] * mat_B[26][22] +
                  mat_A[31][27] * mat_B[27][22] +
                  mat_A[31][28] * mat_B[28][22] +
                  mat_A[31][29] * mat_B[29][22] +
                  mat_A[31][30] * mat_B[30][22] +
                  mat_A[31][31] * mat_B[31][22];
    mat_C[31][23] <= 
                  mat_A[31][0] * mat_B[0][23] +
                  mat_A[31][1] * mat_B[1][23] +
                  mat_A[31][2] * mat_B[2][23] +
                  mat_A[31][3] * mat_B[3][23] +
                  mat_A[31][4] * mat_B[4][23] +
                  mat_A[31][5] * mat_B[5][23] +
                  mat_A[31][6] * mat_B[6][23] +
                  mat_A[31][7] * mat_B[7][23] +
                  mat_A[31][8] * mat_B[8][23] +
                  mat_A[31][9] * mat_B[9][23] +
                  mat_A[31][10] * mat_B[10][23] +
                  mat_A[31][11] * mat_B[11][23] +
                  mat_A[31][12] * mat_B[12][23] +
                  mat_A[31][13] * mat_B[13][23] +
                  mat_A[31][14] * mat_B[14][23] +
                  mat_A[31][15] * mat_B[15][23] +
                  mat_A[31][16] * mat_B[16][23] +
                  mat_A[31][17] * mat_B[17][23] +
                  mat_A[31][18] * mat_B[18][23] +
                  mat_A[31][19] * mat_B[19][23] +
                  mat_A[31][20] * mat_B[20][23] +
                  mat_A[31][21] * mat_B[21][23] +
                  mat_A[31][22] * mat_B[22][23] +
                  mat_A[31][23] * mat_B[23][23] +
                  mat_A[31][24] * mat_B[24][23] +
                  mat_A[31][25] * mat_B[25][23] +
                  mat_A[31][26] * mat_B[26][23] +
                  mat_A[31][27] * mat_B[27][23] +
                  mat_A[31][28] * mat_B[28][23] +
                  mat_A[31][29] * mat_B[29][23] +
                  mat_A[31][30] * mat_B[30][23] +
                  mat_A[31][31] * mat_B[31][23];
    mat_C[31][24] <= 
                  mat_A[31][0] * mat_B[0][24] +
                  mat_A[31][1] * mat_B[1][24] +
                  mat_A[31][2] * mat_B[2][24] +
                  mat_A[31][3] * mat_B[3][24] +
                  mat_A[31][4] * mat_B[4][24] +
                  mat_A[31][5] * mat_B[5][24] +
                  mat_A[31][6] * mat_B[6][24] +
                  mat_A[31][7] * mat_B[7][24] +
                  mat_A[31][8] * mat_B[8][24] +
                  mat_A[31][9] * mat_B[9][24] +
                  mat_A[31][10] * mat_B[10][24] +
                  mat_A[31][11] * mat_B[11][24] +
                  mat_A[31][12] * mat_B[12][24] +
                  mat_A[31][13] * mat_B[13][24] +
                  mat_A[31][14] * mat_B[14][24] +
                  mat_A[31][15] * mat_B[15][24] +
                  mat_A[31][16] * mat_B[16][24] +
                  mat_A[31][17] * mat_B[17][24] +
                  mat_A[31][18] * mat_B[18][24] +
                  mat_A[31][19] * mat_B[19][24] +
                  mat_A[31][20] * mat_B[20][24] +
                  mat_A[31][21] * mat_B[21][24] +
                  mat_A[31][22] * mat_B[22][24] +
                  mat_A[31][23] * mat_B[23][24] +
                  mat_A[31][24] * mat_B[24][24] +
                  mat_A[31][25] * mat_B[25][24] +
                  mat_A[31][26] * mat_B[26][24] +
                  mat_A[31][27] * mat_B[27][24] +
                  mat_A[31][28] * mat_B[28][24] +
                  mat_A[31][29] * mat_B[29][24] +
                  mat_A[31][30] * mat_B[30][24] +
                  mat_A[31][31] * mat_B[31][24];
    mat_C[31][25] <= 
                  mat_A[31][0] * mat_B[0][25] +
                  mat_A[31][1] * mat_B[1][25] +
                  mat_A[31][2] * mat_B[2][25] +
                  mat_A[31][3] * mat_B[3][25] +
                  mat_A[31][4] * mat_B[4][25] +
                  mat_A[31][5] * mat_B[5][25] +
                  mat_A[31][6] * mat_B[6][25] +
                  mat_A[31][7] * mat_B[7][25] +
                  mat_A[31][8] * mat_B[8][25] +
                  mat_A[31][9] * mat_B[9][25] +
                  mat_A[31][10] * mat_B[10][25] +
                  mat_A[31][11] * mat_B[11][25] +
                  mat_A[31][12] * mat_B[12][25] +
                  mat_A[31][13] * mat_B[13][25] +
                  mat_A[31][14] * mat_B[14][25] +
                  mat_A[31][15] * mat_B[15][25] +
                  mat_A[31][16] * mat_B[16][25] +
                  mat_A[31][17] * mat_B[17][25] +
                  mat_A[31][18] * mat_B[18][25] +
                  mat_A[31][19] * mat_B[19][25] +
                  mat_A[31][20] * mat_B[20][25] +
                  mat_A[31][21] * mat_B[21][25] +
                  mat_A[31][22] * mat_B[22][25] +
                  mat_A[31][23] * mat_B[23][25] +
                  mat_A[31][24] * mat_B[24][25] +
                  mat_A[31][25] * mat_B[25][25] +
                  mat_A[31][26] * mat_B[26][25] +
                  mat_A[31][27] * mat_B[27][25] +
                  mat_A[31][28] * mat_B[28][25] +
                  mat_A[31][29] * mat_B[29][25] +
                  mat_A[31][30] * mat_B[30][25] +
                  mat_A[31][31] * mat_B[31][25];
    mat_C[31][26] <= 
                  mat_A[31][0] * mat_B[0][26] +
                  mat_A[31][1] * mat_B[1][26] +
                  mat_A[31][2] * mat_B[2][26] +
                  mat_A[31][3] * mat_B[3][26] +
                  mat_A[31][4] * mat_B[4][26] +
                  mat_A[31][5] * mat_B[5][26] +
                  mat_A[31][6] * mat_B[6][26] +
                  mat_A[31][7] * mat_B[7][26] +
                  mat_A[31][8] * mat_B[8][26] +
                  mat_A[31][9] * mat_B[9][26] +
                  mat_A[31][10] * mat_B[10][26] +
                  mat_A[31][11] * mat_B[11][26] +
                  mat_A[31][12] * mat_B[12][26] +
                  mat_A[31][13] * mat_B[13][26] +
                  mat_A[31][14] * mat_B[14][26] +
                  mat_A[31][15] * mat_B[15][26] +
                  mat_A[31][16] * mat_B[16][26] +
                  mat_A[31][17] * mat_B[17][26] +
                  mat_A[31][18] * mat_B[18][26] +
                  mat_A[31][19] * mat_B[19][26] +
                  mat_A[31][20] * mat_B[20][26] +
                  mat_A[31][21] * mat_B[21][26] +
                  mat_A[31][22] * mat_B[22][26] +
                  mat_A[31][23] * mat_B[23][26] +
                  mat_A[31][24] * mat_B[24][26] +
                  mat_A[31][25] * mat_B[25][26] +
                  mat_A[31][26] * mat_B[26][26] +
                  mat_A[31][27] * mat_B[27][26] +
                  mat_A[31][28] * mat_B[28][26] +
                  mat_A[31][29] * mat_B[29][26] +
                  mat_A[31][30] * mat_B[30][26] +
                  mat_A[31][31] * mat_B[31][26];
    mat_C[31][27] <= 
                  mat_A[31][0] * mat_B[0][27] +
                  mat_A[31][1] * mat_B[1][27] +
                  mat_A[31][2] * mat_B[2][27] +
                  mat_A[31][3] * mat_B[3][27] +
                  mat_A[31][4] * mat_B[4][27] +
                  mat_A[31][5] * mat_B[5][27] +
                  mat_A[31][6] * mat_B[6][27] +
                  mat_A[31][7] * mat_B[7][27] +
                  mat_A[31][8] * mat_B[8][27] +
                  mat_A[31][9] * mat_B[9][27] +
                  mat_A[31][10] * mat_B[10][27] +
                  mat_A[31][11] * mat_B[11][27] +
                  mat_A[31][12] * mat_B[12][27] +
                  mat_A[31][13] * mat_B[13][27] +
                  mat_A[31][14] * mat_B[14][27] +
                  mat_A[31][15] * mat_B[15][27] +
                  mat_A[31][16] * mat_B[16][27] +
                  mat_A[31][17] * mat_B[17][27] +
                  mat_A[31][18] * mat_B[18][27] +
                  mat_A[31][19] * mat_B[19][27] +
                  mat_A[31][20] * mat_B[20][27] +
                  mat_A[31][21] * mat_B[21][27] +
                  mat_A[31][22] * mat_B[22][27] +
                  mat_A[31][23] * mat_B[23][27] +
                  mat_A[31][24] * mat_B[24][27] +
                  mat_A[31][25] * mat_B[25][27] +
                  mat_A[31][26] * mat_B[26][27] +
                  mat_A[31][27] * mat_B[27][27] +
                  mat_A[31][28] * mat_B[28][27] +
                  mat_A[31][29] * mat_B[29][27] +
                  mat_A[31][30] * mat_B[30][27] +
                  mat_A[31][31] * mat_B[31][27];
    mat_C[31][28] <= 
                  mat_A[31][0] * mat_B[0][28] +
                  mat_A[31][1] * mat_B[1][28] +
                  mat_A[31][2] * mat_B[2][28] +
                  mat_A[31][3] * mat_B[3][28] +
                  mat_A[31][4] * mat_B[4][28] +
                  mat_A[31][5] * mat_B[5][28] +
                  mat_A[31][6] * mat_B[6][28] +
                  mat_A[31][7] * mat_B[7][28] +
                  mat_A[31][8] * mat_B[8][28] +
                  mat_A[31][9] * mat_B[9][28] +
                  mat_A[31][10] * mat_B[10][28] +
                  mat_A[31][11] * mat_B[11][28] +
                  mat_A[31][12] * mat_B[12][28] +
                  mat_A[31][13] * mat_B[13][28] +
                  mat_A[31][14] * mat_B[14][28] +
                  mat_A[31][15] * mat_B[15][28] +
                  mat_A[31][16] * mat_B[16][28] +
                  mat_A[31][17] * mat_B[17][28] +
                  mat_A[31][18] * mat_B[18][28] +
                  mat_A[31][19] * mat_B[19][28] +
                  mat_A[31][20] * mat_B[20][28] +
                  mat_A[31][21] * mat_B[21][28] +
                  mat_A[31][22] * mat_B[22][28] +
                  mat_A[31][23] * mat_B[23][28] +
                  mat_A[31][24] * mat_B[24][28] +
                  mat_A[31][25] * mat_B[25][28] +
                  mat_A[31][26] * mat_B[26][28] +
                  mat_A[31][27] * mat_B[27][28] +
                  mat_A[31][28] * mat_B[28][28] +
                  mat_A[31][29] * mat_B[29][28] +
                  mat_A[31][30] * mat_B[30][28] +
                  mat_A[31][31] * mat_B[31][28];
    mat_C[31][29] <= 
                  mat_A[31][0] * mat_B[0][29] +
                  mat_A[31][1] * mat_B[1][29] +
                  mat_A[31][2] * mat_B[2][29] +
                  mat_A[31][3] * mat_B[3][29] +
                  mat_A[31][4] * mat_B[4][29] +
                  mat_A[31][5] * mat_B[5][29] +
                  mat_A[31][6] * mat_B[6][29] +
                  mat_A[31][7] * mat_B[7][29] +
                  mat_A[31][8] * mat_B[8][29] +
                  mat_A[31][9] * mat_B[9][29] +
                  mat_A[31][10] * mat_B[10][29] +
                  mat_A[31][11] * mat_B[11][29] +
                  mat_A[31][12] * mat_B[12][29] +
                  mat_A[31][13] * mat_B[13][29] +
                  mat_A[31][14] * mat_B[14][29] +
                  mat_A[31][15] * mat_B[15][29] +
                  mat_A[31][16] * mat_B[16][29] +
                  mat_A[31][17] * mat_B[17][29] +
                  mat_A[31][18] * mat_B[18][29] +
                  mat_A[31][19] * mat_B[19][29] +
                  mat_A[31][20] * mat_B[20][29] +
                  mat_A[31][21] * mat_B[21][29] +
                  mat_A[31][22] * mat_B[22][29] +
                  mat_A[31][23] * mat_B[23][29] +
                  mat_A[31][24] * mat_B[24][29] +
                  mat_A[31][25] * mat_B[25][29] +
                  mat_A[31][26] * mat_B[26][29] +
                  mat_A[31][27] * mat_B[27][29] +
                  mat_A[31][28] * mat_B[28][29] +
                  mat_A[31][29] * mat_B[29][29] +
                  mat_A[31][30] * mat_B[30][29] +
                  mat_A[31][31] * mat_B[31][29];
    mat_C[31][30] <= 
                  mat_A[31][0] * mat_B[0][30] +
                  mat_A[31][1] * mat_B[1][30] +
                  mat_A[31][2] * mat_B[2][30] +
                  mat_A[31][3] * mat_B[3][30] +
                  mat_A[31][4] * mat_B[4][30] +
                  mat_A[31][5] * mat_B[5][30] +
                  mat_A[31][6] * mat_B[6][30] +
                  mat_A[31][7] * mat_B[7][30] +
                  mat_A[31][8] * mat_B[8][30] +
                  mat_A[31][9] * mat_B[9][30] +
                  mat_A[31][10] * mat_B[10][30] +
                  mat_A[31][11] * mat_B[11][30] +
                  mat_A[31][12] * mat_B[12][30] +
                  mat_A[31][13] * mat_B[13][30] +
                  mat_A[31][14] * mat_B[14][30] +
                  mat_A[31][15] * mat_B[15][30] +
                  mat_A[31][16] * mat_B[16][30] +
                  mat_A[31][17] * mat_B[17][30] +
                  mat_A[31][18] * mat_B[18][30] +
                  mat_A[31][19] * mat_B[19][30] +
                  mat_A[31][20] * mat_B[20][30] +
                  mat_A[31][21] * mat_B[21][30] +
                  mat_A[31][22] * mat_B[22][30] +
                  mat_A[31][23] * mat_B[23][30] +
                  mat_A[31][24] * mat_B[24][30] +
                  mat_A[31][25] * mat_B[25][30] +
                  mat_A[31][26] * mat_B[26][30] +
                  mat_A[31][27] * mat_B[27][30] +
                  mat_A[31][28] * mat_B[28][30] +
                  mat_A[31][29] * mat_B[29][30] +
                  mat_A[31][30] * mat_B[30][30] +
                  mat_A[31][31] * mat_B[31][30];
    mat_C[31][31] <= 
                  mat_A[31][0] * mat_B[0][31] +
                  mat_A[31][1] * mat_B[1][31] +
                  mat_A[31][2] * mat_B[2][31] +
                  mat_A[31][3] * mat_B[3][31] +
                  mat_A[31][4] * mat_B[4][31] +
                  mat_A[31][5] * mat_B[5][31] +
                  mat_A[31][6] * mat_B[6][31] +
                  mat_A[31][7] * mat_B[7][31] +
                  mat_A[31][8] * mat_B[8][31] +
                  mat_A[31][9] * mat_B[9][31] +
                  mat_A[31][10] * mat_B[10][31] +
                  mat_A[31][11] * mat_B[11][31] +
                  mat_A[31][12] * mat_B[12][31] +
                  mat_A[31][13] * mat_B[13][31] +
                  mat_A[31][14] * mat_B[14][31] +
                  mat_A[31][15] * mat_B[15][31] +
                  mat_A[31][16] * mat_B[16][31] +
                  mat_A[31][17] * mat_B[17][31] +
                  mat_A[31][18] * mat_B[18][31] +
                  mat_A[31][19] * mat_B[19][31] +
                  mat_A[31][20] * mat_B[20][31] +
                  mat_A[31][21] * mat_B[21][31] +
                  mat_A[31][22] * mat_B[22][31] +
                  mat_A[31][23] * mat_B[23][31] +
                  mat_A[31][24] * mat_B[24][31] +
                  mat_A[31][25] * mat_B[25][31] +
                  mat_A[31][26] * mat_B[26][31] +
                  mat_A[31][27] * mat_B[27][31] +
                  mat_A[31][28] * mat_B[28][31] +
                  mat_A[31][29] * mat_B[29][31] +
                  mat_A[31][30] * mat_B[30][31] +
                  mat_A[31][31] * mat_B[31][31];
                    end
endmodule
