module multiply_long #(
  parameter mat_size = 2,
  parameter dat_size = 8
) (
  input  logic            start        ,
  input  logic            clk          , //kanske ej behövs
  input  logic [3:0][7:0] mat_A [255:0],
  input  logic [3:0][7:0] mat_B [255:0],
  output logic [3:0][7:0] mat_C [255:0],
  output logic            done
);

  always @(posedge clk)
  begin
    mat_C[0][0] <=
                mat_A[0][0] * mat_B[0][0] +
                mat_A[0][1] * mat_B[8][0] +
                mat_A[0][2] * mat_B[16][0] +
                mat_A[0][3] * mat_B[24][0] +
                mat_A[1][0] * mat_B[32][0] +
                mat_A[1][1] * mat_B[40][0] +
                mat_A[1][2] * mat_B[48][0] +
                mat_A[1][3] * mat_B[56][0] +
                mat_A[2][0] * mat_B[64][0] +
                mat_A[2][1] * mat_B[72][0] +
                mat_A[2][2] * mat_B[80][0] +
                mat_A[2][3] * mat_B[88][0] +
                mat_A[3][0] * mat_B[96][0] +
                mat_A[3][1] * mat_B[104][0] +
                mat_A[3][2] * mat_B[112][0] +
                mat_A[3][3] * mat_B[120][0] +
                mat_A[4][0] * mat_B[128][0] +
                mat_A[4][1] * mat_B[136][0] +
                mat_A[4][2] * mat_B[144][0] +
                mat_A[4][3] * mat_B[152][0] +
                mat_A[5][0] * mat_B[160][0] +
                mat_A[5][1] * mat_B[168][0] +
                mat_A[5][2] * mat_B[176][0] +
                mat_A[5][3] * mat_B[184][0] +
                mat_A[6][0] * mat_B[192][0] +
                mat_A[6][1] * mat_B[200][0] +
                mat_A[6][2] * mat_B[208][0] +
                mat_A[6][3] * mat_B[216][0] +
                mat_A[7][0] * mat_B[224][0] +
                mat_A[7][1] * mat_B[232][0] +
                mat_A[7][2] * mat_B[240][0] +
                mat_A[7][3] * mat_B[248][0];
    mat_C[0][1] <=
                mat_A[0][0] * mat_B[0][1] +
                mat_A[0][1] * mat_B[8][1] +
                mat_A[0][2] * mat_B[16][1] +
                mat_A[0][3] * mat_B[24][1] +
                mat_A[1][0] * mat_B[32][1] +
                mat_A[1][1] * mat_B[40][1] +
                mat_A[1][2] * mat_B[48][1] +
                mat_A[1][3] * mat_B[56][1] +
                mat_A[2][0] * mat_B[64][1] +
                mat_A[2][1] * mat_B[72][1] +
                mat_A[2][2] * mat_B[80][1] +
                mat_A[2][3] * mat_B[88][1] +
                mat_A[3][0] * mat_B[96][1] +
                mat_A[3][1] * mat_B[104][1] +
                mat_A[3][2] * mat_B[112][1] +
                mat_A[3][3] * mat_B[120][1] +
                mat_A[4][0] * mat_B[128][1] +
                mat_A[4][1] * mat_B[136][1] +
                mat_A[4][2] * mat_B[144][1] +
                mat_A[4][3] * mat_B[152][1] +
                mat_A[5][0] * mat_B[160][1] +
                mat_A[5][1] * mat_B[168][1] +
                mat_A[5][2] * mat_B[176][1] +
                mat_A[5][3] * mat_B[184][1] +
                mat_A[6][0] * mat_B[192][1] +
                mat_A[6][1] * mat_B[200][1] +
                mat_A[6][2] * mat_B[208][1] +
                mat_A[6][3] * mat_B[216][1] +
                mat_A[7][0] * mat_B[224][1] +
                mat_A[7][1] * mat_B[232][1] +
                mat_A[7][2] * mat_B[240][1] +
                mat_A[7][3] * mat_B[248][1];
    mat_C[0][2] <=
                mat_A[0][0] * mat_B[0][2] +
                mat_A[0][1] * mat_B[8][2] +
                mat_A[0][2] * mat_B[16][2] +
                mat_A[0][3] * mat_B[24][2] +
                mat_A[1][0] * mat_B[32][2] +
                mat_A[1][1] * mat_B[40][2] +
                mat_A[1][2] * mat_B[48][2] +
                mat_A[1][3] * mat_B[56][2] +
                mat_A[2][0] * mat_B[64][2] +
                mat_A[2][1] * mat_B[72][2] +
                mat_A[2][2] * mat_B[80][2] +
                mat_A[2][3] * mat_B[88][2] +
                mat_A[3][0] * mat_B[96][2] +
                mat_A[3][1] * mat_B[104][2] +
                mat_A[3][2] * mat_B[112][2] +
                mat_A[3][3] * mat_B[120][2] +
                mat_A[4][0] * mat_B[128][2] +
                mat_A[4][1] * mat_B[136][2] +
                mat_A[4][2] * mat_B[144][2] +
                mat_A[4][3] * mat_B[152][2] +
                mat_A[5][0] * mat_B[160][2] +
                mat_A[5][1] * mat_B[168][2] +
                mat_A[5][2] * mat_B[176][2] +
                mat_A[5][3] * mat_B[184][2] +
                mat_A[6][0] * mat_B[192][2] +
                mat_A[6][1] * mat_B[200][2] +
                mat_A[6][2] * mat_B[208][2] +
                mat_A[6][3] * mat_B[216][2] +
                mat_A[7][0] * mat_B[224][2] +
                mat_A[7][1] * mat_B[232][2] +
                mat_A[7][2] * mat_B[240][2] +
                mat_A[7][3] * mat_B[248][2];
    mat_C[0][3] <=
                mat_A[0][0] * mat_B[0][3] +
                mat_A[0][1] * mat_B[8][3] +
                mat_A[0][2] * mat_B[16][3] +
                mat_A[0][3] * mat_B[24][3] +
                mat_A[1][0] * mat_B[32][3] +
                mat_A[1][1] * mat_B[40][3] +
                mat_A[1][2] * mat_B[48][3] +
                mat_A[1][3] * mat_B[56][3] +
                mat_A[2][0] * mat_B[64][3] +
                mat_A[2][1] * mat_B[72][3] +
                mat_A[2][2] * mat_B[80][3] +
                mat_A[2][3] * mat_B[88][3] +
                mat_A[3][0] * mat_B[96][3] +
                mat_A[3][1] * mat_B[104][3] +
                mat_A[3][2] * mat_B[112][3] +
                mat_A[3][3] * mat_B[120][3] +
                mat_A[4][0] * mat_B[128][3] +
                mat_A[4][1] * mat_B[136][3] +
                mat_A[4][2] * mat_B[144][3] +
                mat_A[4][3] * mat_B[152][3] +
                mat_A[5][0] * mat_B[160][3] +
                mat_A[5][1] * mat_B[168][3] +
                mat_A[5][2] * mat_B[176][3] +
                mat_A[5][3] * mat_B[184][3] +
                mat_A[6][0] * mat_B[192][3] +
                mat_A[6][1] * mat_B[200][3] +
                mat_A[6][2] * mat_B[208][3] +
                mat_A[6][3] * mat_B[216][3] +
                mat_A[7][0] * mat_B[224][3] +
                mat_A[7][1] * mat_B[232][3] +
                mat_A[7][2] * mat_B[240][3] +
                mat_A[7][3] * mat_B[248][3];
    mat_C[1][0] <=
                mat_A[0][0] * mat_B[1][0] +
                mat_A[0][1] * mat_B[9][0] +
                mat_A[0][2] * mat_B[17][0] +
                mat_A[0][3] * mat_B[25][0] +
                mat_A[1][0] * mat_B[33][0] +
                mat_A[1][1] * mat_B[41][0] +
                mat_A[1][2] * mat_B[49][0] +
                mat_A[1][3] * mat_B[57][0] +
                mat_A[2][0] * mat_B[65][0] +
                mat_A[2][1] * mat_B[73][0] +
                mat_A[2][2] * mat_B[81][0] +
                mat_A[2][3] * mat_B[89][0] +
                mat_A[3][0] * mat_B[97][0] +
                mat_A[3][1] * mat_B[105][0] +
                mat_A[3][2] * mat_B[113][0] +
                mat_A[3][3] * mat_B[121][0] +
                mat_A[4][0] * mat_B[129][0] +
                mat_A[4][1] * mat_B[137][0] +
                mat_A[4][2] * mat_B[145][0] +
                mat_A[4][3] * mat_B[153][0] +
                mat_A[5][0] * mat_B[161][0] +
                mat_A[5][1] * mat_B[169][0] +
                mat_A[5][2] * mat_B[177][0] +
                mat_A[5][3] * mat_B[185][0] +
                mat_A[6][0] * mat_B[193][0] +
                mat_A[6][1] * mat_B[201][0] +
                mat_A[6][2] * mat_B[209][0] +
                mat_A[6][3] * mat_B[217][0] +
                mat_A[7][0] * mat_B[225][0] +
                mat_A[7][1] * mat_B[233][0] +
                mat_A[7][2] * mat_B[241][0] +
                mat_A[7][3] * mat_B[249][0];
    mat_C[1][1] <=
                mat_A[0][0] * mat_B[1][1] +
                mat_A[0][1] * mat_B[9][1] +
                mat_A[0][2] * mat_B[17][1] +
                mat_A[0][3] * mat_B[25][1] +
                mat_A[1][0] * mat_B[33][1] +
                mat_A[1][1] * mat_B[41][1] +
                mat_A[1][2] * mat_B[49][1] +
                mat_A[1][3] * mat_B[57][1] +
                mat_A[2][0] * mat_B[65][1] +
                mat_A[2][1] * mat_B[73][1] +
                mat_A[2][2] * mat_B[81][1] +
                mat_A[2][3] * mat_B[89][1] +
                mat_A[3][0] * mat_B[97][1] +
                mat_A[3][1] * mat_B[105][1] +
                mat_A[3][2] * mat_B[113][1] +
                mat_A[3][3] * mat_B[121][1] +
                mat_A[4][0] * mat_B[129][1] +
                mat_A[4][1] * mat_B[137][1] +
                mat_A[4][2] * mat_B[145][1] +
                mat_A[4][3] * mat_B[153][1] +
                mat_A[5][0] * mat_B[161][1] +
                mat_A[5][1] * mat_B[169][1] +
                mat_A[5][2] * mat_B[177][1] +
                mat_A[5][3] * mat_B[185][1] +
                mat_A[6][0] * mat_B[193][1] +
                mat_A[6][1] * mat_B[201][1] +
                mat_A[6][2] * mat_B[209][1] +
                mat_A[6][3] * mat_B[217][1] +
                mat_A[7][0] * mat_B[225][1] +
                mat_A[7][1] * mat_B[233][1] +
                mat_A[7][2] * mat_B[241][1] +
                mat_A[7][3] * mat_B[249][1];
    mat_C[1][2] <=
                mat_A[0][0] * mat_B[1][2] +
                mat_A[0][1] * mat_B[9][2] +
                mat_A[0][2] * mat_B[17][2] +
                mat_A[0][3] * mat_B[25][2] +
                mat_A[1][0] * mat_B[33][2] +
                mat_A[1][1] * mat_B[41][2] +
                mat_A[1][2] * mat_B[49][2] +
                mat_A[1][3] * mat_B[57][2] +
                mat_A[2][0] * mat_B[65][2] +
                mat_A[2][1] * mat_B[73][2] +
                mat_A[2][2] * mat_B[81][2] +
                mat_A[2][3] * mat_B[89][2] +
                mat_A[3][0] * mat_B[97][2] +
                mat_A[3][1] * mat_B[105][2] +
                mat_A[3][2] * mat_B[113][2] +
                mat_A[3][3] * mat_B[121][2] +
                mat_A[4][0] * mat_B[129][2] +
                mat_A[4][1] * mat_B[137][2] +
                mat_A[4][2] * mat_B[145][2] +
                mat_A[4][3] * mat_B[153][2] +
                mat_A[5][0] * mat_B[161][2] +
                mat_A[5][1] * mat_B[169][2] +
                mat_A[5][2] * mat_B[177][2] +
                mat_A[5][3] * mat_B[185][2] +
                mat_A[6][0] * mat_B[193][2] +
                mat_A[6][1] * mat_B[201][2] +
                mat_A[6][2] * mat_B[209][2] +
                mat_A[6][3] * mat_B[217][2] +
                mat_A[7][0] * mat_B[225][2] +
                mat_A[7][1] * mat_B[233][2] +
                mat_A[7][2] * mat_B[241][2] +
                mat_A[7][3] * mat_B[249][2];
    mat_C[1][3] <=
                mat_A[0][0] * mat_B[1][3] +
                mat_A[0][1] * mat_B[9][3] +
                mat_A[0][2] * mat_B[17][3] +
                mat_A[0][3] * mat_B[25][3] +
                mat_A[1][0] * mat_B[33][3] +
                mat_A[1][1] * mat_B[41][3] +
                mat_A[1][2] * mat_B[49][3] +
                mat_A[1][3] * mat_B[57][3] +
                mat_A[2][0] * mat_B[65][3] +
                mat_A[2][1] * mat_B[73][3] +
                mat_A[2][2] * mat_B[81][3] +
                mat_A[2][3] * mat_B[89][3] +
                mat_A[3][0] * mat_B[97][3] +
                mat_A[3][1] * mat_B[105][3] +
                mat_A[3][2] * mat_B[113][3] +
                mat_A[3][3] * mat_B[121][3] +
                mat_A[4][0] * mat_B[129][3] +
                mat_A[4][1] * mat_B[137][3] +
                mat_A[4][2] * mat_B[145][3] +
                mat_A[4][3] * mat_B[153][3] +
                mat_A[5][0] * mat_B[161][3] +
                mat_A[5][1] * mat_B[169][3] +
                mat_A[5][2] * mat_B[177][3] +
                mat_A[5][3] * mat_B[185][3] +
                mat_A[6][0] * mat_B[193][3] +
                mat_A[6][1] * mat_B[201][3] +
                mat_A[6][2] * mat_B[209][3] +
                mat_A[6][3] * mat_B[217][3] +
                mat_A[7][0] * mat_B[225][3] +
                mat_A[7][1] * mat_B[233][3] +
                mat_A[7][2] * mat_B[241][3] +
                mat_A[7][3] * mat_B[249][3];
    mat_C[2][0] <=
                mat_A[0][0] * mat_B[2][0] +
                mat_A[0][1] * mat_B[10][0] +
                mat_A[0][2] * mat_B[18][0] +
                mat_A[0][3] * mat_B[26][0] +
                mat_A[1][0] * mat_B[34][0] +
                mat_A[1][1] * mat_B[42][0] +
                mat_A[1][2] * mat_B[50][0] +
                mat_A[1][3] * mat_B[58][0] +
                mat_A[2][0] * mat_B[66][0] +
                mat_A[2][1] * mat_B[74][0] +
                mat_A[2][2] * mat_B[82][0] +
                mat_A[2][3] * mat_B[90][0] +
                mat_A[3][0] * mat_B[98][0] +
                mat_A[3][1] * mat_B[106][0] +
                mat_A[3][2] * mat_B[114][0] +
                mat_A[3][3] * mat_B[122][0] +
                mat_A[4][0] * mat_B[130][0] +
                mat_A[4][1] * mat_B[138][0] +
                mat_A[4][2] * mat_B[146][0] +
                mat_A[4][3] * mat_B[154][0] +
                mat_A[5][0] * mat_B[162][0] +
                mat_A[5][1] * mat_B[170][0] +
                mat_A[5][2] * mat_B[178][0] +
                mat_A[5][3] * mat_B[186][0] +
                mat_A[6][0] * mat_B[194][0] +
                mat_A[6][1] * mat_B[202][0] +
                mat_A[6][2] * mat_B[210][0] +
                mat_A[6][3] * mat_B[218][0] +
                mat_A[7][0] * mat_B[226][0] +
                mat_A[7][1] * mat_B[234][0] +
                mat_A[7][2] * mat_B[242][0] +
                mat_A[7][3] * mat_B[250][0];
    mat_C[2][1] <=
                mat_A[0][0] * mat_B[2][1] +
                mat_A[0][1] * mat_B[10][1] +
                mat_A[0][2] * mat_B[18][1] +
                mat_A[0][3] * mat_B[26][1] +
                mat_A[1][0] * mat_B[34][1] +
                mat_A[1][1] * mat_B[42][1] +
                mat_A[1][2] * mat_B[50][1] +
                mat_A[1][3] * mat_B[58][1] +
                mat_A[2][0] * mat_B[66][1] +
                mat_A[2][1] * mat_B[74][1] +
                mat_A[2][2] * mat_B[82][1] +
                mat_A[2][3] * mat_B[90][1] +
                mat_A[3][0] * mat_B[98][1] +
                mat_A[3][1] * mat_B[106][1] +
                mat_A[3][2] * mat_B[114][1] +
                mat_A[3][3] * mat_B[122][1] +
                mat_A[4][0] * mat_B[130][1] +
                mat_A[4][1] * mat_B[138][1] +
                mat_A[4][2] * mat_B[146][1] +
                mat_A[4][3] * mat_B[154][1] +
                mat_A[5][0] * mat_B[162][1] +
                mat_A[5][1] * mat_B[170][1] +
                mat_A[5][2] * mat_B[178][1] +
                mat_A[5][3] * mat_B[186][1] +
                mat_A[6][0] * mat_B[194][1] +
                mat_A[6][1] * mat_B[202][1] +
                mat_A[6][2] * mat_B[210][1] +
                mat_A[6][3] * mat_B[218][1] +
                mat_A[7][0] * mat_B[226][1] +
                mat_A[7][1] * mat_B[234][1] +
                mat_A[7][2] * mat_B[242][1] +
                mat_A[7][3] * mat_B[250][1];
    mat_C[2][2] <=
                mat_A[0][0] * mat_B[2][2] +
                mat_A[0][1] * mat_B[10][2] +
                mat_A[0][2] * mat_B[18][2] +
                mat_A[0][3] * mat_B[26][2] +
                mat_A[1][0] * mat_B[34][2] +
                mat_A[1][1] * mat_B[42][2] +
                mat_A[1][2] * mat_B[50][2] +
                mat_A[1][3] * mat_B[58][2] +
                mat_A[2][0] * mat_B[66][2] +
                mat_A[2][1] * mat_B[74][2] +
                mat_A[2][2] * mat_B[82][2] +
                mat_A[2][3] * mat_B[90][2] +
                mat_A[3][0] * mat_B[98][2] +
                mat_A[3][1] * mat_B[106][2] +
                mat_A[3][2] * mat_B[114][2] +
                mat_A[3][3] * mat_B[122][2] +
                mat_A[4][0] * mat_B[130][2] +
                mat_A[4][1] * mat_B[138][2] +
                mat_A[4][2] * mat_B[146][2] +
                mat_A[4][3] * mat_B[154][2] +
                mat_A[5][0] * mat_B[162][2] +
                mat_A[5][1] * mat_B[170][2] +
                mat_A[5][2] * mat_B[178][2] +
                mat_A[5][3] * mat_B[186][2] +
                mat_A[6][0] * mat_B[194][2] +
                mat_A[6][1] * mat_B[202][2] +
                mat_A[6][2] * mat_B[210][2] +
                mat_A[6][3] * mat_B[218][2] +
                mat_A[7][0] * mat_B[226][2] +
                mat_A[7][1] * mat_B[234][2] +
                mat_A[7][2] * mat_B[242][2] +
                mat_A[7][3] * mat_B[250][2];
    mat_C[2][3] <=
                mat_A[0][0] * mat_B[2][3] +
                mat_A[0][1] * mat_B[10][3] +
                mat_A[0][2] * mat_B[18][3] +
                mat_A[0][3] * mat_B[26][3] +
                mat_A[1][0] * mat_B[34][3] +
                mat_A[1][1] * mat_B[42][3] +
                mat_A[1][2] * mat_B[50][3] +
                mat_A[1][3] * mat_B[58][3] +
                mat_A[2][0] * mat_B[66][3] +
                mat_A[2][1] * mat_B[74][3] +
                mat_A[2][2] * mat_B[82][3] +
                mat_A[2][3] * mat_B[90][3] +
                mat_A[3][0] * mat_B[98][3] +
                mat_A[3][1] * mat_B[106][3] +
                mat_A[3][2] * mat_B[114][3] +
                mat_A[3][3] * mat_B[122][3] +
                mat_A[4][0] * mat_B[130][3] +
                mat_A[4][1] * mat_B[138][3] +
                mat_A[4][2] * mat_B[146][3] +
                mat_A[4][3] * mat_B[154][3] +
                mat_A[5][0] * mat_B[162][3] +
                mat_A[5][1] * mat_B[170][3] +
                mat_A[5][2] * mat_B[178][3] +
                mat_A[5][3] * mat_B[186][3] +
                mat_A[6][0] * mat_B[194][3] +
                mat_A[6][1] * mat_B[202][3] +
                mat_A[6][2] * mat_B[210][3] +
                mat_A[6][3] * mat_B[218][3] +
                mat_A[7][0] * mat_B[226][3] +
                mat_A[7][1] * mat_B[234][3] +
                mat_A[7][2] * mat_B[242][3] +
                mat_A[7][3] * mat_B[250][3];
    mat_C[3][0] <=
                mat_A[0][0] * mat_B[3][0] +
                mat_A[0][1] * mat_B[11][0] +
                mat_A[0][2] * mat_B[19][0] +
                mat_A[0][3] * mat_B[27][0] +
                mat_A[1][0] * mat_B[35][0] +
                mat_A[1][1] * mat_B[43][0] +
                mat_A[1][2] * mat_B[51][0] +
                mat_A[1][3] * mat_B[59][0] +
                mat_A[2][0] * mat_B[67][0] +
                mat_A[2][1] * mat_B[75][0] +
                mat_A[2][2] * mat_B[83][0] +
                mat_A[2][3] * mat_B[91][0] +
                mat_A[3][0] * mat_B[99][0] +
                mat_A[3][1] * mat_B[107][0] +
                mat_A[3][2] * mat_B[115][0] +
                mat_A[3][3] * mat_B[123][0] +
                mat_A[4][0] * mat_B[131][0] +
                mat_A[4][1] * mat_B[139][0] +
                mat_A[4][2] * mat_B[147][0] +
                mat_A[4][3] * mat_B[155][0] +
                mat_A[5][0] * mat_B[163][0] +
                mat_A[5][1] * mat_B[171][0] +
                mat_A[5][2] * mat_B[179][0] +
                mat_A[5][3] * mat_B[187][0] +
                mat_A[6][0] * mat_B[195][0] +
                mat_A[6][1] * mat_B[203][0] +
                mat_A[6][2] * mat_B[211][0] +
                mat_A[6][3] * mat_B[219][0] +
                mat_A[7][0] * mat_B[227][0] +
                mat_A[7][1] * mat_B[235][0] +
                mat_A[7][2] * mat_B[243][0] +
                mat_A[7][3] * mat_B[251][0];
    mat_C[3][1] <=
                mat_A[0][0] * mat_B[3][1] +
                mat_A[0][1] * mat_B[11][1] +
                mat_A[0][2] * mat_B[19][1] +
                mat_A[0][3] * mat_B[27][1] +
                mat_A[1][0] * mat_B[35][1] +
                mat_A[1][1] * mat_B[43][1] +
                mat_A[1][2] * mat_B[51][1] +
                mat_A[1][3] * mat_B[59][1] +
                mat_A[2][0] * mat_B[67][1] +
                mat_A[2][1] * mat_B[75][1] +
                mat_A[2][2] * mat_B[83][1] +
                mat_A[2][3] * mat_B[91][1] +
                mat_A[3][0] * mat_B[99][1] +
                mat_A[3][1] * mat_B[107][1] +
                mat_A[3][2] * mat_B[115][1] +
                mat_A[3][3] * mat_B[123][1] +
                mat_A[4][0] * mat_B[131][1] +
                mat_A[4][1] * mat_B[139][1] +
                mat_A[4][2] * mat_B[147][1] +
                mat_A[4][3] * mat_B[155][1] +
                mat_A[5][0] * mat_B[163][1] +
                mat_A[5][1] * mat_B[171][1] +
                mat_A[5][2] * mat_B[179][1] +
                mat_A[5][3] * mat_B[187][1] +
                mat_A[6][0] * mat_B[195][1] +
                mat_A[6][1] * mat_B[203][1] +
                mat_A[6][2] * mat_B[211][1] +
                mat_A[6][3] * mat_B[219][1] +
                mat_A[7][0] * mat_B[227][1] +
                mat_A[7][1] * mat_B[235][1] +
                mat_A[7][2] * mat_B[243][1] +
                mat_A[7][3] * mat_B[251][1];
    mat_C[3][2] <=
                mat_A[0][0] * mat_B[3][2] +
                mat_A[0][1] * mat_B[11][2] +
                mat_A[0][2] * mat_B[19][2] +
                mat_A[0][3] * mat_B[27][2] +
                mat_A[1][0] * mat_B[35][2] +
                mat_A[1][1] * mat_B[43][2] +
                mat_A[1][2] * mat_B[51][2] +
                mat_A[1][3] * mat_B[59][2] +
                mat_A[2][0] * mat_B[67][2] +
                mat_A[2][1] * mat_B[75][2] +
                mat_A[2][2] * mat_B[83][2] +
                mat_A[2][3] * mat_B[91][2] +
                mat_A[3][0] * mat_B[99][2] +
                mat_A[3][1] * mat_B[107][2] +
                mat_A[3][2] * mat_B[115][2] +
                mat_A[3][3] * mat_B[123][2] +
                mat_A[4][0] * mat_B[131][2] +
                mat_A[4][1] * mat_B[139][2] +
                mat_A[4][2] * mat_B[147][2] +
                mat_A[4][3] * mat_B[155][2] +
                mat_A[5][0] * mat_B[163][2] +
                mat_A[5][1] * mat_B[171][2] +
                mat_A[5][2] * mat_B[179][2] +
                mat_A[5][3] * mat_B[187][2] +
                mat_A[6][0] * mat_B[195][2] +
                mat_A[6][1] * mat_B[203][2] +
                mat_A[6][2] * mat_B[211][2] +
                mat_A[6][3] * mat_B[219][2] +
                mat_A[7][0] * mat_B[227][2] +
                mat_A[7][1] * mat_B[235][2] +
                mat_A[7][2] * mat_B[243][2] +
                mat_A[7][3] * mat_B[251][2];
    mat_C[3][3] <=
                mat_A[0][0] * mat_B[3][3] +
                mat_A[0][1] * mat_B[11][3] +
                mat_A[0][2] * mat_B[19][3] +
                mat_A[0][3] * mat_B[27][3] +
                mat_A[1][0] * mat_B[35][3] +
                mat_A[1][1] * mat_B[43][3] +
                mat_A[1][2] * mat_B[51][3] +
                mat_A[1][3] * mat_B[59][3] +
                mat_A[2][0] * mat_B[67][3] +
                mat_A[2][1] * mat_B[75][3] +
                mat_A[2][2] * mat_B[83][3] +
                mat_A[2][3] * mat_B[91][3] +
                mat_A[3][0] * mat_B[99][3] +
                mat_A[3][1] * mat_B[107][3] +
                mat_A[3][2] * mat_B[115][3] +
                mat_A[3][3] * mat_B[123][3] +
                mat_A[4][0] * mat_B[131][3] +
                mat_A[4][1] * mat_B[139][3] +
                mat_A[4][2] * mat_B[147][3] +
                mat_A[4][3] * mat_B[155][3] +
                mat_A[5][0] * mat_B[163][3] +
                mat_A[5][1] * mat_B[171][3] +
                mat_A[5][2] * mat_B[179][3] +
                mat_A[5][3] * mat_B[187][3] +
                mat_A[6][0] * mat_B[195][3] +
                mat_A[6][1] * mat_B[203][3] +
                mat_A[6][2] * mat_B[211][3] +
                mat_A[6][3] * mat_B[219][3] +
                mat_A[7][0] * mat_B[227][3] +
                mat_A[7][1] * mat_B[235][3] +
                mat_A[7][2] * mat_B[243][3] +
                mat_A[7][3] * mat_B[251][3];
    mat_C[4][0] <=
                mat_A[0][0] * mat_B[4][0] +
                mat_A[0][1] * mat_B[12][0] +
                mat_A[0][2] * mat_B[20][0] +
                mat_A[0][3] * mat_B[28][0] +
                mat_A[1][0] * mat_B[36][0] +
                mat_A[1][1] * mat_B[44][0] +
                mat_A[1][2] * mat_B[52][0] +
                mat_A[1][3] * mat_B[60][0] +
                mat_A[2][0] * mat_B[68][0] +
                mat_A[2][1] * mat_B[76][0] +
                mat_A[2][2] * mat_B[84][0] +
                mat_A[2][3] * mat_B[92][0] +
                mat_A[3][0] * mat_B[100][0] +
                mat_A[3][1] * mat_B[108][0] +
                mat_A[3][2] * mat_B[116][0] +
                mat_A[3][3] * mat_B[124][0] +
                mat_A[4][0] * mat_B[132][0] +
                mat_A[4][1] * mat_B[140][0] +
                mat_A[4][2] * mat_B[148][0] +
                mat_A[4][3] * mat_B[156][0] +
                mat_A[5][0] * mat_B[164][0] +
                mat_A[5][1] * mat_B[172][0] +
                mat_A[5][2] * mat_B[180][0] +
                mat_A[5][3] * mat_B[188][0] +
                mat_A[6][0] * mat_B[196][0] +
                mat_A[6][1] * mat_B[204][0] +
                mat_A[6][2] * mat_B[212][0] +
                mat_A[6][3] * mat_B[220][0] +
                mat_A[7][0] * mat_B[228][0] +
                mat_A[7][1] * mat_B[236][0] +
                mat_A[7][2] * mat_B[244][0] +
                mat_A[7][3] * mat_B[252][0];
    mat_C[4][1] <=
                mat_A[0][0] * mat_B[4][1] +
                mat_A[0][1] * mat_B[12][1] +
                mat_A[0][2] * mat_B[20][1] +
                mat_A[0][3] * mat_B[28][1] +
                mat_A[1][0] * mat_B[36][1] +
                mat_A[1][1] * mat_B[44][1] +
                mat_A[1][2] * mat_B[52][1] +
                mat_A[1][3] * mat_B[60][1] +
                mat_A[2][0] * mat_B[68][1] +
                mat_A[2][1] * mat_B[76][1] +
                mat_A[2][2] * mat_B[84][1] +
                mat_A[2][3] * mat_B[92][1] +
                mat_A[3][0] * mat_B[100][1] +
                mat_A[3][1] * mat_B[108][1] +
                mat_A[3][2] * mat_B[116][1] +
                mat_A[3][3] * mat_B[124][1] +
                mat_A[4][0] * mat_B[132][1] +
                mat_A[4][1] * mat_B[140][1] +
                mat_A[4][2] * mat_B[148][1] +
                mat_A[4][3] * mat_B[156][1] +
                mat_A[5][0] * mat_B[164][1] +
                mat_A[5][1] * mat_B[172][1] +
                mat_A[5][2] * mat_B[180][1] +
                mat_A[5][3] * mat_B[188][1] +
                mat_A[6][0] * mat_B[196][1] +
                mat_A[6][1] * mat_B[204][1] +
                mat_A[6][2] * mat_B[212][1] +
                mat_A[6][3] * mat_B[220][1] +
                mat_A[7][0] * mat_B[228][1] +
                mat_A[7][1] * mat_B[236][1] +
                mat_A[7][2] * mat_B[244][1] +
                mat_A[7][3] * mat_B[252][1];
    mat_C[4][2] <=
                mat_A[0][0] * mat_B[4][2] +
                mat_A[0][1] * mat_B[12][2] +
                mat_A[0][2] * mat_B[20][2] +
                mat_A[0][3] * mat_B[28][2] +
                mat_A[1][0] * mat_B[36][2] +
                mat_A[1][1] * mat_B[44][2] +
                mat_A[1][2] * mat_B[52][2] +
                mat_A[1][3] * mat_B[60][2] +
                mat_A[2][0] * mat_B[68][2] +
                mat_A[2][1] * mat_B[76][2] +
                mat_A[2][2] * mat_B[84][2] +
                mat_A[2][3] * mat_B[92][2] +
                mat_A[3][0] * mat_B[100][2] +
                mat_A[3][1] * mat_B[108][2] +
                mat_A[3][2] * mat_B[116][2] +
                mat_A[3][3] * mat_B[124][2] +
                mat_A[4][0] * mat_B[132][2] +
                mat_A[4][1] * mat_B[140][2] +
                mat_A[4][2] * mat_B[148][2] +
                mat_A[4][3] * mat_B[156][2] +
                mat_A[5][0] * mat_B[164][2] +
                mat_A[5][1] * mat_B[172][2] +
                mat_A[5][2] * mat_B[180][2] +
                mat_A[5][3] * mat_B[188][2] +
                mat_A[6][0] * mat_B[196][2] +
                mat_A[6][1] * mat_B[204][2] +
                mat_A[6][2] * mat_B[212][2] +
                mat_A[6][3] * mat_B[220][2] +
                mat_A[7][0] * mat_B[228][2] +
                mat_A[7][1] * mat_B[236][2] +
                mat_A[7][2] * mat_B[244][2] +
                mat_A[7][3] * mat_B[252][2];
    mat_C[4][3] <=
                mat_A[0][0] * mat_B[4][3] +
                mat_A[0][1] * mat_B[12][3] +
                mat_A[0][2] * mat_B[20][3] +
                mat_A[0][3] * mat_B[28][3] +
                mat_A[1][0] * mat_B[36][3] +
                mat_A[1][1] * mat_B[44][3] +
                mat_A[1][2] * mat_B[52][3] +
                mat_A[1][3] * mat_B[60][3] +
                mat_A[2][0] * mat_B[68][3] +
                mat_A[2][1] * mat_B[76][3] +
                mat_A[2][2] * mat_B[84][3] +
                mat_A[2][3] * mat_B[92][3] +
                mat_A[3][0] * mat_B[100][3] +
                mat_A[3][1] * mat_B[108][3] +
                mat_A[3][2] * mat_B[116][3] +
                mat_A[3][3] * mat_B[124][3] +
                mat_A[4][0] * mat_B[132][3] +
                mat_A[4][1] * mat_B[140][3] +
                mat_A[4][2] * mat_B[148][3] +
                mat_A[4][3] * mat_B[156][3] +
                mat_A[5][0] * mat_B[164][3] +
                mat_A[5][1] * mat_B[172][3] +
                mat_A[5][2] * mat_B[180][3] +
                mat_A[5][3] * mat_B[188][3] +
                mat_A[6][0] * mat_B[196][3] +
                mat_A[6][1] * mat_B[204][3] +
                mat_A[6][2] * mat_B[212][3] +
                mat_A[6][3] * mat_B[220][3] +
                mat_A[7][0] * mat_B[228][3] +
                mat_A[7][1] * mat_B[236][3] +
                mat_A[7][2] * mat_B[244][3] +
                mat_A[7][3] * mat_B[252][3];
    mat_C[5][0] <=
                mat_A[0][0] * mat_B[5][0] +
                mat_A[0][1] * mat_B[13][0] +
                mat_A[0][2] * mat_B[21][0] +
                mat_A[0][3] * mat_B[29][0] +
                mat_A[1][0] * mat_B[37][0] +
                mat_A[1][1] * mat_B[45][0] +
                mat_A[1][2] * mat_B[53][0] +
                mat_A[1][3] * mat_B[61][0] +
                mat_A[2][0] * mat_B[69][0] +
                mat_A[2][1] * mat_B[77][0] +
                mat_A[2][2] * mat_B[85][0] +
                mat_A[2][3] * mat_B[93][0] +
                mat_A[3][0] * mat_B[101][0] +
                mat_A[3][1] * mat_B[109][0] +
                mat_A[3][2] * mat_B[117][0] +
                mat_A[3][3] * mat_B[125][0] +
                mat_A[4][0] * mat_B[133][0] +
                mat_A[4][1] * mat_B[141][0] +
                mat_A[4][2] * mat_B[149][0] +
                mat_A[4][3] * mat_B[157][0] +
                mat_A[5][0] * mat_B[165][0] +
                mat_A[5][1] * mat_B[173][0] +
                mat_A[5][2] * mat_B[181][0] +
                mat_A[5][3] * mat_B[189][0] +
                mat_A[6][0] * mat_B[197][0] +
                mat_A[6][1] * mat_B[205][0] +
                mat_A[6][2] * mat_B[213][0] +
                mat_A[6][3] * mat_B[221][0] +
                mat_A[7][0] * mat_B[229][0] +
                mat_A[7][1] * mat_B[237][0] +
                mat_A[7][2] * mat_B[245][0] +
                mat_A[7][3] * mat_B[253][0];
    mat_C[5][1] <=
                mat_A[0][0] * mat_B[5][1] +
                mat_A[0][1] * mat_B[13][1] +
                mat_A[0][2] * mat_B[21][1] +
                mat_A[0][3] * mat_B[29][1] +
                mat_A[1][0] * mat_B[37][1] +
                mat_A[1][1] * mat_B[45][1] +
                mat_A[1][2] * mat_B[53][1] +
                mat_A[1][3] * mat_B[61][1] +
                mat_A[2][0] * mat_B[69][1] +
                mat_A[2][1] * mat_B[77][1] +
                mat_A[2][2] * mat_B[85][1] +
                mat_A[2][3] * mat_B[93][1] +
                mat_A[3][0] * mat_B[101][1] +
                mat_A[3][1] * mat_B[109][1] +
                mat_A[3][2] * mat_B[117][1] +
                mat_A[3][3] * mat_B[125][1] +
                mat_A[4][0] * mat_B[133][1] +
                mat_A[4][1] * mat_B[141][1] +
                mat_A[4][2] * mat_B[149][1] +
                mat_A[4][3] * mat_B[157][1] +
                mat_A[5][0] * mat_B[165][1] +
                mat_A[5][1] * mat_B[173][1] +
                mat_A[5][2] * mat_B[181][1] +
                mat_A[5][3] * mat_B[189][1] +
                mat_A[6][0] * mat_B[197][1] +
                mat_A[6][1] * mat_B[205][1] +
                mat_A[6][2] * mat_B[213][1] +
                mat_A[6][3] * mat_B[221][1] +
                mat_A[7][0] * mat_B[229][1] +
                mat_A[7][1] * mat_B[237][1] +
                mat_A[7][2] * mat_B[245][1] +
                mat_A[7][3] * mat_B[253][1];
    mat_C[5][2] <=
                mat_A[0][0] * mat_B[5][2] +
                mat_A[0][1] * mat_B[13][2] +
                mat_A[0][2] * mat_B[21][2] +
                mat_A[0][3] * mat_B[29][2] +
                mat_A[1][0] * mat_B[37][2] +
                mat_A[1][1] * mat_B[45][2] +
                mat_A[1][2] * mat_B[53][2] +
                mat_A[1][3] * mat_B[61][2] +
                mat_A[2][0] * mat_B[69][2] +
                mat_A[2][1] * mat_B[77][2] +
                mat_A[2][2] * mat_B[85][2] +
                mat_A[2][3] * mat_B[93][2] +
                mat_A[3][0] * mat_B[101][2] +
                mat_A[3][1] * mat_B[109][2] +
                mat_A[3][2] * mat_B[117][2] +
                mat_A[3][3] * mat_B[125][2] +
                mat_A[4][0] * mat_B[133][2] +
                mat_A[4][1] * mat_B[141][2] +
                mat_A[4][2] * mat_B[149][2] +
                mat_A[4][3] * mat_B[157][2] +
                mat_A[5][0] * mat_B[165][2] +
                mat_A[5][1] * mat_B[173][2] +
                mat_A[5][2] * mat_B[181][2] +
                mat_A[5][3] * mat_B[189][2] +
                mat_A[6][0] * mat_B[197][2] +
                mat_A[6][1] * mat_B[205][2] +
                mat_A[6][2] * mat_B[213][2] +
                mat_A[6][3] * mat_B[221][2] +
                mat_A[7][0] * mat_B[229][2] +
                mat_A[7][1] * mat_B[237][2] +
                mat_A[7][2] * mat_B[245][2] +
                mat_A[7][3] * mat_B[253][2];
    mat_C[5][3] <=
                mat_A[0][0] * mat_B[5][3] +
                mat_A[0][1] * mat_B[13][3] +
                mat_A[0][2] * mat_B[21][3] +
                mat_A[0][3] * mat_B[29][3] +
                mat_A[1][0] * mat_B[37][3] +
                mat_A[1][1] * mat_B[45][3] +
                mat_A[1][2] * mat_B[53][3] +
                mat_A[1][3] * mat_B[61][3] +
                mat_A[2][0] * mat_B[69][3] +
                mat_A[2][1] * mat_B[77][3] +
                mat_A[2][2] * mat_B[85][3] +
                mat_A[2][3] * mat_B[93][3] +
                mat_A[3][0] * mat_B[101][3] +
                mat_A[3][1] * mat_B[109][3] +
                mat_A[3][2] * mat_B[117][3] +
                mat_A[3][3] * mat_B[125][3] +
                mat_A[4][0] * mat_B[133][3] +
                mat_A[4][1] * mat_B[141][3] +
                mat_A[4][2] * mat_B[149][3] +
                mat_A[4][3] * mat_B[157][3] +
                mat_A[5][0] * mat_B[165][3] +
                mat_A[5][1] * mat_B[173][3] +
                mat_A[5][2] * mat_B[181][3] +
                mat_A[5][3] * mat_B[189][3] +
                mat_A[6][0] * mat_B[197][3] +
                mat_A[6][1] * mat_B[205][3] +
                mat_A[6][2] * mat_B[213][3] +
                mat_A[6][3] * mat_B[221][3] +
                mat_A[7][0] * mat_B[229][3] +
                mat_A[7][1] * mat_B[237][3] +
                mat_A[7][2] * mat_B[245][3] +
                mat_A[7][3] * mat_B[253][3];
    mat_C[6][0] <=
                mat_A[0][0] * mat_B[6][0] +
                mat_A[0][1] * mat_B[14][0] +
                mat_A[0][2] * mat_B[22][0] +
                mat_A[0][3] * mat_B[30][0] +
                mat_A[1][0] * mat_B[38][0] +
                mat_A[1][1] * mat_B[46][0] +
                mat_A[1][2] * mat_B[54][0] +
                mat_A[1][3] * mat_B[62][0] +
                mat_A[2][0] * mat_B[70][0] +
                mat_A[2][1] * mat_B[78][0] +
                mat_A[2][2] * mat_B[86][0] +
                mat_A[2][3] * mat_B[94][0] +
                mat_A[3][0] * mat_B[102][0] +
                mat_A[3][1] * mat_B[110][0] +
                mat_A[3][2] * mat_B[118][0] +
                mat_A[3][3] * mat_B[126][0] +
                mat_A[4][0] * mat_B[134][0] +
                mat_A[4][1] * mat_B[142][0] +
                mat_A[4][2] * mat_B[150][0] +
                mat_A[4][3] * mat_B[158][0] +
                mat_A[5][0] * mat_B[166][0] +
                mat_A[5][1] * mat_B[174][0] +
                mat_A[5][2] * mat_B[182][0] +
                mat_A[5][3] * mat_B[190][0] +
                mat_A[6][0] * mat_B[198][0] +
                mat_A[6][1] * mat_B[206][0] +
                mat_A[6][2] * mat_B[214][0] +
                mat_A[6][3] * mat_B[222][0] +
                mat_A[7][0] * mat_B[230][0] +
                mat_A[7][1] * mat_B[238][0] +
                mat_A[7][2] * mat_B[246][0] +
                mat_A[7][3] * mat_B[254][0];
    mat_C[6][1] <=
                mat_A[0][0] * mat_B[6][1] +
                mat_A[0][1] * mat_B[14][1] +
                mat_A[0][2] * mat_B[22][1] +
                mat_A[0][3] * mat_B[30][1] +
                mat_A[1][0] * mat_B[38][1] +
                mat_A[1][1] * mat_B[46][1] +
                mat_A[1][2] * mat_B[54][1] +
                mat_A[1][3] * mat_B[62][1] +
                mat_A[2][0] * mat_B[70][1] +
                mat_A[2][1] * mat_B[78][1] +
                mat_A[2][2] * mat_B[86][1] +
                mat_A[2][3] * mat_B[94][1] +
                mat_A[3][0] * mat_B[102][1] +
                mat_A[3][1] * mat_B[110][1] +
                mat_A[3][2] * mat_B[118][1] +
                mat_A[3][3] * mat_B[126][1] +
                mat_A[4][0] * mat_B[134][1] +
                mat_A[4][1] * mat_B[142][1] +
                mat_A[4][2] * mat_B[150][1] +
                mat_A[4][3] * mat_B[158][1] +
                mat_A[5][0] * mat_B[166][1] +
                mat_A[5][1] * mat_B[174][1] +
                mat_A[5][2] * mat_B[182][1] +
                mat_A[5][3] * mat_B[190][1] +
                mat_A[6][0] * mat_B[198][1] +
                mat_A[6][1] * mat_B[206][1] +
                mat_A[6][2] * mat_B[214][1] +
                mat_A[6][3] * mat_B[222][1] +
                mat_A[7][0] * mat_B[230][1] +
                mat_A[7][1] * mat_B[238][1] +
                mat_A[7][2] * mat_B[246][1] +
                mat_A[7][3] * mat_B[254][1];
    mat_C[6][2] <=
                mat_A[0][0] * mat_B[6][2] +
                mat_A[0][1] * mat_B[14][2] +
                mat_A[0][2] * mat_B[22][2] +
                mat_A[0][3] * mat_B[30][2] +
                mat_A[1][0] * mat_B[38][2] +
                mat_A[1][1] * mat_B[46][2] +
                mat_A[1][2] * mat_B[54][2] +
                mat_A[1][3] * mat_B[62][2] +
                mat_A[2][0] * mat_B[70][2] +
                mat_A[2][1] * mat_B[78][2] +
                mat_A[2][2] * mat_B[86][2] +
                mat_A[2][3] * mat_B[94][2] +
                mat_A[3][0] * mat_B[102][2] +
                mat_A[3][1] * mat_B[110][2] +
                mat_A[3][2] * mat_B[118][2] +
                mat_A[3][3] * mat_B[126][2] +
                mat_A[4][0] * mat_B[134][2] +
                mat_A[4][1] * mat_B[142][2] +
                mat_A[4][2] * mat_B[150][2] +
                mat_A[4][3] * mat_B[158][2] +
                mat_A[5][0] * mat_B[166][2] +
                mat_A[5][1] * mat_B[174][2] +
                mat_A[5][2] * mat_B[182][2] +
                mat_A[5][3] * mat_B[190][2] +
                mat_A[6][0] * mat_B[198][2] +
                mat_A[6][1] * mat_B[206][2] +
                mat_A[6][2] * mat_B[214][2] +
                mat_A[6][3] * mat_B[222][2] +
                mat_A[7][0] * mat_B[230][2] +
                mat_A[7][1] * mat_B[238][2] +
                mat_A[7][2] * mat_B[246][2] +
                mat_A[7][3] * mat_B[254][2];
    mat_C[6][3] <=
                mat_A[0][0] * mat_B[6][3] +
                mat_A[0][1] * mat_B[14][3] +
                mat_A[0][2] * mat_B[22][3] +
                mat_A[0][3] * mat_B[30][3] +
                mat_A[1][0] * mat_B[38][3] +
                mat_A[1][1] * mat_B[46][3] +
                mat_A[1][2] * mat_B[54][3] +
                mat_A[1][3] * mat_B[62][3] +
                mat_A[2][0] * mat_B[70][3] +
                mat_A[2][1] * mat_B[78][3] +
                mat_A[2][2] * mat_B[86][3] +
                mat_A[2][3] * mat_B[94][3] +
                mat_A[3][0] * mat_B[102][3] +
                mat_A[3][1] * mat_B[110][3] +
                mat_A[3][2] * mat_B[118][3] +
                mat_A[3][3] * mat_B[126][3] +
                mat_A[4][0] * mat_B[134][3] +
                mat_A[4][1] * mat_B[142][3] +
                mat_A[4][2] * mat_B[150][3] +
                mat_A[4][3] * mat_B[158][3] +
                mat_A[5][0] * mat_B[166][3] +
                mat_A[5][1] * mat_B[174][3] +
                mat_A[5][2] * mat_B[182][3] +
                mat_A[5][3] * mat_B[190][3] +
                mat_A[6][0] * mat_B[198][3] +
                mat_A[6][1] * mat_B[206][3] +
                mat_A[6][2] * mat_B[214][3] +
                mat_A[6][3] * mat_B[222][3] +
                mat_A[7][0] * mat_B[230][3] +
                mat_A[7][1] * mat_B[238][3] +
                mat_A[7][2] * mat_B[246][3] +
                mat_A[7][3] * mat_B[254][3];
    mat_C[7][0] <=
                mat_A[0][0] * mat_B[7][0] +
                mat_A[0][1] * mat_B[15][0] +
                mat_A[0][2] * mat_B[23][0] +
                mat_A[0][3] * mat_B[31][0] +
                mat_A[1][0] * mat_B[39][0] +
                mat_A[1][1] * mat_B[47][0] +
                mat_A[1][2] * mat_B[55][0] +
                mat_A[1][3] * mat_B[63][0] +
                mat_A[2][0] * mat_B[71][0] +
                mat_A[2][1] * mat_B[79][0] +
                mat_A[2][2] * mat_B[87][0] +
                mat_A[2][3] * mat_B[95][0] +
                mat_A[3][0] * mat_B[103][0] +
                mat_A[3][1] * mat_B[111][0] +
                mat_A[3][2] * mat_B[119][0] +
                mat_A[3][3] * mat_B[127][0] +
                mat_A[4][0] * mat_B[135][0] +
                mat_A[4][1] * mat_B[143][0] +
                mat_A[4][2] * mat_B[151][0] +
                mat_A[4][3] * mat_B[159][0] +
                mat_A[5][0] * mat_B[167][0] +
                mat_A[5][1] * mat_B[175][0] +
                mat_A[5][2] * mat_B[183][0] +
                mat_A[5][3] * mat_B[191][0] +
                mat_A[6][0] * mat_B[199][0] +
                mat_A[6][1] * mat_B[207][0] +
                mat_A[6][2] * mat_B[215][0] +
                mat_A[6][3] * mat_B[223][0] +
                mat_A[7][0] * mat_B[231][0] +
                mat_A[7][1] * mat_B[239][0] +
                mat_A[7][2] * mat_B[247][0] +
                mat_A[7][3] * mat_B[255][0];
    mat_C[7][1] <=
                mat_A[0][0] * mat_B[7][1] +
                mat_A[0][1] * mat_B[15][1] +
                mat_A[0][2] * mat_B[23][1] +
                mat_A[0][3] * mat_B[31][1] +
                mat_A[1][0] * mat_B[39][1] +
                mat_A[1][1] * mat_B[47][1] +
                mat_A[1][2] * mat_B[55][1] +
                mat_A[1][3] * mat_B[63][1] +
                mat_A[2][0] * mat_B[71][1] +
                mat_A[2][1] * mat_B[79][1] +
                mat_A[2][2] * mat_B[87][1] +
                mat_A[2][3] * mat_B[95][1] +
                mat_A[3][0] * mat_B[103][1] +
                mat_A[3][1] * mat_B[111][1] +
                mat_A[3][2] * mat_B[119][1] +
                mat_A[3][3] * mat_B[127][1] +
                mat_A[4][0] * mat_B[135][1] +
                mat_A[4][1] * mat_B[143][1] +
                mat_A[4][2] * mat_B[151][1] +
                mat_A[4][3] * mat_B[159][1] +
                mat_A[5][0] * mat_B[167][1] +
                mat_A[5][1] * mat_B[175][1] +
                mat_A[5][2] * mat_B[183][1] +
                mat_A[5][3] * mat_B[191][1] +
                mat_A[6][0] * mat_B[199][1] +
                mat_A[6][1] * mat_B[207][1] +
                mat_A[6][2] * mat_B[215][1] +
                mat_A[6][3] * mat_B[223][1] +
                mat_A[7][0] * mat_B[231][1] +
                mat_A[7][1] * mat_B[239][1] +
                mat_A[7][2] * mat_B[247][1] +
                mat_A[7][3] * mat_B[255][1];
    mat_C[7][2] <=
                mat_A[0][0] * mat_B[7][2] +
                mat_A[0][1] * mat_B[15][2] +
                mat_A[0][2] * mat_B[23][2] +
                mat_A[0][3] * mat_B[31][2] +
                mat_A[1][0] * mat_B[39][2] +
                mat_A[1][1] * mat_B[47][2] +
                mat_A[1][2] * mat_B[55][2] +
                mat_A[1][3] * mat_B[63][2] +
                mat_A[2][0] * mat_B[71][2] +
                mat_A[2][1] * mat_B[79][2] +
                mat_A[2][2] * mat_B[87][2] +
                mat_A[2][3] * mat_B[95][2] +
                mat_A[3][0] * mat_B[103][2] +
                mat_A[3][1] * mat_B[111][2] +
                mat_A[3][2] * mat_B[119][2] +
                mat_A[3][3] * mat_B[127][2] +
                mat_A[4][0] * mat_B[135][2] +
                mat_A[4][1] * mat_B[143][2] +
                mat_A[4][2] * mat_B[151][2] +
                mat_A[4][3] * mat_B[159][2] +
                mat_A[5][0] * mat_B[167][2] +
                mat_A[5][1] * mat_B[175][2] +
                mat_A[5][2] * mat_B[183][2] +
                mat_A[5][3] * mat_B[191][2] +
                mat_A[6][0] * mat_B[199][2] +
                mat_A[6][1] * mat_B[207][2] +
                mat_A[6][2] * mat_B[215][2] +
                mat_A[6][3] * mat_B[223][2] +
                mat_A[7][0] * mat_B[231][2] +
                mat_A[7][1] * mat_B[239][2] +
                mat_A[7][2] * mat_B[247][2] +
                mat_A[7][3] * mat_B[255][2];
    mat_C[7][3] <=
                mat_A[0][0] * mat_B[7][3] +
                mat_A[0][1] * mat_B[15][3] +
                mat_A[0][2] * mat_B[23][3] +
                mat_A[0][3] * mat_B[31][3] +
                mat_A[1][0] * mat_B[39][3] +
                mat_A[1][1] * mat_B[47][3] +
                mat_A[1][2] * mat_B[55][3] +
                mat_A[1][3] * mat_B[63][3] +
                mat_A[2][0] * mat_B[71][3] +
                mat_A[2][1] * mat_B[79][3] +
                mat_A[2][2] * mat_B[87][3] +
                mat_A[2][3] * mat_B[95][3] +
                mat_A[3][0] * mat_B[103][3] +
                mat_A[3][1] * mat_B[111][3] +
                mat_A[3][2] * mat_B[119][3] +
                mat_A[3][3] * mat_B[127][3] +
                mat_A[4][0] * mat_B[135][3] +
                mat_A[4][1] * mat_B[143][3] +
                mat_A[4][2] * mat_B[151][3] +
                mat_A[4][3] * mat_B[159][3] +
                mat_A[5][0] * mat_B[167][3] +
                mat_A[5][1] * mat_B[175][3] +
                mat_A[5][2] * mat_B[183][3] +
                mat_A[5][3] * mat_B[191][3] +
                mat_A[6][0] * mat_B[199][3] +
                mat_A[6][1] * mat_B[207][3] +
                mat_A[6][2] * mat_B[215][3] +
                mat_A[6][3] * mat_B[223][3] +
                mat_A[7][0] * mat_B[231][3] +
                mat_A[7][1] * mat_B[239][3] +
                mat_A[7][2] * mat_B[247][3] +
                mat_A[7][3] * mat_B[255][3];
    mat_C[8][0] <=
                mat_A[8][0] * mat_B[0][0] +
                mat_A[8][1] * mat_B[8][0] +
                mat_A[8][2] * mat_B[16][0] +
                mat_A[8][3] * mat_B[24][0] +
                mat_A[9][0] * mat_B[32][0] +
                mat_A[9][1] * mat_B[40][0] +
                mat_A[9][2] * mat_B[48][0] +
                mat_A[9][3] * mat_B[56][0] +
                mat_A[10][0] * mat_B[64][0] +
                mat_A[10][1] * mat_B[72][0] +
                mat_A[10][2] * mat_B[80][0] +
                mat_A[10][3] * mat_B[88][0] +
                mat_A[11][0] * mat_B[96][0] +
                mat_A[11][1] * mat_B[104][0] +
                mat_A[11][2] * mat_B[112][0] +
                mat_A[11][3] * mat_B[120][0] +
                mat_A[12][0] * mat_B[128][0] +
                mat_A[12][1] * mat_B[136][0] +
                mat_A[12][2] * mat_B[144][0] +
                mat_A[12][3] * mat_B[152][0] +
                mat_A[13][0] * mat_B[160][0] +
                mat_A[13][1] * mat_B[168][0] +
                mat_A[13][2] * mat_B[176][0] +
                mat_A[13][3] * mat_B[184][0] +
                mat_A[14][0] * mat_B[192][0] +
                mat_A[14][1] * mat_B[200][0] +
                mat_A[14][2] * mat_B[208][0] +
                mat_A[14][3] * mat_B[216][0] +
                mat_A[15][0] * mat_B[224][0] +
                mat_A[15][1] * mat_B[232][0] +
                mat_A[15][2] * mat_B[240][0] +
                mat_A[15][3] * mat_B[248][0];
    mat_C[8][1] <=
                mat_A[8][0] * mat_B[0][1] +
                mat_A[8][1] * mat_B[8][1] +
                mat_A[8][2] * mat_B[16][1] +
                mat_A[8][3] * mat_B[24][1] +
                mat_A[9][0] * mat_B[32][1] +
                mat_A[9][1] * mat_B[40][1] +
                mat_A[9][2] * mat_B[48][1] +
                mat_A[9][3] * mat_B[56][1] +
                mat_A[10][0] * mat_B[64][1] +
                mat_A[10][1] * mat_B[72][1] +
                mat_A[10][2] * mat_B[80][1] +
                mat_A[10][3] * mat_B[88][1] +
                mat_A[11][0] * mat_B[96][1] +
                mat_A[11][1] * mat_B[104][1] +
                mat_A[11][2] * mat_B[112][1] +
                mat_A[11][3] * mat_B[120][1] +
                mat_A[12][0] * mat_B[128][1] +
                mat_A[12][1] * mat_B[136][1] +
                mat_A[12][2] * mat_B[144][1] +
                mat_A[12][3] * mat_B[152][1] +
                mat_A[13][0] * mat_B[160][1] +
                mat_A[13][1] * mat_B[168][1] +
                mat_A[13][2] * mat_B[176][1] +
                mat_A[13][3] * mat_B[184][1] +
                mat_A[14][0] * mat_B[192][1] +
                mat_A[14][1] * mat_B[200][1] +
                mat_A[14][2] * mat_B[208][1] +
                mat_A[14][3] * mat_B[216][1] +
                mat_A[15][0] * mat_B[224][1] +
                mat_A[15][1] * mat_B[232][1] +
                mat_A[15][2] * mat_B[240][1] +
                mat_A[15][3] * mat_B[248][1];
    mat_C[8][2] <=
                mat_A[8][0] * mat_B[0][2] +
                mat_A[8][1] * mat_B[8][2] +
                mat_A[8][2] * mat_B[16][2] +
                mat_A[8][3] * mat_B[24][2] +
                mat_A[9][0] * mat_B[32][2] +
                mat_A[9][1] * mat_B[40][2] +
                mat_A[9][2] * mat_B[48][2] +
                mat_A[9][3] * mat_B[56][2] +
                mat_A[10][0] * mat_B[64][2] +
                mat_A[10][1] * mat_B[72][2] +
                mat_A[10][2] * mat_B[80][2] +
                mat_A[10][3] * mat_B[88][2] +
                mat_A[11][0] * mat_B[96][2] +
                mat_A[11][1] * mat_B[104][2] +
                mat_A[11][2] * mat_B[112][2] +
                mat_A[11][3] * mat_B[120][2] +
                mat_A[12][0] * mat_B[128][2] +
                mat_A[12][1] * mat_B[136][2] +
                mat_A[12][2] * mat_B[144][2] +
                mat_A[12][3] * mat_B[152][2] +
                mat_A[13][0] * mat_B[160][2] +
                mat_A[13][1] * mat_B[168][2] +
                mat_A[13][2] * mat_B[176][2] +
                mat_A[13][3] * mat_B[184][2] +
                mat_A[14][0] * mat_B[192][2] +
                mat_A[14][1] * mat_B[200][2] +
                mat_A[14][2] * mat_B[208][2] +
                mat_A[14][3] * mat_B[216][2] +
                mat_A[15][0] * mat_B[224][2] +
                mat_A[15][1] * mat_B[232][2] +
                mat_A[15][2] * mat_B[240][2] +
                mat_A[15][3] * mat_B[248][2];
    mat_C[8][3] <=
                mat_A[8][0] * mat_B[0][3] +
                mat_A[8][1] * mat_B[8][3] +
                mat_A[8][2] * mat_B[16][3] +
                mat_A[8][3] * mat_B[24][3] +
                mat_A[9][0] * mat_B[32][3] +
                mat_A[9][1] * mat_B[40][3] +
                mat_A[9][2] * mat_B[48][3] +
                mat_A[9][3] * mat_B[56][3] +
                mat_A[10][0] * mat_B[64][3] +
                mat_A[10][1] * mat_B[72][3] +
                mat_A[10][2] * mat_B[80][3] +
                mat_A[10][3] * mat_B[88][3] +
                mat_A[11][0] * mat_B[96][3] +
                mat_A[11][1] * mat_B[104][3] +
                mat_A[11][2] * mat_B[112][3] +
                mat_A[11][3] * mat_B[120][3] +
                mat_A[12][0] * mat_B[128][3] +
                mat_A[12][1] * mat_B[136][3] +
                mat_A[12][2] * mat_B[144][3] +
                mat_A[12][3] * mat_B[152][3] +
                mat_A[13][0] * mat_B[160][3] +
                mat_A[13][1] * mat_B[168][3] +
                mat_A[13][2] * mat_B[176][3] +
                mat_A[13][3] * mat_B[184][3] +
                mat_A[14][0] * mat_B[192][3] +
                mat_A[14][1] * mat_B[200][3] +
                mat_A[14][2] * mat_B[208][3] +
                mat_A[14][3] * mat_B[216][3] +
                mat_A[15][0] * mat_B[224][3] +
                mat_A[15][1] * mat_B[232][3] +
                mat_A[15][2] * mat_B[240][3] +
                mat_A[15][3] * mat_B[248][3];
    mat_C[9][0] <=
                mat_A[8][0] * mat_B[1][0] +
                mat_A[8][1] * mat_B[9][0] +
                mat_A[8][2] * mat_B[17][0] +
                mat_A[8][3] * mat_B[25][0] +
                mat_A[9][0] * mat_B[33][0] +
                mat_A[9][1] * mat_B[41][0] +
                mat_A[9][2] * mat_B[49][0] +
                mat_A[9][3] * mat_B[57][0] +
                mat_A[10][0] * mat_B[65][0] +
                mat_A[10][1] * mat_B[73][0] +
                mat_A[10][2] * mat_B[81][0] +
                mat_A[10][3] * mat_B[89][0] +
                mat_A[11][0] * mat_B[97][0] +
                mat_A[11][1] * mat_B[105][0] +
                mat_A[11][2] * mat_B[113][0] +
                mat_A[11][3] * mat_B[121][0] +
                mat_A[12][0] * mat_B[129][0] +
                mat_A[12][1] * mat_B[137][0] +
                mat_A[12][2] * mat_B[145][0] +
                mat_A[12][3] * mat_B[153][0] +
                mat_A[13][0] * mat_B[161][0] +
                mat_A[13][1] * mat_B[169][0] +
                mat_A[13][2] * mat_B[177][0] +
                mat_A[13][3] * mat_B[185][0] +
                mat_A[14][0] * mat_B[193][0] +
                mat_A[14][1] * mat_B[201][0] +
                mat_A[14][2] * mat_B[209][0] +
                mat_A[14][3] * mat_B[217][0] +
                mat_A[15][0] * mat_B[225][0] +
                mat_A[15][1] * mat_B[233][0] +
                mat_A[15][2] * mat_B[241][0] +
                mat_A[15][3] * mat_B[249][0];
    mat_C[9][1] <=
                mat_A[8][0] * mat_B[1][1] +
                mat_A[8][1] * mat_B[9][1] +
                mat_A[8][2] * mat_B[17][1] +
                mat_A[8][3] * mat_B[25][1] +
                mat_A[9][0] * mat_B[33][1] +
                mat_A[9][1] * mat_B[41][1] +
                mat_A[9][2] * mat_B[49][1] +
                mat_A[9][3] * mat_B[57][1] +
                mat_A[10][0] * mat_B[65][1] +
                mat_A[10][1] * mat_B[73][1] +
                mat_A[10][2] * mat_B[81][1] +
                mat_A[10][3] * mat_B[89][1] +
                mat_A[11][0] * mat_B[97][1] +
                mat_A[11][1] * mat_B[105][1] +
                mat_A[11][2] * mat_B[113][1] +
                mat_A[11][3] * mat_B[121][1] +
                mat_A[12][0] * mat_B[129][1] +
                mat_A[12][1] * mat_B[137][1] +
                mat_A[12][2] * mat_B[145][1] +
                mat_A[12][3] * mat_B[153][1] +
                mat_A[13][0] * mat_B[161][1] +
                mat_A[13][1] * mat_B[169][1] +
                mat_A[13][2] * mat_B[177][1] +
                mat_A[13][3] * mat_B[185][1] +
                mat_A[14][0] * mat_B[193][1] +
                mat_A[14][1] * mat_B[201][1] +
                mat_A[14][2] * mat_B[209][1] +
                mat_A[14][3] * mat_B[217][1] +
                mat_A[15][0] * mat_B[225][1] +
                mat_A[15][1] * mat_B[233][1] +
                mat_A[15][2] * mat_B[241][1] +
                mat_A[15][3] * mat_B[249][1];
    mat_C[9][2] <=
                mat_A[8][0] * mat_B[1][2] +
                mat_A[8][1] * mat_B[9][2] +
                mat_A[8][2] * mat_B[17][2] +
                mat_A[8][3] * mat_B[25][2] +
                mat_A[9][0] * mat_B[33][2] +
                mat_A[9][1] * mat_B[41][2] +
                mat_A[9][2] * mat_B[49][2] +
                mat_A[9][3] * mat_B[57][2] +
                mat_A[10][0] * mat_B[65][2] +
                mat_A[10][1] * mat_B[73][2] +
                mat_A[10][2] * mat_B[81][2] +
                mat_A[10][3] * mat_B[89][2] +
                mat_A[11][0] * mat_B[97][2] +
                mat_A[11][1] * mat_B[105][2] +
                mat_A[11][2] * mat_B[113][2] +
                mat_A[11][3] * mat_B[121][2] +
                mat_A[12][0] * mat_B[129][2] +
                mat_A[12][1] * mat_B[137][2] +
                mat_A[12][2] * mat_B[145][2] +
                mat_A[12][3] * mat_B[153][2] +
                mat_A[13][0] * mat_B[161][2] +
                mat_A[13][1] * mat_B[169][2] +
                mat_A[13][2] * mat_B[177][2] +
                mat_A[13][3] * mat_B[185][2] +
                mat_A[14][0] * mat_B[193][2] +
                mat_A[14][1] * mat_B[201][2] +
                mat_A[14][2] * mat_B[209][2] +
                mat_A[14][3] * mat_B[217][2] +
                mat_A[15][0] * mat_B[225][2] +
                mat_A[15][1] * mat_B[233][2] +
                mat_A[15][2] * mat_B[241][2] +
                mat_A[15][3] * mat_B[249][2];
    mat_C[9][3] <=
                mat_A[8][0] * mat_B[1][3] +
                mat_A[8][1] * mat_B[9][3] +
                mat_A[8][2] * mat_B[17][3] +
                mat_A[8][3] * mat_B[25][3] +
                mat_A[9][0] * mat_B[33][3] +
                mat_A[9][1] * mat_B[41][3] +
                mat_A[9][2] * mat_B[49][3] +
                mat_A[9][3] * mat_B[57][3] +
                mat_A[10][0] * mat_B[65][3] +
                mat_A[10][1] * mat_B[73][3] +
                mat_A[10][2] * mat_B[81][3] +
                mat_A[10][3] * mat_B[89][3] +
                mat_A[11][0] * mat_B[97][3] +
                mat_A[11][1] * mat_B[105][3] +
                mat_A[11][2] * mat_B[113][3] +
                mat_A[11][3] * mat_B[121][3] +
                mat_A[12][0] * mat_B[129][3] +
                mat_A[12][1] * mat_B[137][3] +
                mat_A[12][2] * mat_B[145][3] +
                mat_A[12][3] * mat_B[153][3] +
                mat_A[13][0] * mat_B[161][3] +
                mat_A[13][1] * mat_B[169][3] +
                mat_A[13][2] * mat_B[177][3] +
                mat_A[13][3] * mat_B[185][3] +
                mat_A[14][0] * mat_B[193][3] +
                mat_A[14][1] * mat_B[201][3] +
                mat_A[14][2] * mat_B[209][3] +
                mat_A[14][3] * mat_B[217][3] +
                mat_A[15][0] * mat_B[225][3] +
                mat_A[15][1] * mat_B[233][3] +
                mat_A[15][2] * mat_B[241][3] +
                mat_A[15][3] * mat_B[249][3];
    mat_C[10][0] <=
                mat_A[8][0] * mat_B[2][0] +
                mat_A[8][1] * mat_B[10][0] +
                mat_A[8][2] * mat_B[18][0] +
                mat_A[8][3] * mat_B[26][0] +
                mat_A[9][0] * mat_B[34][0] +
                mat_A[9][1] * mat_B[42][0] +
                mat_A[9][2] * mat_B[50][0] +
                mat_A[9][3] * mat_B[58][0] +
                mat_A[10][0] * mat_B[66][0] +
                mat_A[10][1] * mat_B[74][0] +
                mat_A[10][2] * mat_B[82][0] +
                mat_A[10][3] * mat_B[90][0] +
                mat_A[11][0] * mat_B[98][0] +
                mat_A[11][1] * mat_B[106][0] +
                mat_A[11][2] * mat_B[114][0] +
                mat_A[11][3] * mat_B[122][0] +
                mat_A[12][0] * mat_B[130][0] +
                mat_A[12][1] * mat_B[138][0] +
                mat_A[12][2] * mat_B[146][0] +
                mat_A[12][3] * mat_B[154][0] +
                mat_A[13][0] * mat_B[162][0] +
                mat_A[13][1] * mat_B[170][0] +
                mat_A[13][2] * mat_B[178][0] +
                mat_A[13][3] * mat_B[186][0] +
                mat_A[14][0] * mat_B[194][0] +
                mat_A[14][1] * mat_B[202][0] +
                mat_A[14][2] * mat_B[210][0] +
                mat_A[14][3] * mat_B[218][0] +
                mat_A[15][0] * mat_B[226][0] +
                mat_A[15][1] * mat_B[234][0] +
                mat_A[15][2] * mat_B[242][0] +
                mat_A[15][3] * mat_B[250][0];
    mat_C[10][1] <=
                mat_A[8][0] * mat_B[2][1] +
                mat_A[8][1] * mat_B[10][1] +
                mat_A[8][2] * mat_B[18][1] +
                mat_A[8][3] * mat_B[26][1] +
                mat_A[9][0] * mat_B[34][1] +
                mat_A[9][1] * mat_B[42][1] +
                mat_A[9][2] * mat_B[50][1] +
                mat_A[9][3] * mat_B[58][1] +
                mat_A[10][0] * mat_B[66][1] +
                mat_A[10][1] * mat_B[74][1] +
                mat_A[10][2] * mat_B[82][1] +
                mat_A[10][3] * mat_B[90][1] +
                mat_A[11][0] * mat_B[98][1] +
                mat_A[11][1] * mat_B[106][1] +
                mat_A[11][2] * mat_B[114][1] +
                mat_A[11][3] * mat_B[122][1] +
                mat_A[12][0] * mat_B[130][1] +
                mat_A[12][1] * mat_B[138][1] +
                mat_A[12][2] * mat_B[146][1] +
                mat_A[12][3] * mat_B[154][1] +
                mat_A[13][0] * mat_B[162][1] +
                mat_A[13][1] * mat_B[170][1] +
                mat_A[13][2] * mat_B[178][1] +
                mat_A[13][3] * mat_B[186][1] +
                mat_A[14][0] * mat_B[194][1] +
                mat_A[14][1] * mat_B[202][1] +
                mat_A[14][2] * mat_B[210][1] +
                mat_A[14][3] * mat_B[218][1] +
                mat_A[15][0] * mat_B[226][1] +
                mat_A[15][1] * mat_B[234][1] +
                mat_A[15][2] * mat_B[242][1] +
                mat_A[15][3] * mat_B[250][1];
    mat_C[10][2] <=
                mat_A[8][0] * mat_B[2][2] +
                mat_A[8][1] * mat_B[10][2] +
                mat_A[8][2] * mat_B[18][2] +
                mat_A[8][3] * mat_B[26][2] +
                mat_A[9][0] * mat_B[34][2] +
                mat_A[9][1] * mat_B[42][2] +
                mat_A[9][2] * mat_B[50][2] +
                mat_A[9][3] * mat_B[58][2] +
                mat_A[10][0] * mat_B[66][2] +
                mat_A[10][1] * mat_B[74][2] +
                mat_A[10][2] * mat_B[82][2] +
                mat_A[10][3] * mat_B[90][2] +
                mat_A[11][0] * mat_B[98][2] +
                mat_A[11][1] * mat_B[106][2] +
                mat_A[11][2] * mat_B[114][2] +
                mat_A[11][3] * mat_B[122][2] +
                mat_A[12][0] * mat_B[130][2] +
                mat_A[12][1] * mat_B[138][2] +
                mat_A[12][2] * mat_B[146][2] +
                mat_A[12][3] * mat_B[154][2] +
                mat_A[13][0] * mat_B[162][2] +
                mat_A[13][1] * mat_B[170][2] +
                mat_A[13][2] * mat_B[178][2] +
                mat_A[13][3] * mat_B[186][2] +
                mat_A[14][0] * mat_B[194][2] +
                mat_A[14][1] * mat_B[202][2] +
                mat_A[14][2] * mat_B[210][2] +
                mat_A[14][3] * mat_B[218][2] +
                mat_A[15][0] * mat_B[226][2] +
                mat_A[15][1] * mat_B[234][2] +
                mat_A[15][2] * mat_B[242][2] +
                mat_A[15][3] * mat_B[250][2];
    mat_C[10][3] <=
                mat_A[8][0] * mat_B[2][3] +
                mat_A[8][1] * mat_B[10][3] +
                mat_A[8][2] * mat_B[18][3] +
                mat_A[8][3] * mat_B[26][3] +
                mat_A[9][0] * mat_B[34][3] +
                mat_A[9][1] * mat_B[42][3] +
                mat_A[9][2] * mat_B[50][3] +
                mat_A[9][3] * mat_B[58][3] +
                mat_A[10][0] * mat_B[66][3] +
                mat_A[10][1] * mat_B[74][3] +
                mat_A[10][2] * mat_B[82][3] +
                mat_A[10][3] * mat_B[90][3] +
                mat_A[11][0] * mat_B[98][3] +
                mat_A[11][1] * mat_B[106][3] +
                mat_A[11][2] * mat_B[114][3] +
                mat_A[11][3] * mat_B[122][3] +
                mat_A[12][0] * mat_B[130][3] +
                mat_A[12][1] * mat_B[138][3] +
                mat_A[12][2] * mat_B[146][3] +
                mat_A[12][3] * mat_B[154][3] +
                mat_A[13][0] * mat_B[162][3] +
                mat_A[13][1] * mat_B[170][3] +
                mat_A[13][2] * mat_B[178][3] +
                mat_A[13][3] * mat_B[186][3] +
                mat_A[14][0] * mat_B[194][3] +
                mat_A[14][1] * mat_B[202][3] +
                mat_A[14][2] * mat_B[210][3] +
                mat_A[14][3] * mat_B[218][3] +
                mat_A[15][0] * mat_B[226][3] +
                mat_A[15][1] * mat_B[234][3] +
                mat_A[15][2] * mat_B[242][3] +
                mat_A[15][3] * mat_B[250][3];
    mat_C[11][0] <=
                mat_A[8][0] * mat_B[3][0] +
                mat_A[8][1] * mat_B[11][0] +
                mat_A[8][2] * mat_B[19][0] +
                mat_A[8][3] * mat_B[27][0] +
                mat_A[9][0] * mat_B[35][0] +
                mat_A[9][1] * mat_B[43][0] +
                mat_A[9][2] * mat_B[51][0] +
                mat_A[9][3] * mat_B[59][0] +
                mat_A[10][0] * mat_B[67][0] +
                mat_A[10][1] * mat_B[75][0] +
                mat_A[10][2] * mat_B[83][0] +
                mat_A[10][3] * mat_B[91][0] +
                mat_A[11][0] * mat_B[99][0] +
                mat_A[11][1] * mat_B[107][0] +
                mat_A[11][2] * mat_B[115][0] +
                mat_A[11][3] * mat_B[123][0] +
                mat_A[12][0] * mat_B[131][0] +
                mat_A[12][1] * mat_B[139][0] +
                mat_A[12][2] * mat_B[147][0] +
                mat_A[12][3] * mat_B[155][0] +
                mat_A[13][0] * mat_B[163][0] +
                mat_A[13][1] * mat_B[171][0] +
                mat_A[13][2] * mat_B[179][0] +
                mat_A[13][3] * mat_B[187][0] +
                mat_A[14][0] * mat_B[195][0] +
                mat_A[14][1] * mat_B[203][0] +
                mat_A[14][2] * mat_B[211][0] +
                mat_A[14][3] * mat_B[219][0] +
                mat_A[15][0] * mat_B[227][0] +
                mat_A[15][1] * mat_B[235][0] +
                mat_A[15][2] * mat_B[243][0] +
                mat_A[15][3] * mat_B[251][0];
    mat_C[11][1] <=
                mat_A[8][0] * mat_B[3][1] +
                mat_A[8][1] * mat_B[11][1] +
                mat_A[8][2] * mat_B[19][1] +
                mat_A[8][3] * mat_B[27][1] +
                mat_A[9][0] * mat_B[35][1] +
                mat_A[9][1] * mat_B[43][1] +
                mat_A[9][2] * mat_B[51][1] +
                mat_A[9][3] * mat_B[59][1] +
                mat_A[10][0] * mat_B[67][1] +
                mat_A[10][1] * mat_B[75][1] +
                mat_A[10][2] * mat_B[83][1] +
                mat_A[10][3] * mat_B[91][1] +
                mat_A[11][0] * mat_B[99][1] +
                mat_A[11][1] * mat_B[107][1] +
                mat_A[11][2] * mat_B[115][1] +
                mat_A[11][3] * mat_B[123][1] +
                mat_A[12][0] * mat_B[131][1] +
                mat_A[12][1] * mat_B[139][1] +
                mat_A[12][2] * mat_B[147][1] +
                mat_A[12][3] * mat_B[155][1] +
                mat_A[13][0] * mat_B[163][1] +
                mat_A[13][1] * mat_B[171][1] +
                mat_A[13][2] * mat_B[179][1] +
                mat_A[13][3] * mat_B[187][1] +
                mat_A[14][0] * mat_B[195][1] +
                mat_A[14][1] * mat_B[203][1] +
                mat_A[14][2] * mat_B[211][1] +
                mat_A[14][3] * mat_B[219][1] +
                mat_A[15][0] * mat_B[227][1] +
                mat_A[15][1] * mat_B[235][1] +
                mat_A[15][2] * mat_B[243][1] +
                mat_A[15][3] * mat_B[251][1];
    mat_C[11][2] <=
                mat_A[8][0] * mat_B[3][2] +
                mat_A[8][1] * mat_B[11][2] +
                mat_A[8][2] * mat_B[19][2] +
                mat_A[8][3] * mat_B[27][2] +
                mat_A[9][0] * mat_B[35][2] +
                mat_A[9][1] * mat_B[43][2] +
                mat_A[9][2] * mat_B[51][2] +
                mat_A[9][3] * mat_B[59][2] +
                mat_A[10][0] * mat_B[67][2] +
                mat_A[10][1] * mat_B[75][2] +
                mat_A[10][2] * mat_B[83][2] +
                mat_A[10][3] * mat_B[91][2] +
                mat_A[11][0] * mat_B[99][2] +
                mat_A[11][1] * mat_B[107][2] +
                mat_A[11][2] * mat_B[115][2] +
                mat_A[11][3] * mat_B[123][2] +
                mat_A[12][0] * mat_B[131][2] +
                mat_A[12][1] * mat_B[139][2] +
                mat_A[12][2] * mat_B[147][2] +
                mat_A[12][3] * mat_B[155][2] +
                mat_A[13][0] * mat_B[163][2] +
                mat_A[13][1] * mat_B[171][2] +
                mat_A[13][2] * mat_B[179][2] +
                mat_A[13][3] * mat_B[187][2] +
                mat_A[14][0] * mat_B[195][2] +
                mat_A[14][1] * mat_B[203][2] +
                mat_A[14][2] * mat_B[211][2] +
                mat_A[14][3] * mat_B[219][2] +
                mat_A[15][0] * mat_B[227][2] +
                mat_A[15][1] * mat_B[235][2] +
                mat_A[15][2] * mat_B[243][2] +
                mat_A[15][3] * mat_B[251][2];
    mat_C[11][3] <=
                mat_A[8][0] * mat_B[3][3] +
                mat_A[8][1] * mat_B[11][3] +
                mat_A[8][2] * mat_B[19][3] +
                mat_A[8][3] * mat_B[27][3] +
                mat_A[9][0] * mat_B[35][3] +
                mat_A[9][1] * mat_B[43][3] +
                mat_A[9][2] * mat_B[51][3] +
                mat_A[9][3] * mat_B[59][3] +
                mat_A[10][0] * mat_B[67][3] +
                mat_A[10][1] * mat_B[75][3] +
                mat_A[10][2] * mat_B[83][3] +
                mat_A[10][3] * mat_B[91][3] +
                mat_A[11][0] * mat_B[99][3] +
                mat_A[11][1] * mat_B[107][3] +
                mat_A[11][2] * mat_B[115][3] +
                mat_A[11][3] * mat_B[123][3] +
                mat_A[12][0] * mat_B[131][3] +
                mat_A[12][1] * mat_B[139][3] +
                mat_A[12][2] * mat_B[147][3] +
                mat_A[12][3] * mat_B[155][3] +
                mat_A[13][0] * mat_B[163][3] +
                mat_A[13][1] * mat_B[171][3] +
                mat_A[13][2] * mat_B[179][3] +
                mat_A[13][3] * mat_B[187][3] +
                mat_A[14][0] * mat_B[195][3] +
                mat_A[14][1] * mat_B[203][3] +
                mat_A[14][2] * mat_B[211][3] +
                mat_A[14][3] * mat_B[219][3] +
                mat_A[15][0] * mat_B[227][3] +
                mat_A[15][1] * mat_B[235][3] +
                mat_A[15][2] * mat_B[243][3] +
                mat_A[15][3] * mat_B[251][3];
    mat_C[12][0] <=
                mat_A[8][0] * mat_B[4][0] +
                mat_A[8][1] * mat_B[12][0] +
                mat_A[8][2] * mat_B[20][0] +
                mat_A[8][3] * mat_B[28][0] +
                mat_A[9][0] * mat_B[36][0] +
                mat_A[9][1] * mat_B[44][0] +
                mat_A[9][2] * mat_B[52][0] +
                mat_A[9][3] * mat_B[60][0] +
                mat_A[10][0] * mat_B[68][0] +
                mat_A[10][1] * mat_B[76][0] +
                mat_A[10][2] * mat_B[84][0] +
                mat_A[10][3] * mat_B[92][0] +
                mat_A[11][0] * mat_B[100][0] +
                mat_A[11][1] * mat_B[108][0] +
                mat_A[11][2] * mat_B[116][0] +
                mat_A[11][3] * mat_B[124][0] +
                mat_A[12][0] * mat_B[132][0] +
                mat_A[12][1] * mat_B[140][0] +
                mat_A[12][2] * mat_B[148][0] +
                mat_A[12][3] * mat_B[156][0] +
                mat_A[13][0] * mat_B[164][0] +
                mat_A[13][1] * mat_B[172][0] +
                mat_A[13][2] * mat_B[180][0] +
                mat_A[13][3] * mat_B[188][0] +
                mat_A[14][0] * mat_B[196][0] +
                mat_A[14][1] * mat_B[204][0] +
                mat_A[14][2] * mat_B[212][0] +
                mat_A[14][3] * mat_B[220][0] +
                mat_A[15][0] * mat_B[228][0] +
                mat_A[15][1] * mat_B[236][0] +
                mat_A[15][2] * mat_B[244][0] +
                mat_A[15][3] * mat_B[252][0];
    mat_C[12][1] <=
                mat_A[8][0] * mat_B[4][1] +
                mat_A[8][1] * mat_B[12][1] +
                mat_A[8][2] * mat_B[20][1] +
                mat_A[8][3] * mat_B[28][1] +
                mat_A[9][0] * mat_B[36][1] +
                mat_A[9][1] * mat_B[44][1] +
                mat_A[9][2] * mat_B[52][1] +
                mat_A[9][3] * mat_B[60][1] +
                mat_A[10][0] * mat_B[68][1] +
                mat_A[10][1] * mat_B[76][1] +
                mat_A[10][2] * mat_B[84][1] +
                mat_A[10][3] * mat_B[92][1] +
                mat_A[11][0] * mat_B[100][1] +
                mat_A[11][1] * mat_B[108][1] +
                mat_A[11][2] * mat_B[116][1] +
                mat_A[11][3] * mat_B[124][1] +
                mat_A[12][0] * mat_B[132][1] +
                mat_A[12][1] * mat_B[140][1] +
                mat_A[12][2] * mat_B[148][1] +
                mat_A[12][3] * mat_B[156][1] +
                mat_A[13][0] * mat_B[164][1] +
                mat_A[13][1] * mat_B[172][1] +
                mat_A[13][2] * mat_B[180][1] +
                mat_A[13][3] * mat_B[188][1] +
                mat_A[14][0] * mat_B[196][1] +
                mat_A[14][1] * mat_B[204][1] +
                mat_A[14][2] * mat_B[212][1] +
                mat_A[14][3] * mat_B[220][1] +
                mat_A[15][0] * mat_B[228][1] +
                mat_A[15][1] * mat_B[236][1] +
                mat_A[15][2] * mat_B[244][1] +
                mat_A[15][3] * mat_B[252][1];
    mat_C[12][2] <=
                mat_A[8][0] * mat_B[4][2] +
                mat_A[8][1] * mat_B[12][2] +
                mat_A[8][2] * mat_B[20][2] +
                mat_A[8][3] * mat_B[28][2] +
                mat_A[9][0] * mat_B[36][2] +
                mat_A[9][1] * mat_B[44][2] +
                mat_A[9][2] * mat_B[52][2] +
                mat_A[9][3] * mat_B[60][2] +
                mat_A[10][0] * mat_B[68][2] +
                mat_A[10][1] * mat_B[76][2] +
                mat_A[10][2] * mat_B[84][2] +
                mat_A[10][3] * mat_B[92][2] +
                mat_A[11][0] * mat_B[100][2] +
                mat_A[11][1] * mat_B[108][2] +
                mat_A[11][2] * mat_B[116][2] +
                mat_A[11][3] * mat_B[124][2] +
                mat_A[12][0] * mat_B[132][2] +
                mat_A[12][1] * mat_B[140][2] +
                mat_A[12][2] * mat_B[148][2] +
                mat_A[12][3] * mat_B[156][2] +
                mat_A[13][0] * mat_B[164][2] +
                mat_A[13][1] * mat_B[172][2] +
                mat_A[13][2] * mat_B[180][2] +
                mat_A[13][3] * mat_B[188][2] +
                mat_A[14][0] * mat_B[196][2] +
                mat_A[14][1] * mat_B[204][2] +
                mat_A[14][2] * mat_B[212][2] +
                mat_A[14][3] * mat_B[220][2] +
                mat_A[15][0] * mat_B[228][2] +
                mat_A[15][1] * mat_B[236][2] +
                mat_A[15][2] * mat_B[244][2] +
                mat_A[15][3] * mat_B[252][2];
    mat_C[12][3] <=
                mat_A[8][0] * mat_B[4][3] +
                mat_A[8][1] * mat_B[12][3] +
                mat_A[8][2] * mat_B[20][3] +
                mat_A[8][3] * mat_B[28][3] +
                mat_A[9][0] * mat_B[36][3] +
                mat_A[9][1] * mat_B[44][3] +
                mat_A[9][2] * mat_B[52][3] +
                mat_A[9][3] * mat_B[60][3] +
                mat_A[10][0] * mat_B[68][3] +
                mat_A[10][1] * mat_B[76][3] +
                mat_A[10][2] * mat_B[84][3] +
                mat_A[10][3] * mat_B[92][3] +
                mat_A[11][0] * mat_B[100][3] +
                mat_A[11][1] * mat_B[108][3] +
                mat_A[11][2] * mat_B[116][3] +
                mat_A[11][3] * mat_B[124][3] +
                mat_A[12][0] * mat_B[132][3] +
                mat_A[12][1] * mat_B[140][3] +
                mat_A[12][2] * mat_B[148][3] +
                mat_A[12][3] * mat_B[156][3] +
                mat_A[13][0] * mat_B[164][3] +
                mat_A[13][1] * mat_B[172][3] +
                mat_A[13][2] * mat_B[180][3] +
                mat_A[13][3] * mat_B[188][3] +
                mat_A[14][0] * mat_B[196][3] +
                mat_A[14][1] * mat_B[204][3] +
                mat_A[14][2] * mat_B[212][3] +
                mat_A[14][3] * mat_B[220][3] +
                mat_A[15][0] * mat_B[228][3] +
                mat_A[15][1] * mat_B[236][3] +
                mat_A[15][2] * mat_B[244][3] +
                mat_A[15][3] * mat_B[252][3];
    mat_C[13][0] <=
                mat_A[8][0] * mat_B[5][0] +
                mat_A[8][1] * mat_B[13][0] +
                mat_A[8][2] * mat_B[21][0] +
                mat_A[8][3] * mat_B[29][0] +
                mat_A[9][0] * mat_B[37][0] +
                mat_A[9][1] * mat_B[45][0] +
                mat_A[9][2] * mat_B[53][0] +
                mat_A[9][3] * mat_B[61][0] +
                mat_A[10][0] * mat_B[69][0] +
                mat_A[10][1] * mat_B[77][0] +
                mat_A[10][2] * mat_B[85][0] +
                mat_A[10][3] * mat_B[93][0] +
                mat_A[11][0] * mat_B[101][0] +
                mat_A[11][1] * mat_B[109][0] +
                mat_A[11][2] * mat_B[117][0] +
                mat_A[11][3] * mat_B[125][0] +
                mat_A[12][0] * mat_B[133][0] +
                mat_A[12][1] * mat_B[141][0] +
                mat_A[12][2] * mat_B[149][0] +
                mat_A[12][3] * mat_B[157][0] +
                mat_A[13][0] * mat_B[165][0] +
                mat_A[13][1] * mat_B[173][0] +
                mat_A[13][2] * mat_B[181][0] +
                mat_A[13][3] * mat_B[189][0] +
                mat_A[14][0] * mat_B[197][0] +
                mat_A[14][1] * mat_B[205][0] +
                mat_A[14][2] * mat_B[213][0] +
                mat_A[14][3] * mat_B[221][0] +
                mat_A[15][0] * mat_B[229][0] +
                mat_A[15][1] * mat_B[237][0] +
                mat_A[15][2] * mat_B[245][0] +
                mat_A[15][3] * mat_B[253][0];
    mat_C[13][1] <=
                mat_A[8][0] * mat_B[5][1] +
                mat_A[8][1] * mat_B[13][1] +
                mat_A[8][2] * mat_B[21][1] +
                mat_A[8][3] * mat_B[29][1] +
                mat_A[9][0] * mat_B[37][1] +
                mat_A[9][1] * mat_B[45][1] +
                mat_A[9][2] * mat_B[53][1] +
                mat_A[9][3] * mat_B[61][1] +
                mat_A[10][0] * mat_B[69][1] +
                mat_A[10][1] * mat_B[77][1] +
                mat_A[10][2] * mat_B[85][1] +
                mat_A[10][3] * mat_B[93][1] +
                mat_A[11][0] * mat_B[101][1] +
                mat_A[11][1] * mat_B[109][1] +
                mat_A[11][2] * mat_B[117][1] +
                mat_A[11][3] * mat_B[125][1] +
                mat_A[12][0] * mat_B[133][1] +
                mat_A[12][1] * mat_B[141][1] +
                mat_A[12][2] * mat_B[149][1] +
                mat_A[12][3] * mat_B[157][1] +
                mat_A[13][0] * mat_B[165][1] +
                mat_A[13][1] * mat_B[173][1] +
                mat_A[13][2] * mat_B[181][1] +
                mat_A[13][3] * mat_B[189][1] +
                mat_A[14][0] * mat_B[197][1] +
                mat_A[14][1] * mat_B[205][1] +
                mat_A[14][2] * mat_B[213][1] +
                mat_A[14][3] * mat_B[221][1] +
                mat_A[15][0] * mat_B[229][1] +
                mat_A[15][1] * mat_B[237][1] +
                mat_A[15][2] * mat_B[245][1] +
                mat_A[15][3] * mat_B[253][1];
    mat_C[13][2] <=
                mat_A[8][0] * mat_B[5][2] +
                mat_A[8][1] * mat_B[13][2] +
                mat_A[8][2] * mat_B[21][2] +
                mat_A[8][3] * mat_B[29][2] +
                mat_A[9][0] * mat_B[37][2] +
                mat_A[9][1] * mat_B[45][2] +
                mat_A[9][2] * mat_B[53][2] +
                mat_A[9][3] * mat_B[61][2] +
                mat_A[10][0] * mat_B[69][2] +
                mat_A[10][1] * mat_B[77][2] +
                mat_A[10][2] * mat_B[85][2] +
                mat_A[10][3] * mat_B[93][2] +
                mat_A[11][0] * mat_B[101][2] +
                mat_A[11][1] * mat_B[109][2] +
                mat_A[11][2] * mat_B[117][2] +
                mat_A[11][3] * mat_B[125][2] +
                mat_A[12][0] * mat_B[133][2] +
                mat_A[12][1] * mat_B[141][2] +
                mat_A[12][2] * mat_B[149][2] +
                mat_A[12][3] * mat_B[157][2] +
                mat_A[13][0] * mat_B[165][2] +
                mat_A[13][1] * mat_B[173][2] +
                mat_A[13][2] * mat_B[181][2] +
                mat_A[13][3] * mat_B[189][2] +
                mat_A[14][0] * mat_B[197][2] +
                mat_A[14][1] * mat_B[205][2] +
                mat_A[14][2] * mat_B[213][2] +
                mat_A[14][3] * mat_B[221][2] +
                mat_A[15][0] * mat_B[229][2] +
                mat_A[15][1] * mat_B[237][2] +
                mat_A[15][2] * mat_B[245][2] +
                mat_A[15][3] * mat_B[253][2];
    mat_C[13][3] <=
                mat_A[8][0] * mat_B[5][3] +
                mat_A[8][1] * mat_B[13][3] +
                mat_A[8][2] * mat_B[21][3] +
                mat_A[8][3] * mat_B[29][3] +
                mat_A[9][0] * mat_B[37][3] +
                mat_A[9][1] * mat_B[45][3] +
                mat_A[9][2] * mat_B[53][3] +
                mat_A[9][3] * mat_B[61][3] +
                mat_A[10][0] * mat_B[69][3] +
                mat_A[10][1] * mat_B[77][3] +
                mat_A[10][2] * mat_B[85][3] +
                mat_A[10][3] * mat_B[93][3] +
                mat_A[11][0] * mat_B[101][3] +
                mat_A[11][1] * mat_B[109][3] +
                mat_A[11][2] * mat_B[117][3] +
                mat_A[11][3] * mat_B[125][3] +
                mat_A[12][0] * mat_B[133][3] +
                mat_A[12][1] * mat_B[141][3] +
                mat_A[12][2] * mat_B[149][3] +
                mat_A[12][3] * mat_B[157][3] +
                mat_A[13][0] * mat_B[165][3] +
                mat_A[13][1] * mat_B[173][3] +
                mat_A[13][2] * mat_B[181][3] +
                mat_A[13][3] * mat_B[189][3] +
                mat_A[14][0] * mat_B[197][3] +
                mat_A[14][1] * mat_B[205][3] +
                mat_A[14][2] * mat_B[213][3] +
                mat_A[14][3] * mat_B[221][3] +
                mat_A[15][0] * mat_B[229][3] +
                mat_A[15][1] * mat_B[237][3] +
                mat_A[15][2] * mat_B[245][3] +
                mat_A[15][3] * mat_B[253][3];
    mat_C[14][0] <=
                mat_A[8][0] * mat_B[6][0] +
                mat_A[8][1] * mat_B[14][0] +
                mat_A[8][2] * mat_B[22][0] +
                mat_A[8][3] * mat_B[30][0] +
                mat_A[9][0] * mat_B[38][0] +
                mat_A[9][1] * mat_B[46][0] +
                mat_A[9][2] * mat_B[54][0] +
                mat_A[9][3] * mat_B[62][0] +
                mat_A[10][0] * mat_B[70][0] +
                mat_A[10][1] * mat_B[78][0] +
                mat_A[10][2] * mat_B[86][0] +
                mat_A[10][3] * mat_B[94][0] +
                mat_A[11][0] * mat_B[102][0] +
                mat_A[11][1] * mat_B[110][0] +
                mat_A[11][2] * mat_B[118][0] +
                mat_A[11][3] * mat_B[126][0] +
                mat_A[12][0] * mat_B[134][0] +
                mat_A[12][1] * mat_B[142][0] +
                mat_A[12][2] * mat_B[150][0] +
                mat_A[12][3] * mat_B[158][0] +
                mat_A[13][0] * mat_B[166][0] +
                mat_A[13][1] * mat_B[174][0] +
                mat_A[13][2] * mat_B[182][0] +
                mat_A[13][3] * mat_B[190][0] +
                mat_A[14][0] * mat_B[198][0] +
                mat_A[14][1] * mat_B[206][0] +
                mat_A[14][2] * mat_B[214][0] +
                mat_A[14][3] * mat_B[222][0] +
                mat_A[15][0] * mat_B[230][0] +
                mat_A[15][1] * mat_B[238][0] +
                mat_A[15][2] * mat_B[246][0] +
                mat_A[15][3] * mat_B[254][0];
    mat_C[14][1] <=
                mat_A[8][0] * mat_B[6][1] +
                mat_A[8][1] * mat_B[14][1] +
                mat_A[8][2] * mat_B[22][1] +
                mat_A[8][3] * mat_B[30][1] +
                mat_A[9][0] * mat_B[38][1] +
                mat_A[9][1] * mat_B[46][1] +
                mat_A[9][2] * mat_B[54][1] +
                mat_A[9][3] * mat_B[62][1] +
                mat_A[10][0] * mat_B[70][1] +
                mat_A[10][1] * mat_B[78][1] +
                mat_A[10][2] * mat_B[86][1] +
                mat_A[10][3] * mat_B[94][1] +
                mat_A[11][0] * mat_B[102][1] +
                mat_A[11][1] * mat_B[110][1] +
                mat_A[11][2] * mat_B[118][1] +
                mat_A[11][3] * mat_B[126][1] +
                mat_A[12][0] * mat_B[134][1] +
                mat_A[12][1] * mat_B[142][1] +
                mat_A[12][2] * mat_B[150][1] +
                mat_A[12][3] * mat_B[158][1] +
                mat_A[13][0] * mat_B[166][1] +
                mat_A[13][1] * mat_B[174][1] +
                mat_A[13][2] * mat_B[182][1] +
                mat_A[13][3] * mat_B[190][1] +
                mat_A[14][0] * mat_B[198][1] +
                mat_A[14][1] * mat_B[206][1] +
                mat_A[14][2] * mat_B[214][1] +
                mat_A[14][3] * mat_B[222][1] +
                mat_A[15][0] * mat_B[230][1] +
                mat_A[15][1] * mat_B[238][1] +
                mat_A[15][2] * mat_B[246][1] +
                mat_A[15][3] * mat_B[254][1];
    mat_C[14][2] <=
                mat_A[8][0] * mat_B[6][2] +
                mat_A[8][1] * mat_B[14][2] +
                mat_A[8][2] * mat_B[22][2] +
                mat_A[8][3] * mat_B[30][2] +
                mat_A[9][0] * mat_B[38][2] +
                mat_A[9][1] * mat_B[46][2] +
                mat_A[9][2] * mat_B[54][2] +
                mat_A[9][3] * mat_B[62][2] +
                mat_A[10][0] * mat_B[70][2] +
                mat_A[10][1] * mat_B[78][2] +
                mat_A[10][2] * mat_B[86][2] +
                mat_A[10][3] * mat_B[94][2] +
                mat_A[11][0] * mat_B[102][2] +
                mat_A[11][1] * mat_B[110][2] +
                mat_A[11][2] * mat_B[118][2] +
                mat_A[11][3] * mat_B[126][2] +
                mat_A[12][0] * mat_B[134][2] +
                mat_A[12][1] * mat_B[142][2] +
                mat_A[12][2] * mat_B[150][2] +
                mat_A[12][3] * mat_B[158][2] +
                mat_A[13][0] * mat_B[166][2] +
                mat_A[13][1] * mat_B[174][2] +
                mat_A[13][2] * mat_B[182][2] +
                mat_A[13][3] * mat_B[190][2] +
                mat_A[14][0] * mat_B[198][2] +
                mat_A[14][1] * mat_B[206][2] +
                mat_A[14][2] * mat_B[214][2] +
                mat_A[14][3] * mat_B[222][2] +
                mat_A[15][0] * mat_B[230][2] +
                mat_A[15][1] * mat_B[238][2] +
                mat_A[15][2] * mat_B[246][2] +
                mat_A[15][3] * mat_B[254][2];
    mat_C[14][3] <=
                mat_A[8][0] * mat_B[6][3] +
                mat_A[8][1] * mat_B[14][3] +
                mat_A[8][2] * mat_B[22][3] +
                mat_A[8][3] * mat_B[30][3] +
                mat_A[9][0] * mat_B[38][3] +
                mat_A[9][1] * mat_B[46][3] +
                mat_A[9][2] * mat_B[54][3] +
                mat_A[9][3] * mat_B[62][3] +
                mat_A[10][0] * mat_B[70][3] +
                mat_A[10][1] * mat_B[78][3] +
                mat_A[10][2] * mat_B[86][3] +
                mat_A[10][3] * mat_B[94][3] +
                mat_A[11][0] * mat_B[102][3] +
                mat_A[11][1] * mat_B[110][3] +
                mat_A[11][2] * mat_B[118][3] +
                mat_A[11][3] * mat_B[126][3] +
                mat_A[12][0] * mat_B[134][3] +
                mat_A[12][1] * mat_B[142][3] +
                mat_A[12][2] * mat_B[150][3] +
                mat_A[12][3] * mat_B[158][3] +
                mat_A[13][0] * mat_B[166][3] +
                mat_A[13][1] * mat_B[174][3] +
                mat_A[13][2] * mat_B[182][3] +
                mat_A[13][3] * mat_B[190][3] +
                mat_A[14][0] * mat_B[198][3] +
                mat_A[14][1] * mat_B[206][3] +
                mat_A[14][2] * mat_B[214][3] +
                mat_A[14][3] * mat_B[222][3] +
                mat_A[15][0] * mat_B[230][3] +
                mat_A[15][1] * mat_B[238][3] +
                mat_A[15][2] * mat_B[246][3] +
                mat_A[15][3] * mat_B[254][3];
    mat_C[15][0] <=
                mat_A[8][0] * mat_B[7][0] +
                mat_A[8][1] * mat_B[15][0] +
                mat_A[8][2] * mat_B[23][0] +
                mat_A[8][3] * mat_B[31][0] +
                mat_A[9][0] * mat_B[39][0] +
                mat_A[9][1] * mat_B[47][0] +
                mat_A[9][2] * mat_B[55][0] +
                mat_A[9][3] * mat_B[63][0] +
                mat_A[10][0] * mat_B[71][0] +
                mat_A[10][1] * mat_B[79][0] +
                mat_A[10][2] * mat_B[87][0] +
                mat_A[10][3] * mat_B[95][0] +
                mat_A[11][0] * mat_B[103][0] +
                mat_A[11][1] * mat_B[111][0] +
                mat_A[11][2] * mat_B[119][0] +
                mat_A[11][3] * mat_B[127][0] +
                mat_A[12][0] * mat_B[135][0] +
                mat_A[12][1] * mat_B[143][0] +
                mat_A[12][2] * mat_B[151][0] +
                mat_A[12][3] * mat_B[159][0] +
                mat_A[13][0] * mat_B[167][0] +
                mat_A[13][1] * mat_B[175][0] +
                mat_A[13][2] * mat_B[183][0] +
                mat_A[13][3] * mat_B[191][0] +
                mat_A[14][0] * mat_B[199][0] +
                mat_A[14][1] * mat_B[207][0] +
                mat_A[14][2] * mat_B[215][0] +
                mat_A[14][3] * mat_B[223][0] +
                mat_A[15][0] * mat_B[231][0] +
                mat_A[15][1] * mat_B[239][0] +
                mat_A[15][2] * mat_B[247][0] +
                mat_A[15][3] * mat_B[255][0];
    mat_C[15][1] <=
                mat_A[8][0] * mat_B[7][1] +
                mat_A[8][1] * mat_B[15][1] +
                mat_A[8][2] * mat_B[23][1] +
                mat_A[8][3] * mat_B[31][1] +
                mat_A[9][0] * mat_B[39][1] +
                mat_A[9][1] * mat_B[47][1] +
                mat_A[9][2] * mat_B[55][1] +
                mat_A[9][3] * mat_B[63][1] +
                mat_A[10][0] * mat_B[71][1] +
                mat_A[10][1] * mat_B[79][1] +
                mat_A[10][2] * mat_B[87][1] +
                mat_A[10][3] * mat_B[95][1] +
                mat_A[11][0] * mat_B[103][1] +
                mat_A[11][1] * mat_B[111][1] +
                mat_A[11][2] * mat_B[119][1] +
                mat_A[11][3] * mat_B[127][1] +
                mat_A[12][0] * mat_B[135][1] +
                mat_A[12][1] * mat_B[143][1] +
                mat_A[12][2] * mat_B[151][1] +
                mat_A[12][3] * mat_B[159][1] +
                mat_A[13][0] * mat_B[167][1] +
                mat_A[13][1] * mat_B[175][1] +
                mat_A[13][2] * mat_B[183][1] +
                mat_A[13][3] * mat_B[191][1] +
                mat_A[14][0] * mat_B[199][1] +
                mat_A[14][1] * mat_B[207][1] +
                mat_A[14][2] * mat_B[215][1] +
                mat_A[14][3] * mat_B[223][1] +
                mat_A[15][0] * mat_B[231][1] +
                mat_A[15][1] * mat_B[239][1] +
                mat_A[15][2] * mat_B[247][1] +
                mat_A[15][3] * mat_B[255][1];
    mat_C[15][2] <=
                mat_A[8][0] * mat_B[7][2] +
                mat_A[8][1] * mat_B[15][2] +
                mat_A[8][2] * mat_B[23][2] +
                mat_A[8][3] * mat_B[31][2] +
                mat_A[9][0] * mat_B[39][2] +
                mat_A[9][1] * mat_B[47][2] +
                mat_A[9][2] * mat_B[55][2] +
                mat_A[9][3] * mat_B[63][2] +
                mat_A[10][0] * mat_B[71][2] +
                mat_A[10][1] * mat_B[79][2] +
                mat_A[10][2] * mat_B[87][2] +
                mat_A[10][3] * mat_B[95][2] +
                mat_A[11][0] * mat_B[103][2] +
                mat_A[11][1] * mat_B[111][2] +
                mat_A[11][2] * mat_B[119][2] +
                mat_A[11][3] * mat_B[127][2] +
                mat_A[12][0] * mat_B[135][2] +
                mat_A[12][1] * mat_B[143][2] +
                mat_A[12][2] * mat_B[151][2] +
                mat_A[12][3] * mat_B[159][2] +
                mat_A[13][0] * mat_B[167][2] +
                mat_A[13][1] * mat_B[175][2] +
                mat_A[13][2] * mat_B[183][2] +
                mat_A[13][3] * mat_B[191][2] +
                mat_A[14][0] * mat_B[199][2] +
                mat_A[14][1] * mat_B[207][2] +
                mat_A[14][2] * mat_B[215][2] +
                mat_A[14][3] * mat_B[223][2] +
                mat_A[15][0] * mat_B[231][2] +
                mat_A[15][1] * mat_B[239][2] +
                mat_A[15][2] * mat_B[247][2] +
                mat_A[15][3] * mat_B[255][2];
    mat_C[15][3] <=
                mat_A[8][0] * mat_B[7][3] +
                mat_A[8][1] * mat_B[15][3] +
                mat_A[8][2] * mat_B[23][3] +
                mat_A[8][3] * mat_B[31][3] +
                mat_A[9][0] * mat_B[39][3] +
                mat_A[9][1] * mat_B[47][3] +
                mat_A[9][2] * mat_B[55][3] +
                mat_A[9][3] * mat_B[63][3] +
                mat_A[10][0] * mat_B[71][3] +
                mat_A[10][1] * mat_B[79][3] +
                mat_A[10][2] * mat_B[87][3] +
                mat_A[10][3] * mat_B[95][3] +
                mat_A[11][0] * mat_B[103][3] +
                mat_A[11][1] * mat_B[111][3] +
                mat_A[11][2] * mat_B[119][3] +
                mat_A[11][3] * mat_B[127][3] +
                mat_A[12][0] * mat_B[135][3] +
                mat_A[12][1] * mat_B[143][3] +
                mat_A[12][2] * mat_B[151][3] +
                mat_A[12][3] * mat_B[159][3] +
                mat_A[13][0] * mat_B[167][3] +
                mat_A[13][1] * mat_B[175][3] +
                mat_A[13][2] * mat_B[183][3] +
                mat_A[13][3] * mat_B[191][3] +
                mat_A[14][0] * mat_B[199][3] +
                mat_A[14][1] * mat_B[207][3] +
                mat_A[14][2] * mat_B[215][3] +
                mat_A[14][3] * mat_B[223][3] +
                mat_A[15][0] * mat_B[231][3] +
                mat_A[15][1] * mat_B[239][3] +
                mat_A[15][2] * mat_B[247][3] +
                mat_A[15][3] * mat_B[255][3];
    mat_C[16][0] <=
                mat_A[16][0] * mat_B[0][0] +
                mat_A[16][1] * mat_B[8][0] +
                mat_A[16][2] * mat_B[16][0] +
                mat_A[16][3] * mat_B[24][0] +
                mat_A[17][0] * mat_B[32][0] +
                mat_A[17][1] * mat_B[40][0] +
                mat_A[17][2] * mat_B[48][0] +
                mat_A[17][3] * mat_B[56][0] +
                mat_A[18][0] * mat_B[64][0] +
                mat_A[18][1] * mat_B[72][0] +
                mat_A[18][2] * mat_B[80][0] +
                mat_A[18][3] * mat_B[88][0] +
                mat_A[19][0] * mat_B[96][0] +
                mat_A[19][1] * mat_B[104][0] +
                mat_A[19][2] * mat_B[112][0] +
                mat_A[19][3] * mat_B[120][0] +
                mat_A[20][0] * mat_B[128][0] +
                mat_A[20][1] * mat_B[136][0] +
                mat_A[20][2] * mat_B[144][0] +
                mat_A[20][3] * mat_B[152][0] +
                mat_A[21][0] * mat_B[160][0] +
                mat_A[21][1] * mat_B[168][0] +
                mat_A[21][2] * mat_B[176][0] +
                mat_A[21][3] * mat_B[184][0] +
                mat_A[22][0] * mat_B[192][0] +
                mat_A[22][1] * mat_B[200][0] +
                mat_A[22][2] * mat_B[208][0] +
                mat_A[22][3] * mat_B[216][0] +
                mat_A[23][0] * mat_B[224][0] +
                mat_A[23][1] * mat_B[232][0] +
                mat_A[23][2] * mat_B[240][0] +
                mat_A[23][3] * mat_B[248][0];
    mat_C[16][1] <=
                mat_A[16][0] * mat_B[0][1] +
                mat_A[16][1] * mat_B[8][1] +
                mat_A[16][2] * mat_B[16][1] +
                mat_A[16][3] * mat_B[24][1] +
                mat_A[17][0] * mat_B[32][1] +
                mat_A[17][1] * mat_B[40][1] +
                mat_A[17][2] * mat_B[48][1] +
                mat_A[17][3] * mat_B[56][1] +
                mat_A[18][0] * mat_B[64][1] +
                mat_A[18][1] * mat_B[72][1] +
                mat_A[18][2] * mat_B[80][1] +
                mat_A[18][3] * mat_B[88][1] +
                mat_A[19][0] * mat_B[96][1] +
                mat_A[19][1] * mat_B[104][1] +
                mat_A[19][2] * mat_B[112][1] +
                mat_A[19][3] * mat_B[120][1] +
                mat_A[20][0] * mat_B[128][1] +
                mat_A[20][1] * mat_B[136][1] +
                mat_A[20][2] * mat_B[144][1] +
                mat_A[20][3] * mat_B[152][1] +
                mat_A[21][0] * mat_B[160][1] +
                mat_A[21][1] * mat_B[168][1] +
                mat_A[21][2] * mat_B[176][1] +
                mat_A[21][3] * mat_B[184][1] +
                mat_A[22][0] * mat_B[192][1] +
                mat_A[22][1] * mat_B[200][1] +
                mat_A[22][2] * mat_B[208][1] +
                mat_A[22][3] * mat_B[216][1] +
                mat_A[23][0] * mat_B[224][1] +
                mat_A[23][1] * mat_B[232][1] +
                mat_A[23][2] * mat_B[240][1] +
                mat_A[23][3] * mat_B[248][1];
    mat_C[16][2] <=
                mat_A[16][0] * mat_B[0][2] +
                mat_A[16][1] * mat_B[8][2] +
                mat_A[16][2] * mat_B[16][2] +
                mat_A[16][3] * mat_B[24][2] +
                mat_A[17][0] * mat_B[32][2] +
                mat_A[17][1] * mat_B[40][2] +
                mat_A[17][2] * mat_B[48][2] +
                mat_A[17][3] * mat_B[56][2] +
                mat_A[18][0] * mat_B[64][2] +
                mat_A[18][1] * mat_B[72][2] +
                mat_A[18][2] * mat_B[80][2] +
                mat_A[18][3] * mat_B[88][2] +
                mat_A[19][0] * mat_B[96][2] +
                mat_A[19][1] * mat_B[104][2] +
                mat_A[19][2] * mat_B[112][2] +
                mat_A[19][3] * mat_B[120][2] +
                mat_A[20][0] * mat_B[128][2] +
                mat_A[20][1] * mat_B[136][2] +
                mat_A[20][2] * mat_B[144][2] +
                mat_A[20][3] * mat_B[152][2] +
                mat_A[21][0] * mat_B[160][2] +
                mat_A[21][1] * mat_B[168][2] +
                mat_A[21][2] * mat_B[176][2] +
                mat_A[21][3] * mat_B[184][2] +
                mat_A[22][0] * mat_B[192][2] +
                mat_A[22][1] * mat_B[200][2] +
                mat_A[22][2] * mat_B[208][2] +
                mat_A[22][3] * mat_B[216][2] +
                mat_A[23][0] * mat_B[224][2] +
                mat_A[23][1] * mat_B[232][2] +
                mat_A[23][2] * mat_B[240][2] +
                mat_A[23][3] * mat_B[248][2];
    mat_C[16][3] <=
                mat_A[16][0] * mat_B[0][3] +
                mat_A[16][1] * mat_B[8][3] +
                mat_A[16][2] * mat_B[16][3] +
                mat_A[16][3] * mat_B[24][3] +
                mat_A[17][0] * mat_B[32][3] +
                mat_A[17][1] * mat_B[40][3] +
                mat_A[17][2] * mat_B[48][3] +
                mat_A[17][3] * mat_B[56][3] +
                mat_A[18][0] * mat_B[64][3] +
                mat_A[18][1] * mat_B[72][3] +
                mat_A[18][2] * mat_B[80][3] +
                mat_A[18][3] * mat_B[88][3] +
                mat_A[19][0] * mat_B[96][3] +
                mat_A[19][1] * mat_B[104][3] +
                mat_A[19][2] * mat_B[112][3] +
                mat_A[19][3] * mat_B[120][3] +
                mat_A[20][0] * mat_B[128][3] +
                mat_A[20][1] * mat_B[136][3] +
                mat_A[20][2] * mat_B[144][3] +
                mat_A[20][3] * mat_B[152][3] +
                mat_A[21][0] * mat_B[160][3] +
                mat_A[21][1] * mat_B[168][3] +
                mat_A[21][2] * mat_B[176][3] +
                mat_A[21][3] * mat_B[184][3] +
                mat_A[22][0] * mat_B[192][3] +
                mat_A[22][1] * mat_B[200][3] +
                mat_A[22][2] * mat_B[208][3] +
                mat_A[22][3] * mat_B[216][3] +
                mat_A[23][0] * mat_B[224][3] +
                mat_A[23][1] * mat_B[232][3] +
                mat_A[23][2] * mat_B[240][3] +
                mat_A[23][3] * mat_B[248][3];
    mat_C[17][0] <=
                mat_A[16][0] * mat_B[1][0] +
                mat_A[16][1] * mat_B[9][0] +
                mat_A[16][2] * mat_B[17][0] +
                mat_A[16][3] * mat_B[25][0] +
                mat_A[17][0] * mat_B[33][0] +
                mat_A[17][1] * mat_B[41][0] +
                mat_A[17][2] * mat_B[49][0] +
                mat_A[17][3] * mat_B[57][0] +
                mat_A[18][0] * mat_B[65][0] +
                mat_A[18][1] * mat_B[73][0] +
                mat_A[18][2] * mat_B[81][0] +
                mat_A[18][3] * mat_B[89][0] +
                mat_A[19][0] * mat_B[97][0] +
                mat_A[19][1] * mat_B[105][0] +
                mat_A[19][2] * mat_B[113][0] +
                mat_A[19][3] * mat_B[121][0] +
                mat_A[20][0] * mat_B[129][0] +
                mat_A[20][1] * mat_B[137][0] +
                mat_A[20][2] * mat_B[145][0] +
                mat_A[20][3] * mat_B[153][0] +
                mat_A[21][0] * mat_B[161][0] +
                mat_A[21][1] * mat_B[169][0] +
                mat_A[21][2] * mat_B[177][0] +
                mat_A[21][3] * mat_B[185][0] +
                mat_A[22][0] * mat_B[193][0] +
                mat_A[22][1] * mat_B[201][0] +
                mat_A[22][2] * mat_B[209][0] +
                mat_A[22][3] * mat_B[217][0] +
                mat_A[23][0] * mat_B[225][0] +
                mat_A[23][1] * mat_B[233][0] +
                mat_A[23][2] * mat_B[241][0] +
                mat_A[23][3] * mat_B[249][0];
    mat_C[17][1] <=
                mat_A[16][0] * mat_B[1][1] +
                mat_A[16][1] * mat_B[9][1] +
                mat_A[16][2] * mat_B[17][1] +
                mat_A[16][3] * mat_B[25][1] +
                mat_A[17][0] * mat_B[33][1] +
                mat_A[17][1] * mat_B[41][1] +
                mat_A[17][2] * mat_B[49][1] +
                mat_A[17][3] * mat_B[57][1] +
                mat_A[18][0] * mat_B[65][1] +
                mat_A[18][1] * mat_B[73][1] +
                mat_A[18][2] * mat_B[81][1] +
                mat_A[18][3] * mat_B[89][1] +
                mat_A[19][0] * mat_B[97][1] +
                mat_A[19][1] * mat_B[105][1] +
                mat_A[19][2] * mat_B[113][1] +
                mat_A[19][3] * mat_B[121][1] +
                mat_A[20][0] * mat_B[129][1] +
                mat_A[20][1] * mat_B[137][1] +
                mat_A[20][2] * mat_B[145][1] +
                mat_A[20][3] * mat_B[153][1] +
                mat_A[21][0] * mat_B[161][1] +
                mat_A[21][1] * mat_B[169][1] +
                mat_A[21][2] * mat_B[177][1] +
                mat_A[21][3] * mat_B[185][1] +
                mat_A[22][0] * mat_B[193][1] +
                mat_A[22][1] * mat_B[201][1] +
                mat_A[22][2] * mat_B[209][1] +
                mat_A[22][3] * mat_B[217][1] +
                mat_A[23][0] * mat_B[225][1] +
                mat_A[23][1] * mat_B[233][1] +
                mat_A[23][2] * mat_B[241][1] +
                mat_A[23][3] * mat_B[249][1];
    mat_C[17][2] <=
                mat_A[16][0] * mat_B[1][2] +
                mat_A[16][1] * mat_B[9][2] +
                mat_A[16][2] * mat_B[17][2] +
                mat_A[16][3] * mat_B[25][2] +
                mat_A[17][0] * mat_B[33][2] +
                mat_A[17][1] * mat_B[41][2] +
                mat_A[17][2] * mat_B[49][2] +
                mat_A[17][3] * mat_B[57][2] +
                mat_A[18][0] * mat_B[65][2] +
                mat_A[18][1] * mat_B[73][2] +
                mat_A[18][2] * mat_B[81][2] +
                mat_A[18][3] * mat_B[89][2] +
                mat_A[19][0] * mat_B[97][2] +
                mat_A[19][1] * mat_B[105][2] +
                mat_A[19][2] * mat_B[113][2] +
                mat_A[19][3] * mat_B[121][2] +
                mat_A[20][0] * mat_B[129][2] +
                mat_A[20][1] * mat_B[137][2] +
                mat_A[20][2] * mat_B[145][2] +
                mat_A[20][3] * mat_B[153][2] +
                mat_A[21][0] * mat_B[161][2] +
                mat_A[21][1] * mat_B[169][2] +
                mat_A[21][2] * mat_B[177][2] +
                mat_A[21][3] * mat_B[185][2] +
                mat_A[22][0] * mat_B[193][2] +
                mat_A[22][1] * mat_B[201][2] +
                mat_A[22][2] * mat_B[209][2] +
                mat_A[22][3] * mat_B[217][2] +
                mat_A[23][0] * mat_B[225][2] +
                mat_A[23][1] * mat_B[233][2] +
                mat_A[23][2] * mat_B[241][2] +
                mat_A[23][3] * mat_B[249][2];
    mat_C[17][3] <=
                mat_A[16][0] * mat_B[1][3] +
                mat_A[16][1] * mat_B[9][3] +
                mat_A[16][2] * mat_B[17][3] +
                mat_A[16][3] * mat_B[25][3] +
                mat_A[17][0] * mat_B[33][3] +
                mat_A[17][1] * mat_B[41][3] +
                mat_A[17][2] * mat_B[49][3] +
                mat_A[17][3] * mat_B[57][3] +
                mat_A[18][0] * mat_B[65][3] +
                mat_A[18][1] * mat_B[73][3] +
                mat_A[18][2] * mat_B[81][3] +
                mat_A[18][3] * mat_B[89][3] +
                mat_A[19][0] * mat_B[97][3] +
                mat_A[19][1] * mat_B[105][3] +
                mat_A[19][2] * mat_B[113][3] +
                mat_A[19][3] * mat_B[121][3] +
                mat_A[20][0] * mat_B[129][3] +
                mat_A[20][1] * mat_B[137][3] +
                mat_A[20][2] * mat_B[145][3] +
                mat_A[20][3] * mat_B[153][3] +
                mat_A[21][0] * mat_B[161][3] +
                mat_A[21][1] * mat_B[169][3] +
                mat_A[21][2] * mat_B[177][3] +
                mat_A[21][3] * mat_B[185][3] +
                mat_A[22][0] * mat_B[193][3] +
                mat_A[22][1] * mat_B[201][3] +
                mat_A[22][2] * mat_B[209][3] +
                mat_A[22][3] * mat_B[217][3] +
                mat_A[23][0] * mat_B[225][3] +
                mat_A[23][1] * mat_B[233][3] +
                mat_A[23][2] * mat_B[241][3] +
                mat_A[23][3] * mat_B[249][3];
    mat_C[18][0] <=
                mat_A[16][0] * mat_B[2][0] +
                mat_A[16][1] * mat_B[10][0] +
                mat_A[16][2] * mat_B[18][0] +
                mat_A[16][3] * mat_B[26][0] +
                mat_A[17][0] * mat_B[34][0] +
                mat_A[17][1] * mat_B[42][0] +
                mat_A[17][2] * mat_B[50][0] +
                mat_A[17][3] * mat_B[58][0] +
                mat_A[18][0] * mat_B[66][0] +
                mat_A[18][1] * mat_B[74][0] +
                mat_A[18][2] * mat_B[82][0] +
                mat_A[18][3] * mat_B[90][0] +
                mat_A[19][0] * mat_B[98][0] +
                mat_A[19][1] * mat_B[106][0] +
                mat_A[19][2] * mat_B[114][0] +
                mat_A[19][3] * mat_B[122][0] +
                mat_A[20][0] * mat_B[130][0] +
                mat_A[20][1] * mat_B[138][0] +
                mat_A[20][2] * mat_B[146][0] +
                mat_A[20][3] * mat_B[154][0] +
                mat_A[21][0] * mat_B[162][0] +
                mat_A[21][1] * mat_B[170][0] +
                mat_A[21][2] * mat_B[178][0] +
                mat_A[21][3] * mat_B[186][0] +
                mat_A[22][0] * mat_B[194][0] +
                mat_A[22][1] * mat_B[202][0] +
                mat_A[22][2] * mat_B[210][0] +
                mat_A[22][3] * mat_B[218][0] +
                mat_A[23][0] * mat_B[226][0] +
                mat_A[23][1] * mat_B[234][0] +
                mat_A[23][2] * mat_B[242][0] +
                mat_A[23][3] * mat_B[250][0];
    mat_C[18][1] <=
                mat_A[16][0] * mat_B[2][1] +
                mat_A[16][1] * mat_B[10][1] +
                mat_A[16][2] * mat_B[18][1] +
                mat_A[16][3] * mat_B[26][1] +
                mat_A[17][0] * mat_B[34][1] +
                mat_A[17][1] * mat_B[42][1] +
                mat_A[17][2] * mat_B[50][1] +
                mat_A[17][3] * mat_B[58][1] +
                mat_A[18][0] * mat_B[66][1] +
                mat_A[18][1] * mat_B[74][1] +
                mat_A[18][2] * mat_B[82][1] +
                mat_A[18][3] * mat_B[90][1] +
                mat_A[19][0] * mat_B[98][1] +
                mat_A[19][1] * mat_B[106][1] +
                mat_A[19][2] * mat_B[114][1] +
                mat_A[19][3] * mat_B[122][1] +
                mat_A[20][0] * mat_B[130][1] +
                mat_A[20][1] * mat_B[138][1] +
                mat_A[20][2] * mat_B[146][1] +
                mat_A[20][3] * mat_B[154][1] +
                mat_A[21][0] * mat_B[162][1] +
                mat_A[21][1] * mat_B[170][1] +
                mat_A[21][2] * mat_B[178][1] +
                mat_A[21][3] * mat_B[186][1] +
                mat_A[22][0] * mat_B[194][1] +
                mat_A[22][1] * mat_B[202][1] +
                mat_A[22][2] * mat_B[210][1] +
                mat_A[22][3] * mat_B[218][1] +
                mat_A[23][0] * mat_B[226][1] +
                mat_A[23][1] * mat_B[234][1] +
                mat_A[23][2] * mat_B[242][1] +
                mat_A[23][3] * mat_B[250][1];
    mat_C[18][2] <=
                mat_A[16][0] * mat_B[2][2] +
                mat_A[16][1] * mat_B[10][2] +
                mat_A[16][2] * mat_B[18][2] +
                mat_A[16][3] * mat_B[26][2] +
                mat_A[17][0] * mat_B[34][2] +
                mat_A[17][1] * mat_B[42][2] +
                mat_A[17][2] * mat_B[50][2] +
                mat_A[17][3] * mat_B[58][2] +
                mat_A[18][0] * mat_B[66][2] +
                mat_A[18][1] * mat_B[74][2] +
                mat_A[18][2] * mat_B[82][2] +
                mat_A[18][3] * mat_B[90][2] +
                mat_A[19][0] * mat_B[98][2] +
                mat_A[19][1] * mat_B[106][2] +
                mat_A[19][2] * mat_B[114][2] +
                mat_A[19][3] * mat_B[122][2] +
                mat_A[20][0] * mat_B[130][2] +
                mat_A[20][1] * mat_B[138][2] +
                mat_A[20][2] * mat_B[146][2] +
                mat_A[20][3] * mat_B[154][2] +
                mat_A[21][0] * mat_B[162][2] +
                mat_A[21][1] * mat_B[170][2] +
                mat_A[21][2] * mat_B[178][2] +
                mat_A[21][3] * mat_B[186][2] +
                mat_A[22][0] * mat_B[194][2] +
                mat_A[22][1] * mat_B[202][2] +
                mat_A[22][2] * mat_B[210][2] +
                mat_A[22][3] * mat_B[218][2] +
                mat_A[23][0] * mat_B[226][2] +
                mat_A[23][1] * mat_B[234][2] +
                mat_A[23][2] * mat_B[242][2] +
                mat_A[23][3] * mat_B[250][2];
    mat_C[18][3] <=
                mat_A[16][0] * mat_B[2][3] +
                mat_A[16][1] * mat_B[10][3] +
                mat_A[16][2] * mat_B[18][3] +
                mat_A[16][3] * mat_B[26][3] +
                mat_A[17][0] * mat_B[34][3] +
                mat_A[17][1] * mat_B[42][3] +
                mat_A[17][2] * mat_B[50][3] +
                mat_A[17][3] * mat_B[58][3] +
                mat_A[18][0] * mat_B[66][3] +
                mat_A[18][1] * mat_B[74][3] +
                mat_A[18][2] * mat_B[82][3] +
                mat_A[18][3] * mat_B[90][3] +
                mat_A[19][0] * mat_B[98][3] +
                mat_A[19][1] * mat_B[106][3] +
                mat_A[19][2] * mat_B[114][3] +
                mat_A[19][3] * mat_B[122][3] +
                mat_A[20][0] * mat_B[130][3] +
                mat_A[20][1] * mat_B[138][3] +
                mat_A[20][2] * mat_B[146][3] +
                mat_A[20][3] * mat_B[154][3] +
                mat_A[21][0] * mat_B[162][3] +
                mat_A[21][1] * mat_B[170][3] +
                mat_A[21][2] * mat_B[178][3] +
                mat_A[21][3] * mat_B[186][3] +
                mat_A[22][0] * mat_B[194][3] +
                mat_A[22][1] * mat_B[202][3] +
                mat_A[22][2] * mat_B[210][3] +
                mat_A[22][3] * mat_B[218][3] +
                mat_A[23][0] * mat_B[226][3] +
                mat_A[23][1] * mat_B[234][3] +
                mat_A[23][2] * mat_B[242][3] +
                mat_A[23][3] * mat_B[250][3];
    mat_C[19][0] <=
                mat_A[16][0] * mat_B[3][0] +
                mat_A[16][1] * mat_B[11][0] +
                mat_A[16][2] * mat_B[19][0] +
                mat_A[16][3] * mat_B[27][0] +
                mat_A[17][0] * mat_B[35][0] +
                mat_A[17][1] * mat_B[43][0] +
                mat_A[17][2] * mat_B[51][0] +
                mat_A[17][3] * mat_B[59][0] +
                mat_A[18][0] * mat_B[67][0] +
                mat_A[18][1] * mat_B[75][0] +
                mat_A[18][2] * mat_B[83][0] +
                mat_A[18][3] * mat_B[91][0] +
                mat_A[19][0] * mat_B[99][0] +
                mat_A[19][1] * mat_B[107][0] +
                mat_A[19][2] * mat_B[115][0] +
                mat_A[19][3] * mat_B[123][0] +
                mat_A[20][0] * mat_B[131][0] +
                mat_A[20][1] * mat_B[139][0] +
                mat_A[20][2] * mat_B[147][0] +
                mat_A[20][3] * mat_B[155][0] +
                mat_A[21][0] * mat_B[163][0] +
                mat_A[21][1] * mat_B[171][0] +
                mat_A[21][2] * mat_B[179][0] +
                mat_A[21][3] * mat_B[187][0] +
                mat_A[22][0] * mat_B[195][0] +
                mat_A[22][1] * mat_B[203][0] +
                mat_A[22][2] * mat_B[211][0] +
                mat_A[22][3] * mat_B[219][0] +
                mat_A[23][0] * mat_B[227][0] +
                mat_A[23][1] * mat_B[235][0] +
                mat_A[23][2] * mat_B[243][0] +
                mat_A[23][3] * mat_B[251][0];
    mat_C[19][1] <=
                mat_A[16][0] * mat_B[3][1] +
                mat_A[16][1] * mat_B[11][1] +
                mat_A[16][2] * mat_B[19][1] +
                mat_A[16][3] * mat_B[27][1] +
                mat_A[17][0] * mat_B[35][1] +
                mat_A[17][1] * mat_B[43][1] +
                mat_A[17][2] * mat_B[51][1] +
                mat_A[17][3] * mat_B[59][1] +
                mat_A[18][0] * mat_B[67][1] +
                mat_A[18][1] * mat_B[75][1] +
                mat_A[18][2] * mat_B[83][1] +
                mat_A[18][3] * mat_B[91][1] +
                mat_A[19][0] * mat_B[99][1] +
                mat_A[19][1] * mat_B[107][1] +
                mat_A[19][2] * mat_B[115][1] +
                mat_A[19][3] * mat_B[123][1] +
                mat_A[20][0] * mat_B[131][1] +
                mat_A[20][1] * mat_B[139][1] +
                mat_A[20][2] * mat_B[147][1] +
                mat_A[20][3] * mat_B[155][1] +
                mat_A[21][0] * mat_B[163][1] +
                mat_A[21][1] * mat_B[171][1] +
                mat_A[21][2] * mat_B[179][1] +
                mat_A[21][3] * mat_B[187][1] +
                mat_A[22][0] * mat_B[195][1] +
                mat_A[22][1] * mat_B[203][1] +
                mat_A[22][2] * mat_B[211][1] +
                mat_A[22][3] * mat_B[219][1] +
                mat_A[23][0] * mat_B[227][1] +
                mat_A[23][1] * mat_B[235][1] +
                mat_A[23][2] * mat_B[243][1] +
                mat_A[23][3] * mat_B[251][1];
    mat_C[19][2] <=
                mat_A[16][0] * mat_B[3][2] +
                mat_A[16][1] * mat_B[11][2] +
                mat_A[16][2] * mat_B[19][2] +
                mat_A[16][3] * mat_B[27][2] +
                mat_A[17][0] * mat_B[35][2] +
                mat_A[17][1] * mat_B[43][2] +
                mat_A[17][2] * mat_B[51][2] +
                mat_A[17][3] * mat_B[59][2] +
                mat_A[18][0] * mat_B[67][2] +
                mat_A[18][1] * mat_B[75][2] +
                mat_A[18][2] * mat_B[83][2] +
                mat_A[18][3] * mat_B[91][2] +
                mat_A[19][0] * mat_B[99][2] +
                mat_A[19][1] * mat_B[107][2] +
                mat_A[19][2] * mat_B[115][2] +
                mat_A[19][3] * mat_B[123][2] +
                mat_A[20][0] * mat_B[131][2] +
                mat_A[20][1] * mat_B[139][2] +
                mat_A[20][2] * mat_B[147][2] +
                mat_A[20][3] * mat_B[155][2] +
                mat_A[21][0] * mat_B[163][2] +
                mat_A[21][1] * mat_B[171][2] +
                mat_A[21][2] * mat_B[179][2] +
                mat_A[21][3] * mat_B[187][2] +
                mat_A[22][0] * mat_B[195][2] +
                mat_A[22][1] * mat_B[203][2] +
                mat_A[22][2] * mat_B[211][2] +
                mat_A[22][3] * mat_B[219][2] +
                mat_A[23][0] * mat_B[227][2] +
                mat_A[23][1] * mat_B[235][2] +
                mat_A[23][2] * mat_B[243][2] +
                mat_A[23][3] * mat_B[251][2];
    mat_C[19][3] <=
                mat_A[16][0] * mat_B[3][3] +
                mat_A[16][1] * mat_B[11][3] +
                mat_A[16][2] * mat_B[19][3] +
                mat_A[16][3] * mat_B[27][3] +
                mat_A[17][0] * mat_B[35][3] +
                mat_A[17][1] * mat_B[43][3] +
                mat_A[17][2] * mat_B[51][3] +
                mat_A[17][3] * mat_B[59][3] +
                mat_A[18][0] * mat_B[67][3] +
                mat_A[18][1] * mat_B[75][3] +
                mat_A[18][2] * mat_B[83][3] +
                mat_A[18][3] * mat_B[91][3] +
                mat_A[19][0] * mat_B[99][3] +
                mat_A[19][1] * mat_B[107][3] +
                mat_A[19][2] * mat_B[115][3] +
                mat_A[19][3] * mat_B[123][3] +
                mat_A[20][0] * mat_B[131][3] +
                mat_A[20][1] * mat_B[139][3] +
                mat_A[20][2] * mat_B[147][3] +
                mat_A[20][3] * mat_B[155][3] +
                mat_A[21][0] * mat_B[163][3] +
                mat_A[21][1] * mat_B[171][3] +
                mat_A[21][2] * mat_B[179][3] +
                mat_A[21][3] * mat_B[187][3] +
                mat_A[22][0] * mat_B[195][3] +
                mat_A[22][1] * mat_B[203][3] +
                mat_A[22][2] * mat_B[211][3] +
                mat_A[22][3] * mat_B[219][3] +
                mat_A[23][0] * mat_B[227][3] +
                mat_A[23][1] * mat_B[235][3] +
                mat_A[23][2] * mat_B[243][3] +
                mat_A[23][3] * mat_B[251][3];
    mat_C[20][0] <=
                mat_A[16][0] * mat_B[4][0] +
                mat_A[16][1] * mat_B[12][0] +
                mat_A[16][2] * mat_B[20][0] +
                mat_A[16][3] * mat_B[28][0] +
                mat_A[17][0] * mat_B[36][0] +
                mat_A[17][1] * mat_B[44][0] +
                mat_A[17][2] * mat_B[52][0] +
                mat_A[17][3] * mat_B[60][0] +
                mat_A[18][0] * mat_B[68][0] +
                mat_A[18][1] * mat_B[76][0] +
                mat_A[18][2] * mat_B[84][0] +
                mat_A[18][3] * mat_B[92][0] +
                mat_A[19][0] * mat_B[100][0] +
                mat_A[19][1] * mat_B[108][0] +
                mat_A[19][2] * mat_B[116][0] +
                mat_A[19][3] * mat_B[124][0] +
                mat_A[20][0] * mat_B[132][0] +
                mat_A[20][1] * mat_B[140][0] +
                mat_A[20][2] * mat_B[148][0] +
                mat_A[20][3] * mat_B[156][0] +
                mat_A[21][0] * mat_B[164][0] +
                mat_A[21][1] * mat_B[172][0] +
                mat_A[21][2] * mat_B[180][0] +
                mat_A[21][3] * mat_B[188][0] +
                mat_A[22][0] * mat_B[196][0] +
                mat_A[22][1] * mat_B[204][0] +
                mat_A[22][2] * mat_B[212][0] +
                mat_A[22][3] * mat_B[220][0] +
                mat_A[23][0] * mat_B[228][0] +
                mat_A[23][1] * mat_B[236][0] +
                mat_A[23][2] * mat_B[244][0] +
                mat_A[23][3] * mat_B[252][0];
    mat_C[20][1] <=
                mat_A[16][0] * mat_B[4][1] +
                mat_A[16][1] * mat_B[12][1] +
                mat_A[16][2] * mat_B[20][1] +
                mat_A[16][3] * mat_B[28][1] +
                mat_A[17][0] * mat_B[36][1] +
                mat_A[17][1] * mat_B[44][1] +
                mat_A[17][2] * mat_B[52][1] +
                mat_A[17][3] * mat_B[60][1] +
                mat_A[18][0] * mat_B[68][1] +
                mat_A[18][1] * mat_B[76][1] +
                mat_A[18][2] * mat_B[84][1] +
                mat_A[18][3] * mat_B[92][1] +
                mat_A[19][0] * mat_B[100][1] +
                mat_A[19][1] * mat_B[108][1] +
                mat_A[19][2] * mat_B[116][1] +
                mat_A[19][3] * mat_B[124][1] +
                mat_A[20][0] * mat_B[132][1] +
                mat_A[20][1] * mat_B[140][1] +
                mat_A[20][2] * mat_B[148][1] +
                mat_A[20][3] * mat_B[156][1] +
                mat_A[21][0] * mat_B[164][1] +
                mat_A[21][1] * mat_B[172][1] +
                mat_A[21][2] * mat_B[180][1] +
                mat_A[21][3] * mat_B[188][1] +
                mat_A[22][0] * mat_B[196][1] +
                mat_A[22][1] * mat_B[204][1] +
                mat_A[22][2] * mat_B[212][1] +
                mat_A[22][3] * mat_B[220][1] +
                mat_A[23][0] * mat_B[228][1] +
                mat_A[23][1] * mat_B[236][1] +
                mat_A[23][2] * mat_B[244][1] +
                mat_A[23][3] * mat_B[252][1];
    mat_C[20][2] <=
                mat_A[16][0] * mat_B[4][2] +
                mat_A[16][1] * mat_B[12][2] +
                mat_A[16][2] * mat_B[20][2] +
                mat_A[16][3] * mat_B[28][2] +
                mat_A[17][0] * mat_B[36][2] +
                mat_A[17][1] * mat_B[44][2] +
                mat_A[17][2] * mat_B[52][2] +
                mat_A[17][3] * mat_B[60][2] +
                mat_A[18][0] * mat_B[68][2] +
                mat_A[18][1] * mat_B[76][2] +
                mat_A[18][2] * mat_B[84][2] +
                mat_A[18][3] * mat_B[92][2] +
                mat_A[19][0] * mat_B[100][2] +
                mat_A[19][1] * mat_B[108][2] +
                mat_A[19][2] * mat_B[116][2] +
                mat_A[19][3] * mat_B[124][2] +
                mat_A[20][0] * mat_B[132][2] +
                mat_A[20][1] * mat_B[140][2] +
                mat_A[20][2] * mat_B[148][2] +
                mat_A[20][3] * mat_B[156][2] +
                mat_A[21][0] * mat_B[164][2] +
                mat_A[21][1] * mat_B[172][2] +
                mat_A[21][2] * mat_B[180][2] +
                mat_A[21][3] * mat_B[188][2] +
                mat_A[22][0] * mat_B[196][2] +
                mat_A[22][1] * mat_B[204][2] +
                mat_A[22][2] * mat_B[212][2] +
                mat_A[22][3] * mat_B[220][2] +
                mat_A[23][0] * mat_B[228][2] +
                mat_A[23][1] * mat_B[236][2] +
                mat_A[23][2] * mat_B[244][2] +
                mat_A[23][3] * mat_B[252][2];
    mat_C[20][3] <=
                mat_A[16][0] * mat_B[4][3] +
                mat_A[16][1] * mat_B[12][3] +
                mat_A[16][2] * mat_B[20][3] +
                mat_A[16][3] * mat_B[28][3] +
                mat_A[17][0] * mat_B[36][3] +
                mat_A[17][1] * mat_B[44][3] +
                mat_A[17][2] * mat_B[52][3] +
                mat_A[17][3] * mat_B[60][3] +
                mat_A[18][0] * mat_B[68][3] +
                mat_A[18][1] * mat_B[76][3] +
                mat_A[18][2] * mat_B[84][3] +
                mat_A[18][3] * mat_B[92][3] +
                mat_A[19][0] * mat_B[100][3] +
                mat_A[19][1] * mat_B[108][3] +
                mat_A[19][2] * mat_B[116][3] +
                mat_A[19][3] * mat_B[124][3] +
                mat_A[20][0] * mat_B[132][3] +
                mat_A[20][1] * mat_B[140][3] +
                mat_A[20][2] * mat_B[148][3] +
                mat_A[20][3] * mat_B[156][3] +
                mat_A[21][0] * mat_B[164][3] +
                mat_A[21][1] * mat_B[172][3] +
                mat_A[21][2] * mat_B[180][3] +
                mat_A[21][3] * mat_B[188][3] +
                mat_A[22][0] * mat_B[196][3] +
                mat_A[22][1] * mat_B[204][3] +
                mat_A[22][2] * mat_B[212][3] +
                mat_A[22][3] * mat_B[220][3] +
                mat_A[23][0] * mat_B[228][3] +
                mat_A[23][1] * mat_B[236][3] +
                mat_A[23][2] * mat_B[244][3] +
                mat_A[23][3] * mat_B[252][3];
    mat_C[21][0] <=
                mat_A[16][0] * mat_B[5][0] +
                mat_A[16][1] * mat_B[13][0] +
                mat_A[16][2] * mat_B[21][0] +
                mat_A[16][3] * mat_B[29][0] +
                mat_A[17][0] * mat_B[37][0] +
                mat_A[17][1] * mat_B[45][0] +
                mat_A[17][2] * mat_B[53][0] +
                mat_A[17][3] * mat_B[61][0] +
                mat_A[18][0] * mat_B[69][0] +
                mat_A[18][1] * mat_B[77][0] +
                mat_A[18][2] * mat_B[85][0] +
                mat_A[18][3] * mat_B[93][0] +
                mat_A[19][0] * mat_B[101][0] +
                mat_A[19][1] * mat_B[109][0] +
                mat_A[19][2] * mat_B[117][0] +
                mat_A[19][3] * mat_B[125][0] +
                mat_A[20][0] * mat_B[133][0] +
                mat_A[20][1] * mat_B[141][0] +
                mat_A[20][2] * mat_B[149][0] +
                mat_A[20][3] * mat_B[157][0] +
                mat_A[21][0] * mat_B[165][0] +
                mat_A[21][1] * mat_B[173][0] +
                mat_A[21][2] * mat_B[181][0] +
                mat_A[21][3] * mat_B[189][0] +
                mat_A[22][0] * mat_B[197][0] +
                mat_A[22][1] * mat_B[205][0] +
                mat_A[22][2] * mat_B[213][0] +
                mat_A[22][3] * mat_B[221][0] +
                mat_A[23][0] * mat_B[229][0] +
                mat_A[23][1] * mat_B[237][0] +
                mat_A[23][2] * mat_B[245][0] +
                mat_A[23][3] * mat_B[253][0];
    mat_C[21][1] <=
                mat_A[16][0] * mat_B[5][1] +
                mat_A[16][1] * mat_B[13][1] +
                mat_A[16][2] * mat_B[21][1] +
                mat_A[16][3] * mat_B[29][1] +
                mat_A[17][0] * mat_B[37][1] +
                mat_A[17][1] * mat_B[45][1] +
                mat_A[17][2] * mat_B[53][1] +
                mat_A[17][3] * mat_B[61][1] +
                mat_A[18][0] * mat_B[69][1] +
                mat_A[18][1] * mat_B[77][1] +
                mat_A[18][2] * mat_B[85][1] +
                mat_A[18][3] * mat_B[93][1] +
                mat_A[19][0] * mat_B[101][1] +
                mat_A[19][1] * mat_B[109][1] +
                mat_A[19][2] * mat_B[117][1] +
                mat_A[19][3] * mat_B[125][1] +
                mat_A[20][0] * mat_B[133][1] +
                mat_A[20][1] * mat_B[141][1] +
                mat_A[20][2] * mat_B[149][1] +
                mat_A[20][3] * mat_B[157][1] +
                mat_A[21][0] * mat_B[165][1] +
                mat_A[21][1] * mat_B[173][1] +
                mat_A[21][2] * mat_B[181][1] +
                mat_A[21][3] * mat_B[189][1] +
                mat_A[22][0] * mat_B[197][1] +
                mat_A[22][1] * mat_B[205][1] +
                mat_A[22][2] * mat_B[213][1] +
                mat_A[22][3] * mat_B[221][1] +
                mat_A[23][0] * mat_B[229][1] +
                mat_A[23][1] * mat_B[237][1] +
                mat_A[23][2] * mat_B[245][1] +
                mat_A[23][3] * mat_B[253][1];
    mat_C[21][2] <=
                mat_A[16][0] * mat_B[5][2] +
                mat_A[16][1] * mat_B[13][2] +
                mat_A[16][2] * mat_B[21][2] +
                mat_A[16][3] * mat_B[29][2] +
                mat_A[17][0] * mat_B[37][2] +
                mat_A[17][1] * mat_B[45][2] +
                mat_A[17][2] * mat_B[53][2] +
                mat_A[17][3] * mat_B[61][2] +
                mat_A[18][0] * mat_B[69][2] +
                mat_A[18][1] * mat_B[77][2] +
                mat_A[18][2] * mat_B[85][2] +
                mat_A[18][3] * mat_B[93][2] +
                mat_A[19][0] * mat_B[101][2] +
                mat_A[19][1] * mat_B[109][2] +
                mat_A[19][2] * mat_B[117][2] +
                mat_A[19][3] * mat_B[125][2] +
                mat_A[20][0] * mat_B[133][2] +
                mat_A[20][1] * mat_B[141][2] +
                mat_A[20][2] * mat_B[149][2] +
                mat_A[20][3] * mat_B[157][2] +
                mat_A[21][0] * mat_B[165][2] +
                mat_A[21][1] * mat_B[173][2] +
                mat_A[21][2] * mat_B[181][2] +
                mat_A[21][3] * mat_B[189][2] +
                mat_A[22][0] * mat_B[197][2] +
                mat_A[22][1] * mat_B[205][2] +
                mat_A[22][2] * mat_B[213][2] +
                mat_A[22][3] * mat_B[221][2] +
                mat_A[23][0] * mat_B[229][2] +
                mat_A[23][1] * mat_B[237][2] +
                mat_A[23][2] * mat_B[245][2] +
                mat_A[23][3] * mat_B[253][2];
    mat_C[21][3] <=
                mat_A[16][0] * mat_B[5][3] +
                mat_A[16][1] * mat_B[13][3] +
                mat_A[16][2] * mat_B[21][3] +
                mat_A[16][3] * mat_B[29][3] +
                mat_A[17][0] * mat_B[37][3] +
                mat_A[17][1] * mat_B[45][3] +
                mat_A[17][2] * mat_B[53][3] +
                mat_A[17][3] * mat_B[61][3] +
                mat_A[18][0] * mat_B[69][3] +
                mat_A[18][1] * mat_B[77][3] +
                mat_A[18][2] * mat_B[85][3] +
                mat_A[18][3] * mat_B[93][3] +
                mat_A[19][0] * mat_B[101][3] +
                mat_A[19][1] * mat_B[109][3] +
                mat_A[19][2] * mat_B[117][3] +
                mat_A[19][3] * mat_B[125][3] +
                mat_A[20][0] * mat_B[133][3] +
                mat_A[20][1] * mat_B[141][3] +
                mat_A[20][2] * mat_B[149][3] +
                mat_A[20][3] * mat_B[157][3] +
                mat_A[21][0] * mat_B[165][3] +
                mat_A[21][1] * mat_B[173][3] +
                mat_A[21][2] * mat_B[181][3] +
                mat_A[21][3] * mat_B[189][3] +
                mat_A[22][0] * mat_B[197][3] +
                mat_A[22][1] * mat_B[205][3] +
                mat_A[22][2] * mat_B[213][3] +
                mat_A[22][3] * mat_B[221][3] +
                mat_A[23][0] * mat_B[229][3] +
                mat_A[23][1] * mat_B[237][3] +
                mat_A[23][2] * mat_B[245][3] +
                mat_A[23][3] * mat_B[253][3];
    mat_C[22][0] <=
                mat_A[16][0] * mat_B[6][0] +
                mat_A[16][1] * mat_B[14][0] +
                mat_A[16][2] * mat_B[22][0] +
                mat_A[16][3] * mat_B[30][0] +
                mat_A[17][0] * mat_B[38][0] +
                mat_A[17][1] * mat_B[46][0] +
                mat_A[17][2] * mat_B[54][0] +
                mat_A[17][3] * mat_B[62][0] +
                mat_A[18][0] * mat_B[70][0] +
                mat_A[18][1] * mat_B[78][0] +
                mat_A[18][2] * mat_B[86][0] +
                mat_A[18][3] * mat_B[94][0] +
                mat_A[19][0] * mat_B[102][0] +
                mat_A[19][1] * mat_B[110][0] +
                mat_A[19][2] * mat_B[118][0] +
                mat_A[19][3] * mat_B[126][0] +
                mat_A[20][0] * mat_B[134][0] +
                mat_A[20][1] * mat_B[142][0] +
                mat_A[20][2] * mat_B[150][0] +
                mat_A[20][3] * mat_B[158][0] +
                mat_A[21][0] * mat_B[166][0] +
                mat_A[21][1] * mat_B[174][0] +
                mat_A[21][2] * mat_B[182][0] +
                mat_A[21][3] * mat_B[190][0] +
                mat_A[22][0] * mat_B[198][0] +
                mat_A[22][1] * mat_B[206][0] +
                mat_A[22][2] * mat_B[214][0] +
                mat_A[22][3] * mat_B[222][0] +
                mat_A[23][0] * mat_B[230][0] +
                mat_A[23][1] * mat_B[238][0] +
                mat_A[23][2] * mat_B[246][0] +
                mat_A[23][3] * mat_B[254][0];
    mat_C[22][1] <=
                mat_A[16][0] * mat_B[6][1] +
                mat_A[16][1] * mat_B[14][1] +
                mat_A[16][2] * mat_B[22][1] +
                mat_A[16][3] * mat_B[30][1] +
                mat_A[17][0] * mat_B[38][1] +
                mat_A[17][1] * mat_B[46][1] +
                mat_A[17][2] * mat_B[54][1] +
                mat_A[17][3] * mat_B[62][1] +
                mat_A[18][0] * mat_B[70][1] +
                mat_A[18][1] * mat_B[78][1] +
                mat_A[18][2] * mat_B[86][1] +
                mat_A[18][3] * mat_B[94][1] +
                mat_A[19][0] * mat_B[102][1] +
                mat_A[19][1] * mat_B[110][1] +
                mat_A[19][2] * mat_B[118][1] +
                mat_A[19][3] * mat_B[126][1] +
                mat_A[20][0] * mat_B[134][1] +
                mat_A[20][1] * mat_B[142][1] +
                mat_A[20][2] * mat_B[150][1] +
                mat_A[20][3] * mat_B[158][1] +
                mat_A[21][0] * mat_B[166][1] +
                mat_A[21][1] * mat_B[174][1] +
                mat_A[21][2] * mat_B[182][1] +
                mat_A[21][3] * mat_B[190][1] +
                mat_A[22][0] * mat_B[198][1] +
                mat_A[22][1] * mat_B[206][1] +
                mat_A[22][2] * mat_B[214][1] +
                mat_A[22][3] * mat_B[222][1] +
                mat_A[23][0] * mat_B[230][1] +
                mat_A[23][1] * mat_B[238][1] +
                mat_A[23][2] * mat_B[246][1] +
                mat_A[23][3] * mat_B[254][1];
    mat_C[22][2] <=
                mat_A[16][0] * mat_B[6][2] +
                mat_A[16][1] * mat_B[14][2] +
                mat_A[16][2] * mat_B[22][2] +
                mat_A[16][3] * mat_B[30][2] +
                mat_A[17][0] * mat_B[38][2] +
                mat_A[17][1] * mat_B[46][2] +
                mat_A[17][2] * mat_B[54][2] +
                mat_A[17][3] * mat_B[62][2] +
                mat_A[18][0] * mat_B[70][2] +
                mat_A[18][1] * mat_B[78][2] +
                mat_A[18][2] * mat_B[86][2] +
                mat_A[18][3] * mat_B[94][2] +
                mat_A[19][0] * mat_B[102][2] +
                mat_A[19][1] * mat_B[110][2] +
                mat_A[19][2] * mat_B[118][2] +
                mat_A[19][3] * mat_B[126][2] +
                mat_A[20][0] * mat_B[134][2] +
                mat_A[20][1] * mat_B[142][2] +
                mat_A[20][2] * mat_B[150][2] +
                mat_A[20][3] * mat_B[158][2] +
                mat_A[21][0] * mat_B[166][2] +
                mat_A[21][1] * mat_B[174][2] +
                mat_A[21][2] * mat_B[182][2] +
                mat_A[21][3] * mat_B[190][2] +
                mat_A[22][0] * mat_B[198][2] +
                mat_A[22][1] * mat_B[206][2] +
                mat_A[22][2] * mat_B[214][2] +
                mat_A[22][3] * mat_B[222][2] +
                mat_A[23][0] * mat_B[230][2] +
                mat_A[23][1] * mat_B[238][2] +
                mat_A[23][2] * mat_B[246][2] +
                mat_A[23][3] * mat_B[254][2];
    mat_C[22][3] <=
                mat_A[16][0] * mat_B[6][3] +
                mat_A[16][1] * mat_B[14][3] +
                mat_A[16][2] * mat_B[22][3] +
                mat_A[16][3] * mat_B[30][3] +
                mat_A[17][0] * mat_B[38][3] +
                mat_A[17][1] * mat_B[46][3] +
                mat_A[17][2] * mat_B[54][3] +
                mat_A[17][3] * mat_B[62][3] +
                mat_A[18][0] * mat_B[70][3] +
                mat_A[18][1] * mat_B[78][3] +
                mat_A[18][2] * mat_B[86][3] +
                mat_A[18][3] * mat_B[94][3] +
                mat_A[19][0] * mat_B[102][3] +
                mat_A[19][1] * mat_B[110][3] +
                mat_A[19][2] * mat_B[118][3] +
                mat_A[19][3] * mat_B[126][3] +
                mat_A[20][0] * mat_B[134][3] +
                mat_A[20][1] * mat_B[142][3] +
                mat_A[20][2] * mat_B[150][3] +
                mat_A[20][3] * mat_B[158][3] +
                mat_A[21][0] * mat_B[166][3] +
                mat_A[21][1] * mat_B[174][3] +
                mat_A[21][2] * mat_B[182][3] +
                mat_A[21][3] * mat_B[190][3] +
                mat_A[22][0] * mat_B[198][3] +
                mat_A[22][1] * mat_B[206][3] +
                mat_A[22][2] * mat_B[214][3] +
                mat_A[22][3] * mat_B[222][3] +
                mat_A[23][0] * mat_B[230][3] +
                mat_A[23][1] * mat_B[238][3] +
                mat_A[23][2] * mat_B[246][3] +
                mat_A[23][3] * mat_B[254][3];
    mat_C[23][0] <=
                mat_A[16][0] * mat_B[7][0] +
                mat_A[16][1] * mat_B[15][0] +
                mat_A[16][2] * mat_B[23][0] +
                mat_A[16][3] * mat_B[31][0] +
                mat_A[17][0] * mat_B[39][0] +
                mat_A[17][1] * mat_B[47][0] +
                mat_A[17][2] * mat_B[55][0] +
                mat_A[17][3] * mat_B[63][0] +
                mat_A[18][0] * mat_B[71][0] +
                mat_A[18][1] * mat_B[79][0] +
                mat_A[18][2] * mat_B[87][0] +
                mat_A[18][3] * mat_B[95][0] +
                mat_A[19][0] * mat_B[103][0] +
                mat_A[19][1] * mat_B[111][0] +
                mat_A[19][2] * mat_B[119][0] +
                mat_A[19][3] * mat_B[127][0] +
                mat_A[20][0] * mat_B[135][0] +
                mat_A[20][1] * mat_B[143][0] +
                mat_A[20][2] * mat_B[151][0] +
                mat_A[20][3] * mat_B[159][0] +
                mat_A[21][0] * mat_B[167][0] +
                mat_A[21][1] * mat_B[175][0] +
                mat_A[21][2] * mat_B[183][0] +
                mat_A[21][3] * mat_B[191][0] +
                mat_A[22][0] * mat_B[199][0] +
                mat_A[22][1] * mat_B[207][0] +
                mat_A[22][2] * mat_B[215][0] +
                mat_A[22][3] * mat_B[223][0] +
                mat_A[23][0] * mat_B[231][0] +
                mat_A[23][1] * mat_B[239][0] +
                mat_A[23][2] * mat_B[247][0] +
                mat_A[23][3] * mat_B[255][0];
    mat_C[23][1] <=
                mat_A[16][0] * mat_B[7][1] +
                mat_A[16][1] * mat_B[15][1] +
                mat_A[16][2] * mat_B[23][1] +
                mat_A[16][3] * mat_B[31][1] +
                mat_A[17][0] * mat_B[39][1] +
                mat_A[17][1] * mat_B[47][1] +
                mat_A[17][2] * mat_B[55][1] +
                mat_A[17][3] * mat_B[63][1] +
                mat_A[18][0] * mat_B[71][1] +
                mat_A[18][1] * mat_B[79][1] +
                mat_A[18][2] * mat_B[87][1] +
                mat_A[18][3] * mat_B[95][1] +
                mat_A[19][0] * mat_B[103][1] +
                mat_A[19][1] * mat_B[111][1] +
                mat_A[19][2] * mat_B[119][1] +
                mat_A[19][3] * mat_B[127][1] +
                mat_A[20][0] * mat_B[135][1] +
                mat_A[20][1] * mat_B[143][1] +
                mat_A[20][2] * mat_B[151][1] +
                mat_A[20][3] * mat_B[159][1] +
                mat_A[21][0] * mat_B[167][1] +
                mat_A[21][1] * mat_B[175][1] +
                mat_A[21][2] * mat_B[183][1] +
                mat_A[21][3] * mat_B[191][1] +
                mat_A[22][0] * mat_B[199][1] +
                mat_A[22][1] * mat_B[207][1] +
                mat_A[22][2] * mat_B[215][1] +
                mat_A[22][3] * mat_B[223][1] +
                mat_A[23][0] * mat_B[231][1] +
                mat_A[23][1] * mat_B[239][1] +
                mat_A[23][2] * mat_B[247][1] +
                mat_A[23][3] * mat_B[255][1];
    mat_C[23][2] <=
                mat_A[16][0] * mat_B[7][2] +
                mat_A[16][1] * mat_B[15][2] +
                mat_A[16][2] * mat_B[23][2] +
                mat_A[16][3] * mat_B[31][2] +
                mat_A[17][0] * mat_B[39][2] +
                mat_A[17][1] * mat_B[47][2] +
                mat_A[17][2] * mat_B[55][2] +
                mat_A[17][3] * mat_B[63][2] +
                mat_A[18][0] * mat_B[71][2] +
                mat_A[18][1] * mat_B[79][2] +
                mat_A[18][2] * mat_B[87][2] +
                mat_A[18][3] * mat_B[95][2] +
                mat_A[19][0] * mat_B[103][2] +
                mat_A[19][1] * mat_B[111][2] +
                mat_A[19][2] * mat_B[119][2] +
                mat_A[19][3] * mat_B[127][2] +
                mat_A[20][0] * mat_B[135][2] +
                mat_A[20][1] * mat_B[143][2] +
                mat_A[20][2] * mat_B[151][2] +
                mat_A[20][3] * mat_B[159][2] +
                mat_A[21][0] * mat_B[167][2] +
                mat_A[21][1] * mat_B[175][2] +
                mat_A[21][2] * mat_B[183][2] +
                mat_A[21][3] * mat_B[191][2] +
                mat_A[22][0] * mat_B[199][2] +
                mat_A[22][1] * mat_B[207][2] +
                mat_A[22][2] * mat_B[215][2] +
                mat_A[22][3] * mat_B[223][2] +
                mat_A[23][0] * mat_B[231][2] +
                mat_A[23][1] * mat_B[239][2] +
                mat_A[23][2] * mat_B[247][2] +
                mat_A[23][3] * mat_B[255][2];
    mat_C[23][3] <=
                mat_A[16][0] * mat_B[7][3] +
                mat_A[16][1] * mat_B[15][3] +
                mat_A[16][2] * mat_B[23][3] +
                mat_A[16][3] * mat_B[31][3] +
                mat_A[17][0] * mat_B[39][3] +
                mat_A[17][1] * mat_B[47][3] +
                mat_A[17][2] * mat_B[55][3] +
                mat_A[17][3] * mat_B[63][3] +
                mat_A[18][0] * mat_B[71][3] +
                mat_A[18][1] * mat_B[79][3] +
                mat_A[18][2] * mat_B[87][3] +
                mat_A[18][3] * mat_B[95][3] +
                mat_A[19][0] * mat_B[103][3] +
                mat_A[19][1] * mat_B[111][3] +
                mat_A[19][2] * mat_B[119][3] +
                mat_A[19][3] * mat_B[127][3] +
                mat_A[20][0] * mat_B[135][3] +
                mat_A[20][1] * mat_B[143][3] +
                mat_A[20][2] * mat_B[151][3] +
                mat_A[20][3] * mat_B[159][3] +
                mat_A[21][0] * mat_B[167][3] +
                mat_A[21][1] * mat_B[175][3] +
                mat_A[21][2] * mat_B[183][3] +
                mat_A[21][3] * mat_B[191][3] +
                mat_A[22][0] * mat_B[199][3] +
                mat_A[22][1] * mat_B[207][3] +
                mat_A[22][2] * mat_B[215][3] +
                mat_A[22][3] * mat_B[223][3] +
                mat_A[23][0] * mat_B[231][3] +
                mat_A[23][1] * mat_B[239][3] +
                mat_A[23][2] * mat_B[247][3] +
                mat_A[23][3] * mat_B[255][3];
    mat_C[24][0] <=
                mat_A[24][0] * mat_B[0][0] +
                mat_A[24][1] * mat_B[8][0] +
                mat_A[24][2] * mat_B[16][0] +
                mat_A[24][3] * mat_B[24][0] +
                mat_A[25][0] * mat_B[32][0] +
                mat_A[25][1] * mat_B[40][0] +
                mat_A[25][2] * mat_B[48][0] +
                mat_A[25][3] * mat_B[56][0] +
                mat_A[26][0] * mat_B[64][0] +
                mat_A[26][1] * mat_B[72][0] +
                mat_A[26][2] * mat_B[80][0] +
                mat_A[26][3] * mat_B[88][0] +
                mat_A[27][0] * mat_B[96][0] +
                mat_A[27][1] * mat_B[104][0] +
                mat_A[27][2] * mat_B[112][0] +
                mat_A[27][3] * mat_B[120][0] +
                mat_A[28][0] * mat_B[128][0] +
                mat_A[28][1] * mat_B[136][0] +
                mat_A[28][2] * mat_B[144][0] +
                mat_A[28][3] * mat_B[152][0] +
                mat_A[29][0] * mat_B[160][0] +
                mat_A[29][1] * mat_B[168][0] +
                mat_A[29][2] * mat_B[176][0] +
                mat_A[29][3] * mat_B[184][0] +
                mat_A[30][0] * mat_B[192][0] +
                mat_A[30][1] * mat_B[200][0] +
                mat_A[30][2] * mat_B[208][0] +
                mat_A[30][3] * mat_B[216][0] +
                mat_A[31][0] * mat_B[224][0] +
                mat_A[31][1] * mat_B[232][0] +
                mat_A[31][2] * mat_B[240][0] +
                mat_A[31][3] * mat_B[248][0];
    mat_C[24][1] <=
                mat_A[24][0] * mat_B[0][1] +
                mat_A[24][1] * mat_B[8][1] +
                mat_A[24][2] * mat_B[16][1] +
                mat_A[24][3] * mat_B[24][1] +
                mat_A[25][0] * mat_B[32][1] +
                mat_A[25][1] * mat_B[40][1] +
                mat_A[25][2] * mat_B[48][1] +
                mat_A[25][3] * mat_B[56][1] +
                mat_A[26][0] * mat_B[64][1] +
                mat_A[26][1] * mat_B[72][1] +
                mat_A[26][2] * mat_B[80][1] +
                mat_A[26][3] * mat_B[88][1] +
                mat_A[27][0] * mat_B[96][1] +
                mat_A[27][1] * mat_B[104][1] +
                mat_A[27][2] * mat_B[112][1] +
                mat_A[27][3] * mat_B[120][1] +
                mat_A[28][0] * mat_B[128][1] +
                mat_A[28][1] * mat_B[136][1] +
                mat_A[28][2] * mat_B[144][1] +
                mat_A[28][3] * mat_B[152][1] +
                mat_A[29][0] * mat_B[160][1] +
                mat_A[29][1] * mat_B[168][1] +
                mat_A[29][2] * mat_B[176][1] +
                mat_A[29][3] * mat_B[184][1] +
                mat_A[30][0] * mat_B[192][1] +
                mat_A[30][1] * mat_B[200][1] +
                mat_A[30][2] * mat_B[208][1] +
                mat_A[30][3] * mat_B[216][1] +
                mat_A[31][0] * mat_B[224][1] +
                mat_A[31][1] * mat_B[232][1] +
                mat_A[31][2] * mat_B[240][1] +
                mat_A[31][3] * mat_B[248][1];
    mat_C[24][2] <=
                mat_A[24][0] * mat_B[0][2] +
                mat_A[24][1] * mat_B[8][2] +
                mat_A[24][2] * mat_B[16][2] +
                mat_A[24][3] * mat_B[24][2] +
                mat_A[25][0] * mat_B[32][2] +
                mat_A[25][1] * mat_B[40][2] +
                mat_A[25][2] * mat_B[48][2] +
                mat_A[25][3] * mat_B[56][2] +
                mat_A[26][0] * mat_B[64][2] +
                mat_A[26][1] * mat_B[72][2] +
                mat_A[26][2] * mat_B[80][2] +
                mat_A[26][3] * mat_B[88][2] +
                mat_A[27][0] * mat_B[96][2] +
                mat_A[27][1] * mat_B[104][2] +
                mat_A[27][2] * mat_B[112][2] +
                mat_A[27][3] * mat_B[120][2] +
                mat_A[28][0] * mat_B[128][2] +
                mat_A[28][1] * mat_B[136][2] +
                mat_A[28][2] * mat_B[144][2] +
                mat_A[28][3] * mat_B[152][2] +
                mat_A[29][0] * mat_B[160][2] +
                mat_A[29][1] * mat_B[168][2] +
                mat_A[29][2] * mat_B[176][2] +
                mat_A[29][3] * mat_B[184][2] +
                mat_A[30][0] * mat_B[192][2] +
                mat_A[30][1] * mat_B[200][2] +
                mat_A[30][2] * mat_B[208][2] +
                mat_A[30][3] * mat_B[216][2] +
                mat_A[31][0] * mat_B[224][2] +
                mat_A[31][1] * mat_B[232][2] +
                mat_A[31][2] * mat_B[240][2] +
                mat_A[31][3] * mat_B[248][2];
    mat_C[24][3] <=
                mat_A[24][0] * mat_B[0][3] +
                mat_A[24][1] * mat_B[8][3] +
                mat_A[24][2] * mat_B[16][3] +
                mat_A[24][3] * mat_B[24][3] +
                mat_A[25][0] * mat_B[32][3] +
                mat_A[25][1] * mat_B[40][3] +
                mat_A[25][2] * mat_B[48][3] +
                mat_A[25][3] * mat_B[56][3] +
                mat_A[26][0] * mat_B[64][3] +
                mat_A[26][1] * mat_B[72][3] +
                mat_A[26][2] * mat_B[80][3] +
                mat_A[26][3] * mat_B[88][3] +
                mat_A[27][0] * mat_B[96][3] +
                mat_A[27][1] * mat_B[104][3] +
                mat_A[27][2] * mat_B[112][3] +
                mat_A[27][3] * mat_B[120][3] +
                mat_A[28][0] * mat_B[128][3] +
                mat_A[28][1] * mat_B[136][3] +
                mat_A[28][2] * mat_B[144][3] +
                mat_A[28][3] * mat_B[152][3] +
                mat_A[29][0] * mat_B[160][3] +
                mat_A[29][1] * mat_B[168][3] +
                mat_A[29][2] * mat_B[176][3] +
                mat_A[29][3] * mat_B[184][3] +
                mat_A[30][0] * mat_B[192][3] +
                mat_A[30][1] * mat_B[200][3] +
                mat_A[30][2] * mat_B[208][3] +
                mat_A[30][3] * mat_B[216][3] +
                mat_A[31][0] * mat_B[224][3] +
                mat_A[31][1] * mat_B[232][3] +
                mat_A[31][2] * mat_B[240][3] +
                mat_A[31][3] * mat_B[248][3];
    mat_C[25][0] <=
                mat_A[24][0] * mat_B[1][0] +
                mat_A[24][1] * mat_B[9][0] +
                mat_A[24][2] * mat_B[17][0] +
                mat_A[24][3] * mat_B[25][0] +
                mat_A[25][0] * mat_B[33][0] +
                mat_A[25][1] * mat_B[41][0] +
                mat_A[25][2] * mat_B[49][0] +
                mat_A[25][3] * mat_B[57][0] +
                mat_A[26][0] * mat_B[65][0] +
                mat_A[26][1] * mat_B[73][0] +
                mat_A[26][2] * mat_B[81][0] +
                mat_A[26][3] * mat_B[89][0] +
                mat_A[27][0] * mat_B[97][0] +
                mat_A[27][1] * mat_B[105][0] +
                mat_A[27][2] * mat_B[113][0] +
                mat_A[27][3] * mat_B[121][0] +
                mat_A[28][0] * mat_B[129][0] +
                mat_A[28][1] * mat_B[137][0] +
                mat_A[28][2] * mat_B[145][0] +
                mat_A[28][3] * mat_B[153][0] +
                mat_A[29][0] * mat_B[161][0] +
                mat_A[29][1] * mat_B[169][0] +
                mat_A[29][2] * mat_B[177][0] +
                mat_A[29][3] * mat_B[185][0] +
                mat_A[30][0] * mat_B[193][0] +
                mat_A[30][1] * mat_B[201][0] +
                mat_A[30][2] * mat_B[209][0] +
                mat_A[30][3] * mat_B[217][0] +
                mat_A[31][0] * mat_B[225][0] +
                mat_A[31][1] * mat_B[233][0] +
                mat_A[31][2] * mat_B[241][0] +
                mat_A[31][3] * mat_B[249][0];
    mat_C[25][1] <=
                mat_A[24][0] * mat_B[1][1] +
                mat_A[24][1] * mat_B[9][1] +
                mat_A[24][2] * mat_B[17][1] +
                mat_A[24][3] * mat_B[25][1] +
                mat_A[25][0] * mat_B[33][1] +
                mat_A[25][1] * mat_B[41][1] +
                mat_A[25][2] * mat_B[49][1] +
                mat_A[25][3] * mat_B[57][1] +
                mat_A[26][0] * mat_B[65][1] +
                mat_A[26][1] * mat_B[73][1] +
                mat_A[26][2] * mat_B[81][1] +
                mat_A[26][3] * mat_B[89][1] +
                mat_A[27][0] * mat_B[97][1] +
                mat_A[27][1] * mat_B[105][1] +
                mat_A[27][2] * mat_B[113][1] +
                mat_A[27][3] * mat_B[121][1] +
                mat_A[28][0] * mat_B[129][1] +
                mat_A[28][1] * mat_B[137][1] +
                mat_A[28][2] * mat_B[145][1] +
                mat_A[28][3] * mat_B[153][1] +
                mat_A[29][0] * mat_B[161][1] +
                mat_A[29][1] * mat_B[169][1] +
                mat_A[29][2] * mat_B[177][1] +
                mat_A[29][3] * mat_B[185][1] +
                mat_A[30][0] * mat_B[193][1] +
                mat_A[30][1] * mat_B[201][1] +
                mat_A[30][2] * mat_B[209][1] +
                mat_A[30][3] * mat_B[217][1] +
                mat_A[31][0] * mat_B[225][1] +
                mat_A[31][1] * mat_B[233][1] +
                mat_A[31][2] * mat_B[241][1] +
                mat_A[31][3] * mat_B[249][1];
    mat_C[25][2] <=
                mat_A[24][0] * mat_B[1][2] +
                mat_A[24][1] * mat_B[9][2] +
                mat_A[24][2] * mat_B[17][2] +
                mat_A[24][3] * mat_B[25][2] +
                mat_A[25][0] * mat_B[33][2] +
                mat_A[25][1] * mat_B[41][2] +
                mat_A[25][2] * mat_B[49][2] +
                mat_A[25][3] * mat_B[57][2] +
                mat_A[26][0] * mat_B[65][2] +
                mat_A[26][1] * mat_B[73][2] +
                mat_A[26][2] * mat_B[81][2] +
                mat_A[26][3] * mat_B[89][2] +
                mat_A[27][0] * mat_B[97][2] +
                mat_A[27][1] * mat_B[105][2] +
                mat_A[27][2] * mat_B[113][2] +
                mat_A[27][3] * mat_B[121][2] +
                mat_A[28][0] * mat_B[129][2] +
                mat_A[28][1] * mat_B[137][2] +
                mat_A[28][2] * mat_B[145][2] +
                mat_A[28][3] * mat_B[153][2] +
                mat_A[29][0] * mat_B[161][2] +
                mat_A[29][1] * mat_B[169][2] +
                mat_A[29][2] * mat_B[177][2] +
                mat_A[29][3] * mat_B[185][2] +
                mat_A[30][0] * mat_B[193][2] +
                mat_A[30][1] * mat_B[201][2] +
                mat_A[30][2] * mat_B[209][2] +
                mat_A[30][3] * mat_B[217][2] +
                mat_A[31][0] * mat_B[225][2] +
                mat_A[31][1] * mat_B[233][2] +
                mat_A[31][2] * mat_B[241][2] +
                mat_A[31][3] * mat_B[249][2];
    mat_C[25][3] <=
                mat_A[24][0] * mat_B[1][3] +
                mat_A[24][1] * mat_B[9][3] +
                mat_A[24][2] * mat_B[17][3] +
                mat_A[24][3] * mat_B[25][3] +
                mat_A[25][0] * mat_B[33][3] +
                mat_A[25][1] * mat_B[41][3] +
                mat_A[25][2] * mat_B[49][3] +
                mat_A[25][3] * mat_B[57][3] +
                mat_A[26][0] * mat_B[65][3] +
                mat_A[26][1] * mat_B[73][3] +
                mat_A[26][2] * mat_B[81][3] +
                mat_A[26][3] * mat_B[89][3] +
                mat_A[27][0] * mat_B[97][3] +
                mat_A[27][1] * mat_B[105][3] +
                mat_A[27][2] * mat_B[113][3] +
                mat_A[27][3] * mat_B[121][3] +
                mat_A[28][0] * mat_B[129][3] +
                mat_A[28][1] * mat_B[137][3] +
                mat_A[28][2] * mat_B[145][3] +
                mat_A[28][3] * mat_B[153][3] +
                mat_A[29][0] * mat_B[161][3] +
                mat_A[29][1] * mat_B[169][3] +
                mat_A[29][2] * mat_B[177][3] +
                mat_A[29][3] * mat_B[185][3] +
                mat_A[30][0] * mat_B[193][3] +
                mat_A[30][1] * mat_B[201][3] +
                mat_A[30][2] * mat_B[209][3] +
                mat_A[30][3] * mat_B[217][3] +
                mat_A[31][0] * mat_B[225][3] +
                mat_A[31][1] * mat_B[233][3] +
                mat_A[31][2] * mat_B[241][3] +
                mat_A[31][3] * mat_B[249][3];
    mat_C[26][0] <=
                mat_A[24][0] * mat_B[2][0] +
                mat_A[24][1] * mat_B[10][0] +
                mat_A[24][2] * mat_B[18][0] +
                mat_A[24][3] * mat_B[26][0] +
                mat_A[25][0] * mat_B[34][0] +
                mat_A[25][1] * mat_B[42][0] +
                mat_A[25][2] * mat_B[50][0] +
                mat_A[25][3] * mat_B[58][0] +
                mat_A[26][0] * mat_B[66][0] +
                mat_A[26][1] * mat_B[74][0] +
                mat_A[26][2] * mat_B[82][0] +
                mat_A[26][3] * mat_B[90][0] +
                mat_A[27][0] * mat_B[98][0] +
                mat_A[27][1] * mat_B[106][0] +
                mat_A[27][2] * mat_B[114][0] +
                mat_A[27][3] * mat_B[122][0] +
                mat_A[28][0] * mat_B[130][0] +
                mat_A[28][1] * mat_B[138][0] +
                mat_A[28][2] * mat_B[146][0] +
                mat_A[28][3] * mat_B[154][0] +
                mat_A[29][0] * mat_B[162][0] +
                mat_A[29][1] * mat_B[170][0] +
                mat_A[29][2] * mat_B[178][0] +
                mat_A[29][3] * mat_B[186][0] +
                mat_A[30][0] * mat_B[194][0] +
                mat_A[30][1] * mat_B[202][0] +
                mat_A[30][2] * mat_B[210][0] +
                mat_A[30][3] * mat_B[218][0] +
                mat_A[31][0] * mat_B[226][0] +
                mat_A[31][1] * mat_B[234][0] +
                mat_A[31][2] * mat_B[242][0] +
                mat_A[31][3] * mat_B[250][0];
    mat_C[26][1] <=
                mat_A[24][0] * mat_B[2][1] +
                mat_A[24][1] * mat_B[10][1] +
                mat_A[24][2] * mat_B[18][1] +
                mat_A[24][3] * mat_B[26][1] +
                mat_A[25][0] * mat_B[34][1] +
                mat_A[25][1] * mat_B[42][1] +
                mat_A[25][2] * mat_B[50][1] +
                mat_A[25][3] * mat_B[58][1] +
                mat_A[26][0] * mat_B[66][1] +
                mat_A[26][1] * mat_B[74][1] +
                mat_A[26][2] * mat_B[82][1] +
                mat_A[26][3] * mat_B[90][1] +
                mat_A[27][0] * mat_B[98][1] +
                mat_A[27][1] * mat_B[106][1] +
                mat_A[27][2] * mat_B[114][1] +
                mat_A[27][3] * mat_B[122][1] +
                mat_A[28][0] * mat_B[130][1] +
                mat_A[28][1] * mat_B[138][1] +
                mat_A[28][2] * mat_B[146][1] +
                mat_A[28][3] * mat_B[154][1] +
                mat_A[29][0] * mat_B[162][1] +
                mat_A[29][1] * mat_B[170][1] +
                mat_A[29][2] * mat_B[178][1] +
                mat_A[29][3] * mat_B[186][1] +
                mat_A[30][0] * mat_B[194][1] +
                mat_A[30][1] * mat_B[202][1] +
                mat_A[30][2] * mat_B[210][1] +
                mat_A[30][3] * mat_B[218][1] +
                mat_A[31][0] * mat_B[226][1] +
                mat_A[31][1] * mat_B[234][1] +
                mat_A[31][2] * mat_B[242][1] +
                mat_A[31][3] * mat_B[250][1];
    mat_C[26][2] <=
                mat_A[24][0] * mat_B[2][2] +
                mat_A[24][1] * mat_B[10][2] +
                mat_A[24][2] * mat_B[18][2] +
                mat_A[24][3] * mat_B[26][2] +
                mat_A[25][0] * mat_B[34][2] +
                mat_A[25][1] * mat_B[42][2] +
                mat_A[25][2] * mat_B[50][2] +
                mat_A[25][3] * mat_B[58][2] +
                mat_A[26][0] * mat_B[66][2] +
                mat_A[26][1] * mat_B[74][2] +
                mat_A[26][2] * mat_B[82][2] +
                mat_A[26][3] * mat_B[90][2] +
                mat_A[27][0] * mat_B[98][2] +
                mat_A[27][1] * mat_B[106][2] +
                mat_A[27][2] * mat_B[114][2] +
                mat_A[27][3] * mat_B[122][2] +
                mat_A[28][0] * mat_B[130][2] +
                mat_A[28][1] * mat_B[138][2] +
                mat_A[28][2] * mat_B[146][2] +
                mat_A[28][3] * mat_B[154][2] +
                mat_A[29][0] * mat_B[162][2] +
                mat_A[29][1] * mat_B[170][2] +
                mat_A[29][2] * mat_B[178][2] +
                mat_A[29][3] * mat_B[186][2] +
                mat_A[30][0] * mat_B[194][2] +
                mat_A[30][1] * mat_B[202][2] +
                mat_A[30][2] * mat_B[210][2] +
                mat_A[30][3] * mat_B[218][2] +
                mat_A[31][0] * mat_B[226][2] +
                mat_A[31][1] * mat_B[234][2] +
                mat_A[31][2] * mat_B[242][2] +
                mat_A[31][3] * mat_B[250][2];
    mat_C[26][3] <=
                mat_A[24][0] * mat_B[2][3] +
                mat_A[24][1] * mat_B[10][3] +
                mat_A[24][2] * mat_B[18][3] +
                mat_A[24][3] * mat_B[26][3] +
                mat_A[25][0] * mat_B[34][3] +
                mat_A[25][1] * mat_B[42][3] +
                mat_A[25][2] * mat_B[50][3] +
                mat_A[25][3] * mat_B[58][3] +
                mat_A[26][0] * mat_B[66][3] +
                mat_A[26][1] * mat_B[74][3] +
                mat_A[26][2] * mat_B[82][3] +
                mat_A[26][3] * mat_B[90][3] +
                mat_A[27][0] * mat_B[98][3] +
                mat_A[27][1] * mat_B[106][3] +
                mat_A[27][2] * mat_B[114][3] +
                mat_A[27][3] * mat_B[122][3] +
                mat_A[28][0] * mat_B[130][3] +
                mat_A[28][1] * mat_B[138][3] +
                mat_A[28][2] * mat_B[146][3] +
                mat_A[28][3] * mat_B[154][3] +
                mat_A[29][0] * mat_B[162][3] +
                mat_A[29][1] * mat_B[170][3] +
                mat_A[29][2] * mat_B[178][3] +
                mat_A[29][3] * mat_B[186][3] +
                mat_A[30][0] * mat_B[194][3] +
                mat_A[30][1] * mat_B[202][3] +
                mat_A[30][2] * mat_B[210][3] +
                mat_A[30][3] * mat_B[218][3] +
                mat_A[31][0] * mat_B[226][3] +
                mat_A[31][1] * mat_B[234][3] +
                mat_A[31][2] * mat_B[242][3] +
                mat_A[31][3] * mat_B[250][3];
    mat_C[27][0] <=
                mat_A[24][0] * mat_B[3][0] +
                mat_A[24][1] * mat_B[11][0] +
                mat_A[24][2] * mat_B[19][0] +
                mat_A[24][3] * mat_B[27][0] +
                mat_A[25][0] * mat_B[35][0] +
                mat_A[25][1] * mat_B[43][0] +
                mat_A[25][2] * mat_B[51][0] +
                mat_A[25][3] * mat_B[59][0] +
                mat_A[26][0] * mat_B[67][0] +
                mat_A[26][1] * mat_B[75][0] +
                mat_A[26][2] * mat_B[83][0] +
                mat_A[26][3] * mat_B[91][0] +
                mat_A[27][0] * mat_B[99][0] +
                mat_A[27][1] * mat_B[107][0] +
                mat_A[27][2] * mat_B[115][0] +
                mat_A[27][3] * mat_B[123][0] +
                mat_A[28][0] * mat_B[131][0] +
                mat_A[28][1] * mat_B[139][0] +
                mat_A[28][2] * mat_B[147][0] +
                mat_A[28][3] * mat_B[155][0] +
                mat_A[29][0] * mat_B[163][0] +
                mat_A[29][1] * mat_B[171][0] +
                mat_A[29][2] * mat_B[179][0] +
                mat_A[29][3] * mat_B[187][0] +
                mat_A[30][0] * mat_B[195][0] +
                mat_A[30][1] * mat_B[203][0] +
                mat_A[30][2] * mat_B[211][0] +
                mat_A[30][3] * mat_B[219][0] +
                mat_A[31][0] * mat_B[227][0] +
                mat_A[31][1] * mat_B[235][0] +
                mat_A[31][2] * mat_B[243][0] +
                mat_A[31][3] * mat_B[251][0];
    mat_C[27][1] <=
                mat_A[24][0] * mat_B[3][1] +
                mat_A[24][1] * mat_B[11][1] +
                mat_A[24][2] * mat_B[19][1] +
                mat_A[24][3] * mat_B[27][1] +
                mat_A[25][0] * mat_B[35][1] +
                mat_A[25][1] * mat_B[43][1] +
                mat_A[25][2] * mat_B[51][1] +
                mat_A[25][3] * mat_B[59][1] +
                mat_A[26][0] * mat_B[67][1] +
                mat_A[26][1] * mat_B[75][1] +
                mat_A[26][2] * mat_B[83][1] +
                mat_A[26][3] * mat_B[91][1] +
                mat_A[27][0] * mat_B[99][1] +
                mat_A[27][1] * mat_B[107][1] +
                mat_A[27][2] * mat_B[115][1] +
                mat_A[27][3] * mat_B[123][1] +
                mat_A[28][0] * mat_B[131][1] +
                mat_A[28][1] * mat_B[139][1] +
                mat_A[28][2] * mat_B[147][1] +
                mat_A[28][3] * mat_B[155][1] +
                mat_A[29][0] * mat_B[163][1] +
                mat_A[29][1] * mat_B[171][1] +
                mat_A[29][2] * mat_B[179][1] +
                mat_A[29][3] * mat_B[187][1] +
                mat_A[30][0] * mat_B[195][1] +
                mat_A[30][1] * mat_B[203][1] +
                mat_A[30][2] * mat_B[211][1] +
                mat_A[30][3] * mat_B[219][1] +
                mat_A[31][0] * mat_B[227][1] +
                mat_A[31][1] * mat_B[235][1] +
                mat_A[31][2] * mat_B[243][1] +
                mat_A[31][3] * mat_B[251][1];
    mat_C[27][2] <=
                mat_A[24][0] * mat_B[3][2] +
                mat_A[24][1] * mat_B[11][2] +
                mat_A[24][2] * mat_B[19][2] +
                mat_A[24][3] * mat_B[27][2] +
                mat_A[25][0] * mat_B[35][2] +
                mat_A[25][1] * mat_B[43][2] +
                mat_A[25][2] * mat_B[51][2] +
                mat_A[25][3] * mat_B[59][2] +
                mat_A[26][0] * mat_B[67][2] +
                mat_A[26][1] * mat_B[75][2] +
                mat_A[26][2] * mat_B[83][2] +
                mat_A[26][3] * mat_B[91][2] +
                mat_A[27][0] * mat_B[99][2] +
                mat_A[27][1] * mat_B[107][2] +
                mat_A[27][2] * mat_B[115][2] +
                mat_A[27][3] * mat_B[123][2] +
                mat_A[28][0] * mat_B[131][2] +
                mat_A[28][1] * mat_B[139][2] +
                mat_A[28][2] * mat_B[147][2] +
                mat_A[28][3] * mat_B[155][2] +
                mat_A[29][0] * mat_B[163][2] +
                mat_A[29][1] * mat_B[171][2] +
                mat_A[29][2] * mat_B[179][2] +
                mat_A[29][3] * mat_B[187][2] +
                mat_A[30][0] * mat_B[195][2] +
                mat_A[30][1] * mat_B[203][2] +
                mat_A[30][2] * mat_B[211][2] +
                mat_A[30][3] * mat_B[219][2] +
                mat_A[31][0] * mat_B[227][2] +
                mat_A[31][1] * mat_B[235][2] +
                mat_A[31][2] * mat_B[243][2] +
                mat_A[31][3] * mat_B[251][2];
    mat_C[27][3] <=
                mat_A[24][0] * mat_B[3][3] +
                mat_A[24][1] * mat_B[11][3] +
                mat_A[24][2] * mat_B[19][3] +
                mat_A[24][3] * mat_B[27][3] +
                mat_A[25][0] * mat_B[35][3] +
                mat_A[25][1] * mat_B[43][3] +
                mat_A[25][2] * mat_B[51][3] +
                mat_A[25][3] * mat_B[59][3] +
                mat_A[26][0] * mat_B[67][3] +
                mat_A[26][1] * mat_B[75][3] +
                mat_A[26][2] * mat_B[83][3] +
                mat_A[26][3] * mat_B[91][3] +
                mat_A[27][0] * mat_B[99][3] +
                mat_A[27][1] * mat_B[107][3] +
                mat_A[27][2] * mat_B[115][3] +
                mat_A[27][3] * mat_B[123][3] +
                mat_A[28][0] * mat_B[131][3] +
                mat_A[28][1] * mat_B[139][3] +
                mat_A[28][2] * mat_B[147][3] +
                mat_A[28][3] * mat_B[155][3] +
                mat_A[29][0] * mat_B[163][3] +
                mat_A[29][1] * mat_B[171][3] +
                mat_A[29][2] * mat_B[179][3] +
                mat_A[29][3] * mat_B[187][3] +
                mat_A[30][0] * mat_B[195][3] +
                mat_A[30][1] * mat_B[203][3] +
                mat_A[30][2] * mat_B[211][3] +
                mat_A[30][3] * mat_B[219][3] +
                mat_A[31][0] * mat_B[227][3] +
                mat_A[31][1] * mat_B[235][3] +
                mat_A[31][2] * mat_B[243][3] +
                mat_A[31][3] * mat_B[251][3];
    mat_C[28][0] <=
                mat_A[24][0] * mat_B[4][0] +
                mat_A[24][1] * mat_B[12][0] +
                mat_A[24][2] * mat_B[20][0] +
                mat_A[24][3] * mat_B[28][0] +
                mat_A[25][0] * mat_B[36][0] +
                mat_A[25][1] * mat_B[44][0] +
                mat_A[25][2] * mat_B[52][0] +
                mat_A[25][3] * mat_B[60][0] +
                mat_A[26][0] * mat_B[68][0] +
                mat_A[26][1] * mat_B[76][0] +
                mat_A[26][2] * mat_B[84][0] +
                mat_A[26][3] * mat_B[92][0] +
                mat_A[27][0] * mat_B[100][0] +
                mat_A[27][1] * mat_B[108][0] +
                mat_A[27][2] * mat_B[116][0] +
                mat_A[27][3] * mat_B[124][0] +
                mat_A[28][0] * mat_B[132][0] +
                mat_A[28][1] * mat_B[140][0] +
                mat_A[28][2] * mat_B[148][0] +
                mat_A[28][3] * mat_B[156][0] +
                mat_A[29][0] * mat_B[164][0] +
                mat_A[29][1] * mat_B[172][0] +
                mat_A[29][2] * mat_B[180][0] +
                mat_A[29][3] * mat_B[188][0] +
                mat_A[30][0] * mat_B[196][0] +
                mat_A[30][1] * mat_B[204][0] +
                mat_A[30][2] * mat_B[212][0] +
                mat_A[30][3] * mat_B[220][0] +
                mat_A[31][0] * mat_B[228][0] +
                mat_A[31][1] * mat_B[236][0] +
                mat_A[31][2] * mat_B[244][0] +
                mat_A[31][3] * mat_B[252][0];
    mat_C[28][1] <=
                mat_A[24][0] * mat_B[4][1] +
                mat_A[24][1] * mat_B[12][1] +
                mat_A[24][2] * mat_B[20][1] +
                mat_A[24][3] * mat_B[28][1] +
                mat_A[25][0] * mat_B[36][1] +
                mat_A[25][1] * mat_B[44][1] +
                mat_A[25][2] * mat_B[52][1] +
                mat_A[25][3] * mat_B[60][1] +
                mat_A[26][0] * mat_B[68][1] +
                mat_A[26][1] * mat_B[76][1] +
                mat_A[26][2] * mat_B[84][1] +
                mat_A[26][3] * mat_B[92][1] +
                mat_A[27][0] * mat_B[100][1] +
                mat_A[27][1] * mat_B[108][1] +
                mat_A[27][2] * mat_B[116][1] +
                mat_A[27][3] * mat_B[124][1] +
                mat_A[28][0] * mat_B[132][1] +
                mat_A[28][1] * mat_B[140][1] +
                mat_A[28][2] * mat_B[148][1] +
                mat_A[28][3] * mat_B[156][1] +
                mat_A[29][0] * mat_B[164][1] +
                mat_A[29][1] * mat_B[172][1] +
                mat_A[29][2] * mat_B[180][1] +
                mat_A[29][3] * mat_B[188][1] +
                mat_A[30][0] * mat_B[196][1] +
                mat_A[30][1] * mat_B[204][1] +
                mat_A[30][2] * mat_B[212][1] +
                mat_A[30][3] * mat_B[220][1] +
                mat_A[31][0] * mat_B[228][1] +
                mat_A[31][1] * mat_B[236][1] +
                mat_A[31][2] * mat_B[244][1] +
                mat_A[31][3] * mat_B[252][1];
    mat_C[28][2] <=
                mat_A[24][0] * mat_B[4][2] +
                mat_A[24][1] * mat_B[12][2] +
                mat_A[24][2] * mat_B[20][2] +
                mat_A[24][3] * mat_B[28][2] +
                mat_A[25][0] * mat_B[36][2] +
                mat_A[25][1] * mat_B[44][2] +
                mat_A[25][2] * mat_B[52][2] +
                mat_A[25][3] * mat_B[60][2] +
                mat_A[26][0] * mat_B[68][2] +
                mat_A[26][1] * mat_B[76][2] +
                mat_A[26][2] * mat_B[84][2] +
                mat_A[26][3] * mat_B[92][2] +
                mat_A[27][0] * mat_B[100][2] +
                mat_A[27][1] * mat_B[108][2] +
                mat_A[27][2] * mat_B[116][2] +
                mat_A[27][3] * mat_B[124][2] +
                mat_A[28][0] * mat_B[132][2] +
                mat_A[28][1] * mat_B[140][2] +
                mat_A[28][2] * mat_B[148][2] +
                mat_A[28][3] * mat_B[156][2] +
                mat_A[29][0] * mat_B[164][2] +
                mat_A[29][1] * mat_B[172][2] +
                mat_A[29][2] * mat_B[180][2] +
                mat_A[29][3] * mat_B[188][2] +
                mat_A[30][0] * mat_B[196][2] +
                mat_A[30][1] * mat_B[204][2] +
                mat_A[30][2] * mat_B[212][2] +
                mat_A[30][3] * mat_B[220][2] +
                mat_A[31][0] * mat_B[228][2] +
                mat_A[31][1] * mat_B[236][2] +
                mat_A[31][2] * mat_B[244][2] +
                mat_A[31][3] * mat_B[252][2];
    mat_C[28][3] <=
                mat_A[24][0] * mat_B[4][3] +
                mat_A[24][1] * mat_B[12][3] +
                mat_A[24][2] * mat_B[20][3] +
                mat_A[24][3] * mat_B[28][3] +
                mat_A[25][0] * mat_B[36][3] +
                mat_A[25][1] * mat_B[44][3] +
                mat_A[25][2] * mat_B[52][3] +
                mat_A[25][3] * mat_B[60][3] +
                mat_A[26][0] * mat_B[68][3] +
                mat_A[26][1] * mat_B[76][3] +
                mat_A[26][2] * mat_B[84][3] +
                mat_A[26][3] * mat_B[92][3] +
                mat_A[27][0] * mat_B[100][3] +
                mat_A[27][1] * mat_B[108][3] +
                mat_A[27][2] * mat_B[116][3] +
                mat_A[27][3] * mat_B[124][3] +
                mat_A[28][0] * mat_B[132][3] +
                mat_A[28][1] * mat_B[140][3] +
                mat_A[28][2] * mat_B[148][3] +
                mat_A[28][3] * mat_B[156][3] +
                mat_A[29][0] * mat_B[164][3] +
                mat_A[29][1] * mat_B[172][3] +
                mat_A[29][2] * mat_B[180][3] +
                mat_A[29][3] * mat_B[188][3] +
                mat_A[30][0] * mat_B[196][3] +
                mat_A[30][1] * mat_B[204][3] +
                mat_A[30][2] * mat_B[212][3] +
                mat_A[30][3] * mat_B[220][3] +
                mat_A[31][0] * mat_B[228][3] +
                mat_A[31][1] * mat_B[236][3] +
                mat_A[31][2] * mat_B[244][3] +
                mat_A[31][3] * mat_B[252][3];
    mat_C[29][0] <=
                mat_A[24][0] * mat_B[5][0] +
                mat_A[24][1] * mat_B[13][0] +
                mat_A[24][2] * mat_B[21][0] +
                mat_A[24][3] * mat_B[29][0] +
                mat_A[25][0] * mat_B[37][0] +
                mat_A[25][1] * mat_B[45][0] +
                mat_A[25][2] * mat_B[53][0] +
                mat_A[25][3] * mat_B[61][0] +
                mat_A[26][0] * mat_B[69][0] +
                mat_A[26][1] * mat_B[77][0] +
                mat_A[26][2] * mat_B[85][0] +
                mat_A[26][3] * mat_B[93][0] +
                mat_A[27][0] * mat_B[101][0] +
                mat_A[27][1] * mat_B[109][0] +
                mat_A[27][2] * mat_B[117][0] +
                mat_A[27][3] * mat_B[125][0] +
                mat_A[28][0] * mat_B[133][0] +
                mat_A[28][1] * mat_B[141][0] +
                mat_A[28][2] * mat_B[149][0] +
                mat_A[28][3] * mat_B[157][0] +
                mat_A[29][0] * mat_B[165][0] +
                mat_A[29][1] * mat_B[173][0] +
                mat_A[29][2] * mat_B[181][0] +
                mat_A[29][3] * mat_B[189][0] +
                mat_A[30][0] * mat_B[197][0] +
                mat_A[30][1] * mat_B[205][0] +
                mat_A[30][2] * mat_B[213][0] +
                mat_A[30][3] * mat_B[221][0] +
                mat_A[31][0] * mat_B[229][0] +
                mat_A[31][1] * mat_B[237][0] +
                mat_A[31][2] * mat_B[245][0] +
                mat_A[31][3] * mat_B[253][0];
    mat_C[29][1] <=
                mat_A[24][0] * mat_B[5][1] +
                mat_A[24][1] * mat_B[13][1] +
                mat_A[24][2] * mat_B[21][1] +
                mat_A[24][3] * mat_B[29][1] +
                mat_A[25][0] * mat_B[37][1] +
                mat_A[25][1] * mat_B[45][1] +
                mat_A[25][2] * mat_B[53][1] +
                mat_A[25][3] * mat_B[61][1] +
                mat_A[26][0] * mat_B[69][1] +
                mat_A[26][1] * mat_B[77][1] +
                mat_A[26][2] * mat_B[85][1] +
                mat_A[26][3] * mat_B[93][1] +
                mat_A[27][0] * mat_B[101][1] +
                mat_A[27][1] * mat_B[109][1] +
                mat_A[27][2] * mat_B[117][1] +
                mat_A[27][3] * mat_B[125][1] +
                mat_A[28][0] * mat_B[133][1] +
                mat_A[28][1] * mat_B[141][1] +
                mat_A[28][2] * mat_B[149][1] +
                mat_A[28][3] * mat_B[157][1] +
                mat_A[29][0] * mat_B[165][1] +
                mat_A[29][1] * mat_B[173][1] +
                mat_A[29][2] * mat_B[181][1] +
                mat_A[29][3] * mat_B[189][1] +
                mat_A[30][0] * mat_B[197][1] +
                mat_A[30][1] * mat_B[205][1] +
                mat_A[30][2] * mat_B[213][1] +
                mat_A[30][3] * mat_B[221][1] +
                mat_A[31][0] * mat_B[229][1] +
                mat_A[31][1] * mat_B[237][1] +
                mat_A[31][2] * mat_B[245][1] +
                mat_A[31][3] * mat_B[253][1];
    mat_C[29][2] <=
                mat_A[24][0] * mat_B[5][2] +
                mat_A[24][1] * mat_B[13][2] +
                mat_A[24][2] * mat_B[21][2] +
                mat_A[24][3] * mat_B[29][2] +
                mat_A[25][0] * mat_B[37][2] +
                mat_A[25][1] * mat_B[45][2] +
                mat_A[25][2] * mat_B[53][2] +
                mat_A[25][3] * mat_B[61][2] +
                mat_A[26][0] * mat_B[69][2] +
                mat_A[26][1] * mat_B[77][2] +
                mat_A[26][2] * mat_B[85][2] +
                mat_A[26][3] * mat_B[93][2] +
                mat_A[27][0] * mat_B[101][2] +
                mat_A[27][1] * mat_B[109][2] +
                mat_A[27][2] * mat_B[117][2] +
                mat_A[27][3] * mat_B[125][2] +
                mat_A[28][0] * mat_B[133][2] +
                mat_A[28][1] * mat_B[141][2] +
                mat_A[28][2] * mat_B[149][2] +
                mat_A[28][3] * mat_B[157][2] +
                mat_A[29][0] * mat_B[165][2] +
                mat_A[29][1] * mat_B[173][2] +
                mat_A[29][2] * mat_B[181][2] +
                mat_A[29][3] * mat_B[189][2] +
                mat_A[30][0] * mat_B[197][2] +
                mat_A[30][1] * mat_B[205][2] +
                mat_A[30][2] * mat_B[213][2] +
                mat_A[30][3] * mat_B[221][2] +
                mat_A[31][0] * mat_B[229][2] +
                mat_A[31][1] * mat_B[237][2] +
                mat_A[31][2] * mat_B[245][2] +
                mat_A[31][3] * mat_B[253][2];
    mat_C[29][3] <=
                mat_A[24][0] * mat_B[5][3] +
                mat_A[24][1] * mat_B[13][3] +
                mat_A[24][2] * mat_B[21][3] +
                mat_A[24][3] * mat_B[29][3] +
                mat_A[25][0] * mat_B[37][3] +
                mat_A[25][1] * mat_B[45][3] +
                mat_A[25][2] * mat_B[53][3] +
                mat_A[25][3] * mat_B[61][3] +
                mat_A[26][0] * mat_B[69][3] +
                mat_A[26][1] * mat_B[77][3] +
                mat_A[26][2] * mat_B[85][3] +
                mat_A[26][3] * mat_B[93][3] +
                mat_A[27][0] * mat_B[101][3] +
                mat_A[27][1] * mat_B[109][3] +
                mat_A[27][2] * mat_B[117][3] +
                mat_A[27][3] * mat_B[125][3] +
                mat_A[28][0] * mat_B[133][3] +
                mat_A[28][1] * mat_B[141][3] +
                mat_A[28][2] * mat_B[149][3] +
                mat_A[28][3] * mat_B[157][3] +
                mat_A[29][0] * mat_B[165][3] +
                mat_A[29][1] * mat_B[173][3] +
                mat_A[29][2] * mat_B[181][3] +
                mat_A[29][3] * mat_B[189][3] +
                mat_A[30][0] * mat_B[197][3] +
                mat_A[30][1] * mat_B[205][3] +
                mat_A[30][2] * mat_B[213][3] +
                mat_A[30][3] * mat_B[221][3] +
                mat_A[31][0] * mat_B[229][3] +
                mat_A[31][1] * mat_B[237][3] +
                mat_A[31][2] * mat_B[245][3] +
                mat_A[31][3] * mat_B[253][3];
    mat_C[30][0] <=
                mat_A[24][0] * mat_B[6][0] +
                mat_A[24][1] * mat_B[14][0] +
                mat_A[24][2] * mat_B[22][0] +
                mat_A[24][3] * mat_B[30][0] +
                mat_A[25][0] * mat_B[38][0] +
                mat_A[25][1] * mat_B[46][0] +
                mat_A[25][2] * mat_B[54][0] +
                mat_A[25][3] * mat_B[62][0] +
                mat_A[26][0] * mat_B[70][0] +
                mat_A[26][1] * mat_B[78][0] +
                mat_A[26][2] * mat_B[86][0] +
                mat_A[26][3] * mat_B[94][0] +
                mat_A[27][0] * mat_B[102][0] +
                mat_A[27][1] * mat_B[110][0] +
                mat_A[27][2] * mat_B[118][0] +
                mat_A[27][3] * mat_B[126][0] +
                mat_A[28][0] * mat_B[134][0] +
                mat_A[28][1] * mat_B[142][0] +
                mat_A[28][2] * mat_B[150][0] +
                mat_A[28][3] * mat_B[158][0] +
                mat_A[29][0] * mat_B[166][0] +
                mat_A[29][1] * mat_B[174][0] +
                mat_A[29][2] * mat_B[182][0] +
                mat_A[29][3] * mat_B[190][0] +
                mat_A[30][0] * mat_B[198][0] +
                mat_A[30][1] * mat_B[206][0] +
                mat_A[30][2] * mat_B[214][0] +
                mat_A[30][3] * mat_B[222][0] +
                mat_A[31][0] * mat_B[230][0] +
                mat_A[31][1] * mat_B[238][0] +
                mat_A[31][2] * mat_B[246][0] +
                mat_A[31][3] * mat_B[254][0];
    mat_C[30][1] <=
                mat_A[24][0] * mat_B[6][1] +
                mat_A[24][1] * mat_B[14][1] +
                mat_A[24][2] * mat_B[22][1] +
                mat_A[24][3] * mat_B[30][1] +
                mat_A[25][0] * mat_B[38][1] +
                mat_A[25][1] * mat_B[46][1] +
                mat_A[25][2] * mat_B[54][1] +
                mat_A[25][3] * mat_B[62][1] +
                mat_A[26][0] * mat_B[70][1] +
                mat_A[26][1] * mat_B[78][1] +
                mat_A[26][2] * mat_B[86][1] +
                mat_A[26][3] * mat_B[94][1] +
                mat_A[27][0] * mat_B[102][1] +
                mat_A[27][1] * mat_B[110][1] +
                mat_A[27][2] * mat_B[118][1] +
                mat_A[27][3] * mat_B[126][1] +
                mat_A[28][0] * mat_B[134][1] +
                mat_A[28][1] * mat_B[142][1] +
                mat_A[28][2] * mat_B[150][1] +
                mat_A[28][3] * mat_B[158][1] +
                mat_A[29][0] * mat_B[166][1] +
                mat_A[29][1] * mat_B[174][1] +
                mat_A[29][2] * mat_B[182][1] +
                mat_A[29][3] * mat_B[190][1] +
                mat_A[30][0] * mat_B[198][1] +
                mat_A[30][1] * mat_B[206][1] +
                mat_A[30][2] * mat_B[214][1] +
                mat_A[30][3] * mat_B[222][1] +
                mat_A[31][0] * mat_B[230][1] +
                mat_A[31][1] * mat_B[238][1] +
                mat_A[31][2] * mat_B[246][1] +
                mat_A[31][3] * mat_B[254][1];
    mat_C[30][2] <=
                mat_A[24][0] * mat_B[6][2] +
                mat_A[24][1] * mat_B[14][2] +
                mat_A[24][2] * mat_B[22][2] +
                mat_A[24][3] * mat_B[30][2] +
                mat_A[25][0] * mat_B[38][2] +
                mat_A[25][1] * mat_B[46][2] +
                mat_A[25][2] * mat_B[54][2] +
                mat_A[25][3] * mat_B[62][2] +
                mat_A[26][0] * mat_B[70][2] +
                mat_A[26][1] * mat_B[78][2] +
                mat_A[26][2] * mat_B[86][2] +
                mat_A[26][3] * mat_B[94][2] +
                mat_A[27][0] * mat_B[102][2] +
                mat_A[27][1] * mat_B[110][2] +
                mat_A[27][2] * mat_B[118][2] +
                mat_A[27][3] * mat_B[126][2] +
                mat_A[28][0] * mat_B[134][2] +
                mat_A[28][1] * mat_B[142][2] +
                mat_A[28][2] * mat_B[150][2] +
                mat_A[28][3] * mat_B[158][2] +
                mat_A[29][0] * mat_B[166][2] +
                mat_A[29][1] * mat_B[174][2] +
                mat_A[29][2] * mat_B[182][2] +
                mat_A[29][3] * mat_B[190][2] +
                mat_A[30][0] * mat_B[198][2] +
                mat_A[30][1] * mat_B[206][2] +
                mat_A[30][2] * mat_B[214][2] +
                mat_A[30][3] * mat_B[222][2] +
                mat_A[31][0] * mat_B[230][2] +
                mat_A[31][1] * mat_B[238][2] +
                mat_A[31][2] * mat_B[246][2] +
                mat_A[31][3] * mat_B[254][2];
    mat_C[30][3] <=
                mat_A[24][0] * mat_B[6][3] +
                mat_A[24][1] * mat_B[14][3] +
                mat_A[24][2] * mat_B[22][3] +
                mat_A[24][3] * mat_B[30][3] +
                mat_A[25][0] * mat_B[38][3] +
                mat_A[25][1] * mat_B[46][3] +
                mat_A[25][2] * mat_B[54][3] +
                mat_A[25][3] * mat_B[62][3] +
                mat_A[26][0] * mat_B[70][3] +
                mat_A[26][1] * mat_B[78][3] +
                mat_A[26][2] * mat_B[86][3] +
                mat_A[26][3] * mat_B[94][3] +
                mat_A[27][0] * mat_B[102][3] +
                mat_A[27][1] * mat_B[110][3] +
                mat_A[27][2] * mat_B[118][3] +
                mat_A[27][3] * mat_B[126][3] +
                mat_A[28][0] * mat_B[134][3] +
                mat_A[28][1] * mat_B[142][3] +
                mat_A[28][2] * mat_B[150][3] +
                mat_A[28][3] * mat_B[158][3] +
                mat_A[29][0] * mat_B[166][3] +
                mat_A[29][1] * mat_B[174][3] +
                mat_A[29][2] * mat_B[182][3] +
                mat_A[29][3] * mat_B[190][3] +
                mat_A[30][0] * mat_B[198][3] +
                mat_A[30][1] * mat_B[206][3] +
                mat_A[30][2] * mat_B[214][3] +
                mat_A[30][3] * mat_B[222][3] +
                mat_A[31][0] * mat_B[230][3] +
                mat_A[31][1] * mat_B[238][3] +
                mat_A[31][2] * mat_B[246][3] +
                mat_A[31][3] * mat_B[254][3];
    mat_C[31][0] <=
                mat_A[24][0] * mat_B[7][0] +
                mat_A[24][1] * mat_B[15][0] +
                mat_A[24][2] * mat_B[23][0] +
                mat_A[24][3] * mat_B[31][0] +
                mat_A[25][0] * mat_B[39][0] +
                mat_A[25][1] * mat_B[47][0] +
                mat_A[25][2] * mat_B[55][0] +
                mat_A[25][3] * mat_B[63][0] +
                mat_A[26][0] * mat_B[71][0] +
                mat_A[26][1] * mat_B[79][0] +
                mat_A[26][2] * mat_B[87][0] +
                mat_A[26][3] * mat_B[95][0] +
                mat_A[27][0] * mat_B[103][0] +
                mat_A[27][1] * mat_B[111][0] +
                mat_A[27][2] * mat_B[119][0] +
                mat_A[27][3] * mat_B[127][0] +
                mat_A[28][0] * mat_B[135][0] +
                mat_A[28][1] * mat_B[143][0] +
                mat_A[28][2] * mat_B[151][0] +
                mat_A[28][3] * mat_B[159][0] +
                mat_A[29][0] * mat_B[167][0] +
                mat_A[29][1] * mat_B[175][0] +
                mat_A[29][2] * mat_B[183][0] +
                mat_A[29][3] * mat_B[191][0] +
                mat_A[30][0] * mat_B[199][0] +
                mat_A[30][1] * mat_B[207][0] +
                mat_A[30][2] * mat_B[215][0] +
                mat_A[30][3] * mat_B[223][0] +
                mat_A[31][0] * mat_B[231][0] +
                mat_A[31][1] * mat_B[239][0] +
                mat_A[31][2] * mat_B[247][0] +
                mat_A[31][3] * mat_B[255][0];
    mat_C[31][1] <=
                mat_A[24][0] * mat_B[7][1] +
                mat_A[24][1] * mat_B[15][1] +
                mat_A[24][2] * mat_B[23][1] +
                mat_A[24][3] * mat_B[31][1] +
                mat_A[25][0] * mat_B[39][1] +
                mat_A[25][1] * mat_B[47][1] +
                mat_A[25][2] * mat_B[55][1] +
                mat_A[25][3] * mat_B[63][1] +
                mat_A[26][0] * mat_B[71][1] +
                mat_A[26][1] * mat_B[79][1] +
                mat_A[26][2] * mat_B[87][1] +
                mat_A[26][3] * mat_B[95][1] +
                mat_A[27][0] * mat_B[103][1] +
                mat_A[27][1] * mat_B[111][1] +
                mat_A[27][2] * mat_B[119][1] +
                mat_A[27][3] * mat_B[127][1] +
                mat_A[28][0] * mat_B[135][1] +
                mat_A[28][1] * mat_B[143][1] +
                mat_A[28][2] * mat_B[151][1] +
                mat_A[28][3] * mat_B[159][1] +
                mat_A[29][0] * mat_B[167][1] +
                mat_A[29][1] * mat_B[175][1] +
                mat_A[29][2] * mat_B[183][1] +
                mat_A[29][3] * mat_B[191][1] +
                mat_A[30][0] * mat_B[199][1] +
                mat_A[30][1] * mat_B[207][1] +
                mat_A[30][2] * mat_B[215][1] +
                mat_A[30][3] * mat_B[223][1] +
                mat_A[31][0] * mat_B[231][1] +
                mat_A[31][1] * mat_B[239][1] +
                mat_A[31][2] * mat_B[247][1] +
                mat_A[31][3] * mat_B[255][1];
    mat_C[31][2] <=
                mat_A[24][0] * mat_B[7][2] +
                mat_A[24][1] * mat_B[15][2] +
                mat_A[24][2] * mat_B[23][2] +
                mat_A[24][3] * mat_B[31][2] +
                mat_A[25][0] * mat_B[39][2] +
                mat_A[25][1] * mat_B[47][2] +
                mat_A[25][2] * mat_B[55][2] +
                mat_A[25][3] * mat_B[63][2] +
                mat_A[26][0] * mat_B[71][2] +
                mat_A[26][1] * mat_B[79][2] +
                mat_A[26][2] * mat_B[87][2] +
                mat_A[26][3] * mat_B[95][2] +
                mat_A[27][0] * mat_B[103][2] +
                mat_A[27][1] * mat_B[111][2] +
                mat_A[27][2] * mat_B[119][2] +
                mat_A[27][3] * mat_B[127][2] +
                mat_A[28][0] * mat_B[135][2] +
                mat_A[28][1] * mat_B[143][2] +
                mat_A[28][2] * mat_B[151][2] +
                mat_A[28][3] * mat_B[159][2] +
                mat_A[29][0] * mat_B[167][2] +
                mat_A[29][1] * mat_B[175][2] +
                mat_A[29][2] * mat_B[183][2] +
                mat_A[29][3] * mat_B[191][2] +
                mat_A[30][0] * mat_B[199][2] +
                mat_A[30][1] * mat_B[207][2] +
                mat_A[30][2] * mat_B[215][2] +
                mat_A[30][3] * mat_B[223][2] +
                mat_A[31][0] * mat_B[231][2] +
                mat_A[31][1] * mat_B[239][2] +
                mat_A[31][2] * mat_B[247][2] +
                mat_A[31][3] * mat_B[255][2];
    mat_C[31][3] <=
                mat_A[24][0] * mat_B[7][3] +
                mat_A[24][1] * mat_B[15][3] +
                mat_A[24][2] * mat_B[23][3] +
                mat_A[24][3] * mat_B[31][3] +
                mat_A[25][0] * mat_B[39][3] +
                mat_A[25][1] * mat_B[47][3] +
                mat_A[25][2] * mat_B[55][3] +
                mat_A[25][3] * mat_B[63][3] +
                mat_A[26][0] * mat_B[71][3] +
                mat_A[26][1] * mat_B[79][3] +
                mat_A[26][2] * mat_B[87][3] +
                mat_A[26][3] * mat_B[95][3] +
                mat_A[27][0] * mat_B[103][3] +
                mat_A[27][1] * mat_B[111][3] +
                mat_A[27][2] * mat_B[119][3] +
                mat_A[27][3] * mat_B[127][3] +
                mat_A[28][0] * mat_B[135][3] +
                mat_A[28][1] * mat_B[143][3] +
                mat_A[28][2] * mat_B[151][3] +
                mat_A[28][3] * mat_B[159][3] +
                mat_A[29][0] * mat_B[167][3] +
                mat_A[29][1] * mat_B[175][3] +
                mat_A[29][2] * mat_B[183][3] +
                mat_A[29][3] * mat_B[191][3] +
                mat_A[30][0] * mat_B[199][3] +
                mat_A[30][1] * mat_B[207][3] +
                mat_A[30][2] * mat_B[215][3] +
                mat_A[30][3] * mat_B[223][3] +
                mat_A[31][0] * mat_B[231][3] +
                mat_A[31][1] * mat_B[239][3] +
                mat_A[31][2] * mat_B[247][3] +
                mat_A[31][3] * mat_B[255][3];
    mat_C[32][0] <=
                mat_A[32][0] * mat_B[0][0] +
                mat_A[32][1] * mat_B[8][0] +
                mat_A[32][2] * mat_B[16][0] +
                mat_A[32][3] * mat_B[24][0] +
                mat_A[33][0] * mat_B[32][0] +
                mat_A[33][1] * mat_B[40][0] +
                mat_A[33][2] * mat_B[48][0] +
                mat_A[33][3] * mat_B[56][0] +
                mat_A[34][0] * mat_B[64][0] +
                mat_A[34][1] * mat_B[72][0] +
                mat_A[34][2] * mat_B[80][0] +
                mat_A[34][3] * mat_B[88][0] +
                mat_A[35][0] * mat_B[96][0] +
                mat_A[35][1] * mat_B[104][0] +
                mat_A[35][2] * mat_B[112][0] +
                mat_A[35][3] * mat_B[120][0] +
                mat_A[36][0] * mat_B[128][0] +
                mat_A[36][1] * mat_B[136][0] +
                mat_A[36][2] * mat_B[144][0] +
                mat_A[36][3] * mat_B[152][0] +
                mat_A[37][0] * mat_B[160][0] +
                mat_A[37][1] * mat_B[168][0] +
                mat_A[37][2] * mat_B[176][0] +
                mat_A[37][3] * mat_B[184][0] +
                mat_A[38][0] * mat_B[192][0] +
                mat_A[38][1] * mat_B[200][0] +
                mat_A[38][2] * mat_B[208][0] +
                mat_A[38][3] * mat_B[216][0] +
                mat_A[39][0] * mat_B[224][0] +
                mat_A[39][1] * mat_B[232][0] +
                mat_A[39][2] * mat_B[240][0] +
                mat_A[39][3] * mat_B[248][0];
    mat_C[32][1] <=
                mat_A[32][0] * mat_B[0][1] +
                mat_A[32][1] * mat_B[8][1] +
                mat_A[32][2] * mat_B[16][1] +
                mat_A[32][3] * mat_B[24][1] +
                mat_A[33][0] * mat_B[32][1] +
                mat_A[33][1] * mat_B[40][1] +
                mat_A[33][2] * mat_B[48][1] +
                mat_A[33][3] * mat_B[56][1] +
                mat_A[34][0] * mat_B[64][1] +
                mat_A[34][1] * mat_B[72][1] +
                mat_A[34][2] * mat_B[80][1] +
                mat_A[34][3] * mat_B[88][1] +
                mat_A[35][0] * mat_B[96][1] +
                mat_A[35][1] * mat_B[104][1] +
                mat_A[35][2] * mat_B[112][1] +
                mat_A[35][3] * mat_B[120][1] +
                mat_A[36][0] * mat_B[128][1] +
                mat_A[36][1] * mat_B[136][1] +
                mat_A[36][2] * mat_B[144][1] +
                mat_A[36][3] * mat_B[152][1] +
                mat_A[37][0] * mat_B[160][1] +
                mat_A[37][1] * mat_B[168][1] +
                mat_A[37][2] * mat_B[176][1] +
                mat_A[37][3] * mat_B[184][1] +
                mat_A[38][0] * mat_B[192][1] +
                mat_A[38][1] * mat_B[200][1] +
                mat_A[38][2] * mat_B[208][1] +
                mat_A[38][3] * mat_B[216][1] +
                mat_A[39][0] * mat_B[224][1] +
                mat_A[39][1] * mat_B[232][1] +
                mat_A[39][2] * mat_B[240][1] +
                mat_A[39][3] * mat_B[248][1];
    mat_C[32][2] <=
                mat_A[32][0] * mat_B[0][2] +
                mat_A[32][1] * mat_B[8][2] +
                mat_A[32][2] * mat_B[16][2] +
                mat_A[32][3] * mat_B[24][2] +
                mat_A[33][0] * mat_B[32][2] +
                mat_A[33][1] * mat_B[40][2] +
                mat_A[33][2] * mat_B[48][2] +
                mat_A[33][3] * mat_B[56][2] +
                mat_A[34][0] * mat_B[64][2] +
                mat_A[34][1] * mat_B[72][2] +
                mat_A[34][2] * mat_B[80][2] +
                mat_A[34][3] * mat_B[88][2] +
                mat_A[35][0] * mat_B[96][2] +
                mat_A[35][1] * mat_B[104][2] +
                mat_A[35][2] * mat_B[112][2] +
                mat_A[35][3] * mat_B[120][2] +
                mat_A[36][0] * mat_B[128][2] +
                mat_A[36][1] * mat_B[136][2] +
                mat_A[36][2] * mat_B[144][2] +
                mat_A[36][3] * mat_B[152][2] +
                mat_A[37][0] * mat_B[160][2] +
                mat_A[37][1] * mat_B[168][2] +
                mat_A[37][2] * mat_B[176][2] +
                mat_A[37][3] * mat_B[184][2] +
                mat_A[38][0] * mat_B[192][2] +
                mat_A[38][1] * mat_B[200][2] +
                mat_A[38][2] * mat_B[208][2] +
                mat_A[38][3] * mat_B[216][2] +
                mat_A[39][0] * mat_B[224][2] +
                mat_A[39][1] * mat_B[232][2] +
                mat_A[39][2] * mat_B[240][2] +
                mat_A[39][3] * mat_B[248][2];
    mat_C[32][3] <=
                mat_A[32][0] * mat_B[0][3] +
                mat_A[32][1] * mat_B[8][3] +
                mat_A[32][2] * mat_B[16][3] +
                mat_A[32][3] * mat_B[24][3] +
                mat_A[33][0] * mat_B[32][3] +
                mat_A[33][1] * mat_B[40][3] +
                mat_A[33][2] * mat_B[48][3] +
                mat_A[33][3] * mat_B[56][3] +
                mat_A[34][0] * mat_B[64][3] +
                mat_A[34][1] * mat_B[72][3] +
                mat_A[34][2] * mat_B[80][3] +
                mat_A[34][3] * mat_B[88][3] +
                mat_A[35][0] * mat_B[96][3] +
                mat_A[35][1] * mat_B[104][3] +
                mat_A[35][2] * mat_B[112][3] +
                mat_A[35][3] * mat_B[120][3] +
                mat_A[36][0] * mat_B[128][3] +
                mat_A[36][1] * mat_B[136][3] +
                mat_A[36][2] * mat_B[144][3] +
                mat_A[36][3] * mat_B[152][3] +
                mat_A[37][0] * mat_B[160][3] +
                mat_A[37][1] * mat_B[168][3] +
                mat_A[37][2] * mat_B[176][3] +
                mat_A[37][3] * mat_B[184][3] +
                mat_A[38][0] * mat_B[192][3] +
                mat_A[38][1] * mat_B[200][3] +
                mat_A[38][2] * mat_B[208][3] +
                mat_A[38][3] * mat_B[216][3] +
                mat_A[39][0] * mat_B[224][3] +
                mat_A[39][1] * mat_B[232][3] +
                mat_A[39][2] * mat_B[240][3] +
                mat_A[39][3] * mat_B[248][3];
    mat_C[33][0] <=
                mat_A[32][0] * mat_B[1][0] +
                mat_A[32][1] * mat_B[9][0] +
                mat_A[32][2] * mat_B[17][0] +
                mat_A[32][3] * mat_B[25][0] +
                mat_A[33][0] * mat_B[33][0] +
                mat_A[33][1] * mat_B[41][0] +
                mat_A[33][2] * mat_B[49][0] +
                mat_A[33][3] * mat_B[57][0] +
                mat_A[34][0] * mat_B[65][0] +
                mat_A[34][1] * mat_B[73][0] +
                mat_A[34][2] * mat_B[81][0] +
                mat_A[34][3] * mat_B[89][0] +
                mat_A[35][0] * mat_B[97][0] +
                mat_A[35][1] * mat_B[105][0] +
                mat_A[35][2] * mat_B[113][0] +
                mat_A[35][3] * mat_B[121][0] +
                mat_A[36][0] * mat_B[129][0] +
                mat_A[36][1] * mat_B[137][0] +
                mat_A[36][2] * mat_B[145][0] +
                mat_A[36][3] * mat_B[153][0] +
                mat_A[37][0] * mat_B[161][0] +
                mat_A[37][1] * mat_B[169][0] +
                mat_A[37][2] * mat_B[177][0] +
                mat_A[37][3] * mat_B[185][0] +
                mat_A[38][0] * mat_B[193][0] +
                mat_A[38][1] * mat_B[201][0] +
                mat_A[38][2] * mat_B[209][0] +
                mat_A[38][3] * mat_B[217][0] +
                mat_A[39][0] * mat_B[225][0] +
                mat_A[39][1] * mat_B[233][0] +
                mat_A[39][2] * mat_B[241][0] +
                mat_A[39][3] * mat_B[249][0];
    mat_C[33][1] <=
                mat_A[32][0] * mat_B[1][1] +
                mat_A[32][1] * mat_B[9][1] +
                mat_A[32][2] * mat_B[17][1] +
                mat_A[32][3] * mat_B[25][1] +
                mat_A[33][0] * mat_B[33][1] +
                mat_A[33][1] * mat_B[41][1] +
                mat_A[33][2] * mat_B[49][1] +
                mat_A[33][3] * mat_B[57][1] +
                mat_A[34][0] * mat_B[65][1] +
                mat_A[34][1] * mat_B[73][1] +
                mat_A[34][2] * mat_B[81][1] +
                mat_A[34][3] * mat_B[89][1] +
                mat_A[35][0] * mat_B[97][1] +
                mat_A[35][1] * mat_B[105][1] +
                mat_A[35][2] * mat_B[113][1] +
                mat_A[35][3] * mat_B[121][1] +
                mat_A[36][0] * mat_B[129][1] +
                mat_A[36][1] * mat_B[137][1] +
                mat_A[36][2] * mat_B[145][1] +
                mat_A[36][3] * mat_B[153][1] +
                mat_A[37][0] * mat_B[161][1] +
                mat_A[37][1] * mat_B[169][1] +
                mat_A[37][2] * mat_B[177][1] +
                mat_A[37][3] * mat_B[185][1] +
                mat_A[38][0] * mat_B[193][1] +
                mat_A[38][1] * mat_B[201][1] +
                mat_A[38][2] * mat_B[209][1] +
                mat_A[38][3] * mat_B[217][1] +
                mat_A[39][0] * mat_B[225][1] +
                mat_A[39][1] * mat_B[233][1] +
                mat_A[39][2] * mat_B[241][1] +
                mat_A[39][3] * mat_B[249][1];
    mat_C[33][2] <=
                mat_A[32][0] * mat_B[1][2] +
                mat_A[32][1] * mat_B[9][2] +
                mat_A[32][2] * mat_B[17][2] +
                mat_A[32][3] * mat_B[25][2] +
                mat_A[33][0] * mat_B[33][2] +
                mat_A[33][1] * mat_B[41][2] +
                mat_A[33][2] * mat_B[49][2] +
                mat_A[33][3] * mat_B[57][2] +
                mat_A[34][0] * mat_B[65][2] +
                mat_A[34][1] * mat_B[73][2] +
                mat_A[34][2] * mat_B[81][2] +
                mat_A[34][3] * mat_B[89][2] +
                mat_A[35][0] * mat_B[97][2] +
                mat_A[35][1] * mat_B[105][2] +
                mat_A[35][2] * mat_B[113][2] +
                mat_A[35][3] * mat_B[121][2] +
                mat_A[36][0] * mat_B[129][2] +
                mat_A[36][1] * mat_B[137][2] +
                mat_A[36][2] * mat_B[145][2] +
                mat_A[36][3] * mat_B[153][2] +
                mat_A[37][0] * mat_B[161][2] +
                mat_A[37][1] * mat_B[169][2] +
                mat_A[37][2] * mat_B[177][2] +
                mat_A[37][3] * mat_B[185][2] +
                mat_A[38][0] * mat_B[193][2] +
                mat_A[38][1] * mat_B[201][2] +
                mat_A[38][2] * mat_B[209][2] +
                mat_A[38][3] * mat_B[217][2] +
                mat_A[39][0] * mat_B[225][2] +
                mat_A[39][1] * mat_B[233][2] +
                mat_A[39][2] * mat_B[241][2] +
                mat_A[39][3] * mat_B[249][2];
    mat_C[33][3] <=
                mat_A[32][0] * mat_B[1][3] +
                mat_A[32][1] * mat_B[9][3] +
                mat_A[32][2] * mat_B[17][3] +
                mat_A[32][3] * mat_B[25][3] +
                mat_A[33][0] * mat_B[33][3] +
                mat_A[33][1] * mat_B[41][3] +
                mat_A[33][2] * mat_B[49][3] +
                mat_A[33][3] * mat_B[57][3] +
                mat_A[34][0] * mat_B[65][3] +
                mat_A[34][1] * mat_B[73][3] +
                mat_A[34][2] * mat_B[81][3] +
                mat_A[34][3] * mat_B[89][3] +
                mat_A[35][0] * mat_B[97][3] +
                mat_A[35][1] * mat_B[105][3] +
                mat_A[35][2] * mat_B[113][3] +
                mat_A[35][3] * mat_B[121][3] +
                mat_A[36][0] * mat_B[129][3] +
                mat_A[36][1] * mat_B[137][3] +
                mat_A[36][2] * mat_B[145][3] +
                mat_A[36][3] * mat_B[153][3] +
                mat_A[37][0] * mat_B[161][3] +
                mat_A[37][1] * mat_B[169][3] +
                mat_A[37][2] * mat_B[177][3] +
                mat_A[37][3] * mat_B[185][3] +
                mat_A[38][0] * mat_B[193][3] +
                mat_A[38][1] * mat_B[201][3] +
                mat_A[38][2] * mat_B[209][3] +
                mat_A[38][3] * mat_B[217][3] +
                mat_A[39][0] * mat_B[225][3] +
                mat_A[39][1] * mat_B[233][3] +
                mat_A[39][2] * mat_B[241][3] +
                mat_A[39][3] * mat_B[249][3];
    mat_C[34][0] <=
                mat_A[32][0] * mat_B[2][0] +
                mat_A[32][1] * mat_B[10][0] +
                mat_A[32][2] * mat_B[18][0] +
                mat_A[32][3] * mat_B[26][0] +
                mat_A[33][0] * mat_B[34][0] +
                mat_A[33][1] * mat_B[42][0] +
                mat_A[33][2] * mat_B[50][0] +
                mat_A[33][3] * mat_B[58][0] +
                mat_A[34][0] * mat_B[66][0] +
                mat_A[34][1] * mat_B[74][0] +
                mat_A[34][2] * mat_B[82][0] +
                mat_A[34][3] * mat_B[90][0] +
                mat_A[35][0] * mat_B[98][0] +
                mat_A[35][1] * mat_B[106][0] +
                mat_A[35][2] * mat_B[114][0] +
                mat_A[35][3] * mat_B[122][0] +
                mat_A[36][0] * mat_B[130][0] +
                mat_A[36][1] * mat_B[138][0] +
                mat_A[36][2] * mat_B[146][0] +
                mat_A[36][3] * mat_B[154][0] +
                mat_A[37][0] * mat_B[162][0] +
                mat_A[37][1] * mat_B[170][0] +
                mat_A[37][2] * mat_B[178][0] +
                mat_A[37][3] * mat_B[186][0] +
                mat_A[38][0] * mat_B[194][0] +
                mat_A[38][1] * mat_B[202][0] +
                mat_A[38][2] * mat_B[210][0] +
                mat_A[38][3] * mat_B[218][0] +
                mat_A[39][0] * mat_B[226][0] +
                mat_A[39][1] * mat_B[234][0] +
                mat_A[39][2] * mat_B[242][0] +
                mat_A[39][3] * mat_B[250][0];
    mat_C[34][1] <=
                mat_A[32][0] * mat_B[2][1] +
                mat_A[32][1] * mat_B[10][1] +
                mat_A[32][2] * mat_B[18][1] +
                mat_A[32][3] * mat_B[26][1] +
                mat_A[33][0] * mat_B[34][1] +
                mat_A[33][1] * mat_B[42][1] +
                mat_A[33][2] * mat_B[50][1] +
                mat_A[33][3] * mat_B[58][1] +
                mat_A[34][0] * mat_B[66][1] +
                mat_A[34][1] * mat_B[74][1] +
                mat_A[34][2] * mat_B[82][1] +
                mat_A[34][3] * mat_B[90][1] +
                mat_A[35][0] * mat_B[98][1] +
                mat_A[35][1] * mat_B[106][1] +
                mat_A[35][2] * mat_B[114][1] +
                mat_A[35][3] * mat_B[122][1] +
                mat_A[36][0] * mat_B[130][1] +
                mat_A[36][1] * mat_B[138][1] +
                mat_A[36][2] * mat_B[146][1] +
                mat_A[36][3] * mat_B[154][1] +
                mat_A[37][0] * mat_B[162][1] +
                mat_A[37][1] * mat_B[170][1] +
                mat_A[37][2] * mat_B[178][1] +
                mat_A[37][3] * mat_B[186][1] +
                mat_A[38][0] * mat_B[194][1] +
                mat_A[38][1] * mat_B[202][1] +
                mat_A[38][2] * mat_B[210][1] +
                mat_A[38][3] * mat_B[218][1] +
                mat_A[39][0] * mat_B[226][1] +
                mat_A[39][1] * mat_B[234][1] +
                mat_A[39][2] * mat_B[242][1] +
                mat_A[39][3] * mat_B[250][1];
    mat_C[34][2] <=
                mat_A[32][0] * mat_B[2][2] +
                mat_A[32][1] * mat_B[10][2] +
                mat_A[32][2] * mat_B[18][2] +
                mat_A[32][3] * mat_B[26][2] +
                mat_A[33][0] * mat_B[34][2] +
                mat_A[33][1] * mat_B[42][2] +
                mat_A[33][2] * mat_B[50][2] +
                mat_A[33][3] * mat_B[58][2] +
                mat_A[34][0] * mat_B[66][2] +
                mat_A[34][1] * mat_B[74][2] +
                mat_A[34][2] * mat_B[82][2] +
                mat_A[34][3] * mat_B[90][2] +
                mat_A[35][0] * mat_B[98][2] +
                mat_A[35][1] * mat_B[106][2] +
                mat_A[35][2] * mat_B[114][2] +
                mat_A[35][3] * mat_B[122][2] +
                mat_A[36][0] * mat_B[130][2] +
                mat_A[36][1] * mat_B[138][2] +
                mat_A[36][2] * mat_B[146][2] +
                mat_A[36][3] * mat_B[154][2] +
                mat_A[37][0] * mat_B[162][2] +
                mat_A[37][1] * mat_B[170][2] +
                mat_A[37][2] * mat_B[178][2] +
                mat_A[37][3] * mat_B[186][2] +
                mat_A[38][0] * mat_B[194][2] +
                mat_A[38][1] * mat_B[202][2] +
                mat_A[38][2] * mat_B[210][2] +
                mat_A[38][3] * mat_B[218][2] +
                mat_A[39][0] * mat_B[226][2] +
                mat_A[39][1] * mat_B[234][2] +
                mat_A[39][2] * mat_B[242][2] +
                mat_A[39][3] * mat_B[250][2];
    mat_C[34][3] <=
                mat_A[32][0] * mat_B[2][3] +
                mat_A[32][1] * mat_B[10][3] +
                mat_A[32][2] * mat_B[18][3] +
                mat_A[32][3] * mat_B[26][3] +
                mat_A[33][0] * mat_B[34][3] +
                mat_A[33][1] * mat_B[42][3] +
                mat_A[33][2] * mat_B[50][3] +
                mat_A[33][3] * mat_B[58][3] +
                mat_A[34][0] * mat_B[66][3] +
                mat_A[34][1] * mat_B[74][3] +
                mat_A[34][2] * mat_B[82][3] +
                mat_A[34][3] * mat_B[90][3] +
                mat_A[35][0] * mat_B[98][3] +
                mat_A[35][1] * mat_B[106][3] +
                mat_A[35][2] * mat_B[114][3] +
                mat_A[35][3] * mat_B[122][3] +
                mat_A[36][0] * mat_B[130][3] +
                mat_A[36][1] * mat_B[138][3] +
                mat_A[36][2] * mat_B[146][3] +
                mat_A[36][3] * mat_B[154][3] +
                mat_A[37][0] * mat_B[162][3] +
                mat_A[37][1] * mat_B[170][3] +
                mat_A[37][2] * mat_B[178][3] +
                mat_A[37][3] * mat_B[186][3] +
                mat_A[38][0] * mat_B[194][3] +
                mat_A[38][1] * mat_B[202][3] +
                mat_A[38][2] * mat_B[210][3] +
                mat_A[38][3] * mat_B[218][3] +
                mat_A[39][0] * mat_B[226][3] +
                mat_A[39][1] * mat_B[234][3] +
                mat_A[39][2] * mat_B[242][3] +
                mat_A[39][3] * mat_B[250][3];
    mat_C[35][0] <=
                mat_A[32][0] * mat_B[3][0] +
                mat_A[32][1] * mat_B[11][0] +
                mat_A[32][2] * mat_B[19][0] +
                mat_A[32][3] * mat_B[27][0] +
                mat_A[33][0] * mat_B[35][0] +
                mat_A[33][1] * mat_B[43][0] +
                mat_A[33][2] * mat_B[51][0] +
                mat_A[33][3] * mat_B[59][0] +
                mat_A[34][0] * mat_B[67][0] +
                mat_A[34][1] * mat_B[75][0] +
                mat_A[34][2] * mat_B[83][0] +
                mat_A[34][3] * mat_B[91][0] +
                mat_A[35][0] * mat_B[99][0] +
                mat_A[35][1] * mat_B[107][0] +
                mat_A[35][2] * mat_B[115][0] +
                mat_A[35][3] * mat_B[123][0] +
                mat_A[36][0] * mat_B[131][0] +
                mat_A[36][1] * mat_B[139][0] +
                mat_A[36][2] * mat_B[147][0] +
                mat_A[36][3] * mat_B[155][0] +
                mat_A[37][0] * mat_B[163][0] +
                mat_A[37][1] * mat_B[171][0] +
                mat_A[37][2] * mat_B[179][0] +
                mat_A[37][3] * mat_B[187][0] +
                mat_A[38][0] * mat_B[195][0] +
                mat_A[38][1] * mat_B[203][0] +
                mat_A[38][2] * mat_B[211][0] +
                mat_A[38][3] * mat_B[219][0] +
                mat_A[39][0] * mat_B[227][0] +
                mat_A[39][1] * mat_B[235][0] +
                mat_A[39][2] * mat_B[243][0] +
                mat_A[39][3] * mat_B[251][0];
    mat_C[35][1] <=
                mat_A[32][0] * mat_B[3][1] +
                mat_A[32][1] * mat_B[11][1] +
                mat_A[32][2] * mat_B[19][1] +
                mat_A[32][3] * mat_B[27][1] +
                mat_A[33][0] * mat_B[35][1] +
                mat_A[33][1] * mat_B[43][1] +
                mat_A[33][2] * mat_B[51][1] +
                mat_A[33][3] * mat_B[59][1] +
                mat_A[34][0] * mat_B[67][1] +
                mat_A[34][1] * mat_B[75][1] +
                mat_A[34][2] * mat_B[83][1] +
                mat_A[34][3] * mat_B[91][1] +
                mat_A[35][0] * mat_B[99][1] +
                mat_A[35][1] * mat_B[107][1] +
                mat_A[35][2] * mat_B[115][1] +
                mat_A[35][3] * mat_B[123][1] +
                mat_A[36][0] * mat_B[131][1] +
                mat_A[36][1] * mat_B[139][1] +
                mat_A[36][2] * mat_B[147][1] +
                mat_A[36][3] * mat_B[155][1] +
                mat_A[37][0] * mat_B[163][1] +
                mat_A[37][1] * mat_B[171][1] +
                mat_A[37][2] * mat_B[179][1] +
                mat_A[37][3] * mat_B[187][1] +
                mat_A[38][0] * mat_B[195][1] +
                mat_A[38][1] * mat_B[203][1] +
                mat_A[38][2] * mat_B[211][1] +
                mat_A[38][3] * mat_B[219][1] +
                mat_A[39][0] * mat_B[227][1] +
                mat_A[39][1] * mat_B[235][1] +
                mat_A[39][2] * mat_B[243][1] +
                mat_A[39][3] * mat_B[251][1];
    mat_C[35][2] <=
                mat_A[32][0] * mat_B[3][2] +
                mat_A[32][1] * mat_B[11][2] +
                mat_A[32][2] * mat_B[19][2] +
                mat_A[32][3] * mat_B[27][2] +
                mat_A[33][0] * mat_B[35][2] +
                mat_A[33][1] * mat_B[43][2] +
                mat_A[33][2] * mat_B[51][2] +
                mat_A[33][3] * mat_B[59][2] +
                mat_A[34][0] * mat_B[67][2] +
                mat_A[34][1] * mat_B[75][2] +
                mat_A[34][2] * mat_B[83][2] +
                mat_A[34][3] * mat_B[91][2] +
                mat_A[35][0] * mat_B[99][2] +
                mat_A[35][1] * mat_B[107][2] +
                mat_A[35][2] * mat_B[115][2] +
                mat_A[35][3] * mat_B[123][2] +
                mat_A[36][0] * mat_B[131][2] +
                mat_A[36][1] * mat_B[139][2] +
                mat_A[36][2] * mat_B[147][2] +
                mat_A[36][3] * mat_B[155][2] +
                mat_A[37][0] * mat_B[163][2] +
                mat_A[37][1] * mat_B[171][2] +
                mat_A[37][2] * mat_B[179][2] +
                mat_A[37][3] * mat_B[187][2] +
                mat_A[38][0] * mat_B[195][2] +
                mat_A[38][1] * mat_B[203][2] +
                mat_A[38][2] * mat_B[211][2] +
                mat_A[38][3] * mat_B[219][2] +
                mat_A[39][0] * mat_B[227][2] +
                mat_A[39][1] * mat_B[235][2] +
                mat_A[39][2] * mat_B[243][2] +
                mat_A[39][3] * mat_B[251][2];
    mat_C[35][3] <=
                mat_A[32][0] * mat_B[3][3] +
                mat_A[32][1] * mat_B[11][3] +
                mat_A[32][2] * mat_B[19][3] +
                mat_A[32][3] * mat_B[27][3] +
                mat_A[33][0] * mat_B[35][3] +
                mat_A[33][1] * mat_B[43][3] +
                mat_A[33][2] * mat_B[51][3] +
                mat_A[33][3] * mat_B[59][3] +
                mat_A[34][0] * mat_B[67][3] +
                mat_A[34][1] * mat_B[75][3] +
                mat_A[34][2] * mat_B[83][3] +
                mat_A[34][3] * mat_B[91][3] +
                mat_A[35][0] * mat_B[99][3] +
                mat_A[35][1] * mat_B[107][3] +
                mat_A[35][2] * mat_B[115][3] +
                mat_A[35][3] * mat_B[123][3] +
                mat_A[36][0] * mat_B[131][3] +
                mat_A[36][1] * mat_B[139][3] +
                mat_A[36][2] * mat_B[147][3] +
                mat_A[36][3] * mat_B[155][3] +
                mat_A[37][0] * mat_B[163][3] +
                mat_A[37][1] * mat_B[171][3] +
                mat_A[37][2] * mat_B[179][3] +
                mat_A[37][3] * mat_B[187][3] +
                mat_A[38][0] * mat_B[195][3] +
                mat_A[38][1] * mat_B[203][3] +
                mat_A[38][2] * mat_B[211][3] +
                mat_A[38][3] * mat_B[219][3] +
                mat_A[39][0] * mat_B[227][3] +
                mat_A[39][1] * mat_B[235][3] +
                mat_A[39][2] * mat_B[243][3] +
                mat_A[39][3] * mat_B[251][3];
    mat_C[36][0] <=
                mat_A[32][0] * mat_B[4][0] +
                mat_A[32][1] * mat_B[12][0] +
                mat_A[32][2] * mat_B[20][0] +
                mat_A[32][3] * mat_B[28][0] +
                mat_A[33][0] * mat_B[36][0] +
                mat_A[33][1] * mat_B[44][0] +
                mat_A[33][2] * mat_B[52][0] +
                mat_A[33][3] * mat_B[60][0] +
                mat_A[34][0] * mat_B[68][0] +
                mat_A[34][1] * mat_B[76][0] +
                mat_A[34][2] * mat_B[84][0] +
                mat_A[34][3] * mat_B[92][0] +
                mat_A[35][0] * mat_B[100][0] +
                mat_A[35][1] * mat_B[108][0] +
                mat_A[35][2] * mat_B[116][0] +
                mat_A[35][3] * mat_B[124][0] +
                mat_A[36][0] * mat_B[132][0] +
                mat_A[36][1] * mat_B[140][0] +
                mat_A[36][2] * mat_B[148][0] +
                mat_A[36][3] * mat_B[156][0] +
                mat_A[37][0] * mat_B[164][0] +
                mat_A[37][1] * mat_B[172][0] +
                mat_A[37][2] * mat_B[180][0] +
                mat_A[37][3] * mat_B[188][0] +
                mat_A[38][0] * mat_B[196][0] +
                mat_A[38][1] * mat_B[204][0] +
                mat_A[38][2] * mat_B[212][0] +
                mat_A[38][3] * mat_B[220][0] +
                mat_A[39][0] * mat_B[228][0] +
                mat_A[39][1] * mat_B[236][0] +
                mat_A[39][2] * mat_B[244][0] +
                mat_A[39][3] * mat_B[252][0];
    mat_C[36][1] <=
                mat_A[32][0] * mat_B[4][1] +
                mat_A[32][1] * mat_B[12][1] +
                mat_A[32][2] * mat_B[20][1] +
                mat_A[32][3] * mat_B[28][1] +
                mat_A[33][0] * mat_B[36][1] +
                mat_A[33][1] * mat_B[44][1] +
                mat_A[33][2] * mat_B[52][1] +
                mat_A[33][3] * mat_B[60][1] +
                mat_A[34][0] * mat_B[68][1] +
                mat_A[34][1] * mat_B[76][1] +
                mat_A[34][2] * mat_B[84][1] +
                mat_A[34][3] * mat_B[92][1] +
                mat_A[35][0] * mat_B[100][1] +
                mat_A[35][1] * mat_B[108][1] +
                mat_A[35][2] * mat_B[116][1] +
                mat_A[35][3] * mat_B[124][1] +
                mat_A[36][0] * mat_B[132][1] +
                mat_A[36][1] * mat_B[140][1] +
                mat_A[36][2] * mat_B[148][1] +
                mat_A[36][3] * mat_B[156][1] +
                mat_A[37][0] * mat_B[164][1] +
                mat_A[37][1] * mat_B[172][1] +
                mat_A[37][2] * mat_B[180][1] +
                mat_A[37][3] * mat_B[188][1] +
                mat_A[38][0] * mat_B[196][1] +
                mat_A[38][1] * mat_B[204][1] +
                mat_A[38][2] * mat_B[212][1] +
                mat_A[38][3] * mat_B[220][1] +
                mat_A[39][0] * mat_B[228][1] +
                mat_A[39][1] * mat_B[236][1] +
                mat_A[39][2] * mat_B[244][1] +
                mat_A[39][3] * mat_B[252][1];
    mat_C[36][2] <=
                mat_A[32][0] * mat_B[4][2] +
                mat_A[32][1] * mat_B[12][2] +
                mat_A[32][2] * mat_B[20][2] +
                mat_A[32][3] * mat_B[28][2] +
                mat_A[33][0] * mat_B[36][2] +
                mat_A[33][1] * mat_B[44][2] +
                mat_A[33][2] * mat_B[52][2] +
                mat_A[33][3] * mat_B[60][2] +
                mat_A[34][0] * mat_B[68][2] +
                mat_A[34][1] * mat_B[76][2] +
                mat_A[34][2] * mat_B[84][2] +
                mat_A[34][3] * mat_B[92][2] +
                mat_A[35][0] * mat_B[100][2] +
                mat_A[35][1] * mat_B[108][2] +
                mat_A[35][2] * mat_B[116][2] +
                mat_A[35][3] * mat_B[124][2] +
                mat_A[36][0] * mat_B[132][2] +
                mat_A[36][1] * mat_B[140][2] +
                mat_A[36][2] * mat_B[148][2] +
                mat_A[36][3] * mat_B[156][2] +
                mat_A[37][0] * mat_B[164][2] +
                mat_A[37][1] * mat_B[172][2] +
                mat_A[37][2] * mat_B[180][2] +
                mat_A[37][3] * mat_B[188][2] +
                mat_A[38][0] * mat_B[196][2] +
                mat_A[38][1] * mat_B[204][2] +
                mat_A[38][2] * mat_B[212][2] +
                mat_A[38][3] * mat_B[220][2] +
                mat_A[39][0] * mat_B[228][2] +
                mat_A[39][1] * mat_B[236][2] +
                mat_A[39][2] * mat_B[244][2] +
                mat_A[39][3] * mat_B[252][2];
    mat_C[36][3] <=
                mat_A[32][0] * mat_B[4][3] +
                mat_A[32][1] * mat_B[12][3] +
                mat_A[32][2] * mat_B[20][3] +
                mat_A[32][3] * mat_B[28][3] +
                mat_A[33][0] * mat_B[36][3] +
                mat_A[33][1] * mat_B[44][3] +
                mat_A[33][2] * mat_B[52][3] +
                mat_A[33][3] * mat_B[60][3] +
                mat_A[34][0] * mat_B[68][3] +
                mat_A[34][1] * mat_B[76][3] +
                mat_A[34][2] * mat_B[84][3] +
                mat_A[34][3] * mat_B[92][3] +
                mat_A[35][0] * mat_B[100][3] +
                mat_A[35][1] * mat_B[108][3] +
                mat_A[35][2] * mat_B[116][3] +
                mat_A[35][3] * mat_B[124][3] +
                mat_A[36][0] * mat_B[132][3] +
                mat_A[36][1] * mat_B[140][3] +
                mat_A[36][2] * mat_B[148][3] +
                mat_A[36][3] * mat_B[156][3] +
                mat_A[37][0] * mat_B[164][3] +
                mat_A[37][1] * mat_B[172][3] +
                mat_A[37][2] * mat_B[180][3] +
                mat_A[37][3] * mat_B[188][3] +
                mat_A[38][0] * mat_B[196][3] +
                mat_A[38][1] * mat_B[204][3] +
                mat_A[38][2] * mat_B[212][3] +
                mat_A[38][3] * mat_B[220][3] +
                mat_A[39][0] * mat_B[228][3] +
                mat_A[39][1] * mat_B[236][3] +
                mat_A[39][2] * mat_B[244][3] +
                mat_A[39][3] * mat_B[252][3];
    mat_C[37][0] <=
                mat_A[32][0] * mat_B[5][0] +
                mat_A[32][1] * mat_B[13][0] +
                mat_A[32][2] * mat_B[21][0] +
                mat_A[32][3] * mat_B[29][0] +
                mat_A[33][0] * mat_B[37][0] +
                mat_A[33][1] * mat_B[45][0] +
                mat_A[33][2] * mat_B[53][0] +
                mat_A[33][3] * mat_B[61][0] +
                mat_A[34][0] * mat_B[69][0] +
                mat_A[34][1] * mat_B[77][0] +
                mat_A[34][2] * mat_B[85][0] +
                mat_A[34][3] * mat_B[93][0] +
                mat_A[35][0] * mat_B[101][0] +
                mat_A[35][1] * mat_B[109][0] +
                mat_A[35][2] * mat_B[117][0] +
                mat_A[35][3] * mat_B[125][0] +
                mat_A[36][0] * mat_B[133][0] +
                mat_A[36][1] * mat_B[141][0] +
                mat_A[36][2] * mat_B[149][0] +
                mat_A[36][3] * mat_B[157][0] +
                mat_A[37][0] * mat_B[165][0] +
                mat_A[37][1] * mat_B[173][0] +
                mat_A[37][2] * mat_B[181][0] +
                mat_A[37][3] * mat_B[189][0] +
                mat_A[38][0] * mat_B[197][0] +
                mat_A[38][1] * mat_B[205][0] +
                mat_A[38][2] * mat_B[213][0] +
                mat_A[38][3] * mat_B[221][0] +
                mat_A[39][0] * mat_B[229][0] +
                mat_A[39][1] * mat_B[237][0] +
                mat_A[39][2] * mat_B[245][0] +
                mat_A[39][3] * mat_B[253][0];
    mat_C[37][1] <=
                mat_A[32][0] * mat_B[5][1] +
                mat_A[32][1] * mat_B[13][1] +
                mat_A[32][2] * mat_B[21][1] +
                mat_A[32][3] * mat_B[29][1] +
                mat_A[33][0] * mat_B[37][1] +
                mat_A[33][1] * mat_B[45][1] +
                mat_A[33][2] * mat_B[53][1] +
                mat_A[33][3] * mat_B[61][1] +
                mat_A[34][0] * mat_B[69][1] +
                mat_A[34][1] * mat_B[77][1] +
                mat_A[34][2] * mat_B[85][1] +
                mat_A[34][3] * mat_B[93][1] +
                mat_A[35][0] * mat_B[101][1] +
                mat_A[35][1] * mat_B[109][1] +
                mat_A[35][2] * mat_B[117][1] +
                mat_A[35][3] * mat_B[125][1] +
                mat_A[36][0] * mat_B[133][1] +
                mat_A[36][1] * mat_B[141][1] +
                mat_A[36][2] * mat_B[149][1] +
                mat_A[36][3] * mat_B[157][1] +
                mat_A[37][0] * mat_B[165][1] +
                mat_A[37][1] * mat_B[173][1] +
                mat_A[37][2] * mat_B[181][1] +
                mat_A[37][3] * mat_B[189][1] +
                mat_A[38][0] * mat_B[197][1] +
                mat_A[38][1] * mat_B[205][1] +
                mat_A[38][2] * mat_B[213][1] +
                mat_A[38][3] * mat_B[221][1] +
                mat_A[39][0] * mat_B[229][1] +
                mat_A[39][1] * mat_B[237][1] +
                mat_A[39][2] * mat_B[245][1] +
                mat_A[39][3] * mat_B[253][1];
    mat_C[37][2] <=
                mat_A[32][0] * mat_B[5][2] +
                mat_A[32][1] * mat_B[13][2] +
                mat_A[32][2] * mat_B[21][2] +
                mat_A[32][3] * mat_B[29][2] +
                mat_A[33][0] * mat_B[37][2] +
                mat_A[33][1] * mat_B[45][2] +
                mat_A[33][2] * mat_B[53][2] +
                mat_A[33][3] * mat_B[61][2] +
                mat_A[34][0] * mat_B[69][2] +
                mat_A[34][1] * mat_B[77][2] +
                mat_A[34][2] * mat_B[85][2] +
                mat_A[34][3] * mat_B[93][2] +
                mat_A[35][0] * mat_B[101][2] +
                mat_A[35][1] * mat_B[109][2] +
                mat_A[35][2] * mat_B[117][2] +
                mat_A[35][3] * mat_B[125][2] +
                mat_A[36][0] * mat_B[133][2] +
                mat_A[36][1] * mat_B[141][2] +
                mat_A[36][2] * mat_B[149][2] +
                mat_A[36][3] * mat_B[157][2] +
                mat_A[37][0] * mat_B[165][2] +
                mat_A[37][1] * mat_B[173][2] +
                mat_A[37][2] * mat_B[181][2] +
                mat_A[37][3] * mat_B[189][2] +
                mat_A[38][0] * mat_B[197][2] +
                mat_A[38][1] * mat_B[205][2] +
                mat_A[38][2] * mat_B[213][2] +
                mat_A[38][3] * mat_B[221][2] +
                mat_A[39][0] * mat_B[229][2] +
                mat_A[39][1] * mat_B[237][2] +
                mat_A[39][2] * mat_B[245][2] +
                mat_A[39][3] * mat_B[253][2];
    mat_C[37][3] <=
                mat_A[32][0] * mat_B[5][3] +
                mat_A[32][1] * mat_B[13][3] +
                mat_A[32][2] * mat_B[21][3] +
                mat_A[32][3] * mat_B[29][3] +
                mat_A[33][0] * mat_B[37][3] +
                mat_A[33][1] * mat_B[45][3] +
                mat_A[33][2] * mat_B[53][3] +
                mat_A[33][3] * mat_B[61][3] +
                mat_A[34][0] * mat_B[69][3] +
                mat_A[34][1] * mat_B[77][3] +
                mat_A[34][2] * mat_B[85][3] +
                mat_A[34][3] * mat_B[93][3] +
                mat_A[35][0] * mat_B[101][3] +
                mat_A[35][1] * mat_B[109][3] +
                mat_A[35][2] * mat_B[117][3] +
                mat_A[35][3] * mat_B[125][3] +
                mat_A[36][0] * mat_B[133][3] +
                mat_A[36][1] * mat_B[141][3] +
                mat_A[36][2] * mat_B[149][3] +
                mat_A[36][3] * mat_B[157][3] +
                mat_A[37][0] * mat_B[165][3] +
                mat_A[37][1] * mat_B[173][3] +
                mat_A[37][2] * mat_B[181][3] +
                mat_A[37][3] * mat_B[189][3] +
                mat_A[38][0] * mat_B[197][3] +
                mat_A[38][1] * mat_B[205][3] +
                mat_A[38][2] * mat_B[213][3] +
                mat_A[38][3] * mat_B[221][3] +
                mat_A[39][0] * mat_B[229][3] +
                mat_A[39][1] * mat_B[237][3] +
                mat_A[39][2] * mat_B[245][3] +
                mat_A[39][3] * mat_B[253][3];
    mat_C[38][0] <=
                mat_A[32][0] * mat_B[6][0] +
                mat_A[32][1] * mat_B[14][0] +
                mat_A[32][2] * mat_B[22][0] +
                mat_A[32][3] * mat_B[30][0] +
                mat_A[33][0] * mat_B[38][0] +
                mat_A[33][1] * mat_B[46][0] +
                mat_A[33][2] * mat_B[54][0] +
                mat_A[33][3] * mat_B[62][0] +
                mat_A[34][0] * mat_B[70][0] +
                mat_A[34][1] * mat_B[78][0] +
                mat_A[34][2] * mat_B[86][0] +
                mat_A[34][3] * mat_B[94][0] +
                mat_A[35][0] * mat_B[102][0] +
                mat_A[35][1] * mat_B[110][0] +
                mat_A[35][2] * mat_B[118][0] +
                mat_A[35][3] * mat_B[126][0] +
                mat_A[36][0] * mat_B[134][0] +
                mat_A[36][1] * mat_B[142][0] +
                mat_A[36][2] * mat_B[150][0] +
                mat_A[36][3] * mat_B[158][0] +
                mat_A[37][0] * mat_B[166][0] +
                mat_A[37][1] * mat_B[174][0] +
                mat_A[37][2] * mat_B[182][0] +
                mat_A[37][3] * mat_B[190][0] +
                mat_A[38][0] * mat_B[198][0] +
                mat_A[38][1] * mat_B[206][0] +
                mat_A[38][2] * mat_B[214][0] +
                mat_A[38][3] * mat_B[222][0] +
                mat_A[39][0] * mat_B[230][0] +
                mat_A[39][1] * mat_B[238][0] +
                mat_A[39][2] * mat_B[246][0] +
                mat_A[39][3] * mat_B[254][0];
    mat_C[38][1] <=
                mat_A[32][0] * mat_B[6][1] +
                mat_A[32][1] * mat_B[14][1] +
                mat_A[32][2] * mat_B[22][1] +
                mat_A[32][3] * mat_B[30][1] +
                mat_A[33][0] * mat_B[38][1] +
                mat_A[33][1] * mat_B[46][1] +
                mat_A[33][2] * mat_B[54][1] +
                mat_A[33][3] * mat_B[62][1] +
                mat_A[34][0] * mat_B[70][1] +
                mat_A[34][1] * mat_B[78][1] +
                mat_A[34][2] * mat_B[86][1] +
                mat_A[34][3] * mat_B[94][1] +
                mat_A[35][0] * mat_B[102][1] +
                mat_A[35][1] * mat_B[110][1] +
                mat_A[35][2] * mat_B[118][1] +
                mat_A[35][3] * mat_B[126][1] +
                mat_A[36][0] * mat_B[134][1] +
                mat_A[36][1] * mat_B[142][1] +
                mat_A[36][2] * mat_B[150][1] +
                mat_A[36][3] * mat_B[158][1] +
                mat_A[37][0] * mat_B[166][1] +
                mat_A[37][1] * mat_B[174][1] +
                mat_A[37][2] * mat_B[182][1] +
                mat_A[37][3] * mat_B[190][1] +
                mat_A[38][0] * mat_B[198][1] +
                mat_A[38][1] * mat_B[206][1] +
                mat_A[38][2] * mat_B[214][1] +
                mat_A[38][3] * mat_B[222][1] +
                mat_A[39][0] * mat_B[230][1] +
                mat_A[39][1] * mat_B[238][1] +
                mat_A[39][2] * mat_B[246][1] +
                mat_A[39][3] * mat_B[254][1];
    mat_C[38][2] <=
                mat_A[32][0] * mat_B[6][2] +
                mat_A[32][1] * mat_B[14][2] +
                mat_A[32][2] * mat_B[22][2] +
                mat_A[32][3] * mat_B[30][2] +
                mat_A[33][0] * mat_B[38][2] +
                mat_A[33][1] * mat_B[46][2] +
                mat_A[33][2] * mat_B[54][2] +
                mat_A[33][3] * mat_B[62][2] +
                mat_A[34][0] * mat_B[70][2] +
                mat_A[34][1] * mat_B[78][2] +
                mat_A[34][2] * mat_B[86][2] +
                mat_A[34][3] * mat_B[94][2] +
                mat_A[35][0] * mat_B[102][2] +
                mat_A[35][1] * mat_B[110][2] +
                mat_A[35][2] * mat_B[118][2] +
                mat_A[35][3] * mat_B[126][2] +
                mat_A[36][0] * mat_B[134][2] +
                mat_A[36][1] * mat_B[142][2] +
                mat_A[36][2] * mat_B[150][2] +
                mat_A[36][3] * mat_B[158][2] +
                mat_A[37][0] * mat_B[166][2] +
                mat_A[37][1] * mat_B[174][2] +
                mat_A[37][2] * mat_B[182][2] +
                mat_A[37][3] * mat_B[190][2] +
                mat_A[38][0] * mat_B[198][2] +
                mat_A[38][1] * mat_B[206][2] +
                mat_A[38][2] * mat_B[214][2] +
                mat_A[38][3] * mat_B[222][2] +
                mat_A[39][0] * mat_B[230][2] +
                mat_A[39][1] * mat_B[238][2] +
                mat_A[39][2] * mat_B[246][2] +
                mat_A[39][3] * mat_B[254][2];
    mat_C[38][3] <=
                mat_A[32][0] * mat_B[6][3] +
                mat_A[32][1] * mat_B[14][3] +
                mat_A[32][2] * mat_B[22][3] +
                mat_A[32][3] * mat_B[30][3] +
                mat_A[33][0] * mat_B[38][3] +
                mat_A[33][1] * mat_B[46][3] +
                mat_A[33][2] * mat_B[54][3] +
                mat_A[33][3] * mat_B[62][3] +
                mat_A[34][0] * mat_B[70][3] +
                mat_A[34][1] * mat_B[78][3] +
                mat_A[34][2] * mat_B[86][3] +
                mat_A[34][3] * mat_B[94][3] +
                mat_A[35][0] * mat_B[102][3] +
                mat_A[35][1] * mat_B[110][3] +
                mat_A[35][2] * mat_B[118][3] +
                mat_A[35][3] * mat_B[126][3] +
                mat_A[36][0] * mat_B[134][3] +
                mat_A[36][1] * mat_B[142][3] +
                mat_A[36][2] * mat_B[150][3] +
                mat_A[36][3] * mat_B[158][3] +
                mat_A[37][0] * mat_B[166][3] +
                mat_A[37][1] * mat_B[174][3] +
                mat_A[37][2] * mat_B[182][3] +
                mat_A[37][3] * mat_B[190][3] +
                mat_A[38][0] * mat_B[198][3] +
                mat_A[38][1] * mat_B[206][3] +
                mat_A[38][2] * mat_B[214][3] +
                mat_A[38][3] * mat_B[222][3] +
                mat_A[39][0] * mat_B[230][3] +
                mat_A[39][1] * mat_B[238][3] +
                mat_A[39][2] * mat_B[246][3] +
                mat_A[39][3] * mat_B[254][3];
    mat_C[39][0] <=
                mat_A[32][0] * mat_B[7][0] +
                mat_A[32][1] * mat_B[15][0] +
                mat_A[32][2] * mat_B[23][0] +
                mat_A[32][3] * mat_B[31][0] +
                mat_A[33][0] * mat_B[39][0] +
                mat_A[33][1] * mat_B[47][0] +
                mat_A[33][2] * mat_B[55][0] +
                mat_A[33][3] * mat_B[63][0] +
                mat_A[34][0] * mat_B[71][0] +
                mat_A[34][1] * mat_B[79][0] +
                mat_A[34][2] * mat_B[87][0] +
                mat_A[34][3] * mat_B[95][0] +
                mat_A[35][0] * mat_B[103][0] +
                mat_A[35][1] * mat_B[111][0] +
                mat_A[35][2] * mat_B[119][0] +
                mat_A[35][3] * mat_B[127][0] +
                mat_A[36][0] * mat_B[135][0] +
                mat_A[36][1] * mat_B[143][0] +
                mat_A[36][2] * mat_B[151][0] +
                mat_A[36][3] * mat_B[159][0] +
                mat_A[37][0] * mat_B[167][0] +
                mat_A[37][1] * mat_B[175][0] +
                mat_A[37][2] * mat_B[183][0] +
                mat_A[37][3] * mat_B[191][0] +
                mat_A[38][0] * mat_B[199][0] +
                mat_A[38][1] * mat_B[207][0] +
                mat_A[38][2] * mat_B[215][0] +
                mat_A[38][3] * mat_B[223][0] +
                mat_A[39][0] * mat_B[231][0] +
                mat_A[39][1] * mat_B[239][0] +
                mat_A[39][2] * mat_B[247][0] +
                mat_A[39][3] * mat_B[255][0];
    mat_C[39][1] <=
                mat_A[32][0] * mat_B[7][1] +
                mat_A[32][1] * mat_B[15][1] +
                mat_A[32][2] * mat_B[23][1] +
                mat_A[32][3] * mat_B[31][1] +
                mat_A[33][0] * mat_B[39][1] +
                mat_A[33][1] * mat_B[47][1] +
                mat_A[33][2] * mat_B[55][1] +
                mat_A[33][3] * mat_B[63][1] +
                mat_A[34][0] * mat_B[71][1] +
                mat_A[34][1] * mat_B[79][1] +
                mat_A[34][2] * mat_B[87][1] +
                mat_A[34][3] * mat_B[95][1] +
                mat_A[35][0] * mat_B[103][1] +
                mat_A[35][1] * mat_B[111][1] +
                mat_A[35][2] * mat_B[119][1] +
                mat_A[35][3] * mat_B[127][1] +
                mat_A[36][0] * mat_B[135][1] +
                mat_A[36][1] * mat_B[143][1] +
                mat_A[36][2] * mat_B[151][1] +
                mat_A[36][3] * mat_B[159][1] +
                mat_A[37][0] * mat_B[167][1] +
                mat_A[37][1] * mat_B[175][1] +
                mat_A[37][2] * mat_B[183][1] +
                mat_A[37][3] * mat_B[191][1] +
                mat_A[38][0] * mat_B[199][1] +
                mat_A[38][1] * mat_B[207][1] +
                mat_A[38][2] * mat_B[215][1] +
                mat_A[38][3] * mat_B[223][1] +
                mat_A[39][0] * mat_B[231][1] +
                mat_A[39][1] * mat_B[239][1] +
                mat_A[39][2] * mat_B[247][1] +
                mat_A[39][3] * mat_B[255][1];
    mat_C[39][2] <=
                mat_A[32][0] * mat_B[7][2] +
                mat_A[32][1] * mat_B[15][2] +
                mat_A[32][2] * mat_B[23][2] +
                mat_A[32][3] * mat_B[31][2] +
                mat_A[33][0] * mat_B[39][2] +
                mat_A[33][1] * mat_B[47][2] +
                mat_A[33][2] * mat_B[55][2] +
                mat_A[33][3] * mat_B[63][2] +
                mat_A[34][0] * mat_B[71][2] +
                mat_A[34][1] * mat_B[79][2] +
                mat_A[34][2] * mat_B[87][2] +
                mat_A[34][3] * mat_B[95][2] +
                mat_A[35][0] * mat_B[103][2] +
                mat_A[35][1] * mat_B[111][2] +
                mat_A[35][2] * mat_B[119][2] +
                mat_A[35][3] * mat_B[127][2] +
                mat_A[36][0] * mat_B[135][2] +
                mat_A[36][1] * mat_B[143][2] +
                mat_A[36][2] * mat_B[151][2] +
                mat_A[36][3] * mat_B[159][2] +
                mat_A[37][0] * mat_B[167][2] +
                mat_A[37][1] * mat_B[175][2] +
                mat_A[37][2] * mat_B[183][2] +
                mat_A[37][3] * mat_B[191][2] +
                mat_A[38][0] * mat_B[199][2] +
                mat_A[38][1] * mat_B[207][2] +
                mat_A[38][2] * mat_B[215][2] +
                mat_A[38][3] * mat_B[223][2] +
                mat_A[39][0] * mat_B[231][2] +
                mat_A[39][1] * mat_B[239][2] +
                mat_A[39][2] * mat_B[247][2] +
                mat_A[39][3] * mat_B[255][2];
    mat_C[39][3] <=
                mat_A[32][0] * mat_B[7][3] +
                mat_A[32][1] * mat_B[15][3] +
                mat_A[32][2] * mat_B[23][3] +
                mat_A[32][3] * mat_B[31][3] +
                mat_A[33][0] * mat_B[39][3] +
                mat_A[33][1] * mat_B[47][3] +
                mat_A[33][2] * mat_B[55][3] +
                mat_A[33][3] * mat_B[63][3] +
                mat_A[34][0] * mat_B[71][3] +
                mat_A[34][1] * mat_B[79][3] +
                mat_A[34][2] * mat_B[87][3] +
                mat_A[34][3] * mat_B[95][3] +
                mat_A[35][0] * mat_B[103][3] +
                mat_A[35][1] * mat_B[111][3] +
                mat_A[35][2] * mat_B[119][3] +
                mat_A[35][3] * mat_B[127][3] +
                mat_A[36][0] * mat_B[135][3] +
                mat_A[36][1] * mat_B[143][3] +
                mat_A[36][2] * mat_B[151][3] +
                mat_A[36][3] * mat_B[159][3] +
                mat_A[37][0] * mat_B[167][3] +
                mat_A[37][1] * mat_B[175][3] +
                mat_A[37][2] * mat_B[183][3] +
                mat_A[37][3] * mat_B[191][3] +
                mat_A[38][0] * mat_B[199][3] +
                mat_A[38][1] * mat_B[207][3] +
                mat_A[38][2] * mat_B[215][3] +
                mat_A[38][3] * mat_B[223][3] +
                mat_A[39][0] * mat_B[231][3] +
                mat_A[39][1] * mat_B[239][3] +
                mat_A[39][2] * mat_B[247][3] +
                mat_A[39][3] * mat_B[255][3];
    mat_C[40][0] <=
                mat_A[40][0] * mat_B[0][0] +
                mat_A[40][1] * mat_B[8][0] +
                mat_A[40][2] * mat_B[16][0] +
                mat_A[40][3] * mat_B[24][0] +
                mat_A[41][0] * mat_B[32][0] +
                mat_A[41][1] * mat_B[40][0] +
                mat_A[41][2] * mat_B[48][0] +
                mat_A[41][3] * mat_B[56][0] +
                mat_A[42][0] * mat_B[64][0] +
                mat_A[42][1] * mat_B[72][0] +
                mat_A[42][2] * mat_B[80][0] +
                mat_A[42][3] * mat_B[88][0] +
                mat_A[43][0] * mat_B[96][0] +
                mat_A[43][1] * mat_B[104][0] +
                mat_A[43][2] * mat_B[112][0] +
                mat_A[43][3] * mat_B[120][0] +
                mat_A[44][0] * mat_B[128][0] +
                mat_A[44][1] * mat_B[136][0] +
                mat_A[44][2] * mat_B[144][0] +
                mat_A[44][3] * mat_B[152][0] +
                mat_A[45][0] * mat_B[160][0] +
                mat_A[45][1] * mat_B[168][0] +
                mat_A[45][2] * mat_B[176][0] +
                mat_A[45][3] * mat_B[184][0] +
                mat_A[46][0] * mat_B[192][0] +
                mat_A[46][1] * mat_B[200][0] +
                mat_A[46][2] * mat_B[208][0] +
                mat_A[46][3] * mat_B[216][0] +
                mat_A[47][0] * mat_B[224][0] +
                mat_A[47][1] * mat_B[232][0] +
                mat_A[47][2] * mat_B[240][0] +
                mat_A[47][3] * mat_B[248][0];
    mat_C[40][1] <=
                mat_A[40][0] * mat_B[0][1] +
                mat_A[40][1] * mat_B[8][1] +
                mat_A[40][2] * mat_B[16][1] +
                mat_A[40][3] * mat_B[24][1] +
                mat_A[41][0] * mat_B[32][1] +
                mat_A[41][1] * mat_B[40][1] +
                mat_A[41][2] * mat_B[48][1] +
                mat_A[41][3] * mat_B[56][1] +
                mat_A[42][0] * mat_B[64][1] +
                mat_A[42][1] * mat_B[72][1] +
                mat_A[42][2] * mat_B[80][1] +
                mat_A[42][3] * mat_B[88][1] +
                mat_A[43][0] * mat_B[96][1] +
                mat_A[43][1] * mat_B[104][1] +
                mat_A[43][2] * mat_B[112][1] +
                mat_A[43][3] * mat_B[120][1] +
                mat_A[44][0] * mat_B[128][1] +
                mat_A[44][1] * mat_B[136][1] +
                mat_A[44][2] * mat_B[144][1] +
                mat_A[44][3] * mat_B[152][1] +
                mat_A[45][0] * mat_B[160][1] +
                mat_A[45][1] * mat_B[168][1] +
                mat_A[45][2] * mat_B[176][1] +
                mat_A[45][3] * mat_B[184][1] +
                mat_A[46][0] * mat_B[192][1] +
                mat_A[46][1] * mat_B[200][1] +
                mat_A[46][2] * mat_B[208][1] +
                mat_A[46][3] * mat_B[216][1] +
                mat_A[47][0] * mat_B[224][1] +
                mat_A[47][1] * mat_B[232][1] +
                mat_A[47][2] * mat_B[240][1] +
                mat_A[47][3] * mat_B[248][1];
    mat_C[40][2] <=
                mat_A[40][0] * mat_B[0][2] +
                mat_A[40][1] * mat_B[8][2] +
                mat_A[40][2] * mat_B[16][2] +
                mat_A[40][3] * mat_B[24][2] +
                mat_A[41][0] * mat_B[32][2] +
                mat_A[41][1] * mat_B[40][2] +
                mat_A[41][2] * mat_B[48][2] +
                mat_A[41][3] * mat_B[56][2] +
                mat_A[42][0] * mat_B[64][2] +
                mat_A[42][1] * mat_B[72][2] +
                mat_A[42][2] * mat_B[80][2] +
                mat_A[42][3] * mat_B[88][2] +
                mat_A[43][0] * mat_B[96][2] +
                mat_A[43][1] * mat_B[104][2] +
                mat_A[43][2] * mat_B[112][2] +
                mat_A[43][3] * mat_B[120][2] +
                mat_A[44][0] * mat_B[128][2] +
                mat_A[44][1] * mat_B[136][2] +
                mat_A[44][2] * mat_B[144][2] +
                mat_A[44][3] * mat_B[152][2] +
                mat_A[45][0] * mat_B[160][2] +
                mat_A[45][1] * mat_B[168][2] +
                mat_A[45][2] * mat_B[176][2] +
                mat_A[45][3] * mat_B[184][2] +
                mat_A[46][0] * mat_B[192][2] +
                mat_A[46][1] * mat_B[200][2] +
                mat_A[46][2] * mat_B[208][2] +
                mat_A[46][3] * mat_B[216][2] +
                mat_A[47][0] * mat_B[224][2] +
                mat_A[47][1] * mat_B[232][2] +
                mat_A[47][2] * mat_B[240][2] +
                mat_A[47][3] * mat_B[248][2];
    mat_C[40][3] <=
                mat_A[40][0] * mat_B[0][3] +
                mat_A[40][1] * mat_B[8][3] +
                mat_A[40][2] * mat_B[16][3] +
                mat_A[40][3] * mat_B[24][3] +
                mat_A[41][0] * mat_B[32][3] +
                mat_A[41][1] * mat_B[40][3] +
                mat_A[41][2] * mat_B[48][3] +
                mat_A[41][3] * mat_B[56][3] +
                mat_A[42][0] * mat_B[64][3] +
                mat_A[42][1] * mat_B[72][3] +
                mat_A[42][2] * mat_B[80][3] +
                mat_A[42][3] * mat_B[88][3] +
                mat_A[43][0] * mat_B[96][3] +
                mat_A[43][1] * mat_B[104][3] +
                mat_A[43][2] * mat_B[112][3] +
                mat_A[43][3] * mat_B[120][3] +
                mat_A[44][0] * mat_B[128][3] +
                mat_A[44][1] * mat_B[136][3] +
                mat_A[44][2] * mat_B[144][3] +
                mat_A[44][3] * mat_B[152][3] +
                mat_A[45][0] * mat_B[160][3] +
                mat_A[45][1] * mat_B[168][3] +
                mat_A[45][2] * mat_B[176][3] +
                mat_A[45][3] * mat_B[184][3] +
                mat_A[46][0] * mat_B[192][3] +
                mat_A[46][1] * mat_B[200][3] +
                mat_A[46][2] * mat_B[208][3] +
                mat_A[46][3] * mat_B[216][3] +
                mat_A[47][0] * mat_B[224][3] +
                mat_A[47][1] * mat_B[232][3] +
                mat_A[47][2] * mat_B[240][3] +
                mat_A[47][3] * mat_B[248][3];
    mat_C[41][0] <=
                mat_A[40][0] * mat_B[1][0] +
                mat_A[40][1] * mat_B[9][0] +
                mat_A[40][2] * mat_B[17][0] +
                mat_A[40][3] * mat_B[25][0] +
                mat_A[41][0] * mat_B[33][0] +
                mat_A[41][1] * mat_B[41][0] +
                mat_A[41][2] * mat_B[49][0] +
                mat_A[41][3] * mat_B[57][0] +
                mat_A[42][0] * mat_B[65][0] +
                mat_A[42][1] * mat_B[73][0] +
                mat_A[42][2] * mat_B[81][0] +
                mat_A[42][3] * mat_B[89][0] +
                mat_A[43][0] * mat_B[97][0] +
                mat_A[43][1] * mat_B[105][0] +
                mat_A[43][2] * mat_B[113][0] +
                mat_A[43][3] * mat_B[121][0] +
                mat_A[44][0] * mat_B[129][0] +
                mat_A[44][1] * mat_B[137][0] +
                mat_A[44][2] * mat_B[145][0] +
                mat_A[44][3] * mat_B[153][0] +
                mat_A[45][0] * mat_B[161][0] +
                mat_A[45][1] * mat_B[169][0] +
                mat_A[45][2] * mat_B[177][0] +
                mat_A[45][3] * mat_B[185][0] +
                mat_A[46][0] * mat_B[193][0] +
                mat_A[46][1] * mat_B[201][0] +
                mat_A[46][2] * mat_B[209][0] +
                mat_A[46][3] * mat_B[217][0] +
                mat_A[47][0] * mat_B[225][0] +
                mat_A[47][1] * mat_B[233][0] +
                mat_A[47][2] * mat_B[241][0] +
                mat_A[47][3] * mat_B[249][0];
    mat_C[41][1] <=
                mat_A[40][0] * mat_B[1][1] +
                mat_A[40][1] * mat_B[9][1] +
                mat_A[40][2] * mat_B[17][1] +
                mat_A[40][3] * mat_B[25][1] +
                mat_A[41][0] * mat_B[33][1] +
                mat_A[41][1] * mat_B[41][1] +
                mat_A[41][2] * mat_B[49][1] +
                mat_A[41][3] * mat_B[57][1] +
                mat_A[42][0] * mat_B[65][1] +
                mat_A[42][1] * mat_B[73][1] +
                mat_A[42][2] * mat_B[81][1] +
                mat_A[42][3] * mat_B[89][1] +
                mat_A[43][0] * mat_B[97][1] +
                mat_A[43][1] * mat_B[105][1] +
                mat_A[43][2] * mat_B[113][1] +
                mat_A[43][3] * mat_B[121][1] +
                mat_A[44][0] * mat_B[129][1] +
                mat_A[44][1] * mat_B[137][1] +
                mat_A[44][2] * mat_B[145][1] +
                mat_A[44][3] * mat_B[153][1] +
                mat_A[45][0] * mat_B[161][1] +
                mat_A[45][1] * mat_B[169][1] +
                mat_A[45][2] * mat_B[177][1] +
                mat_A[45][3] * mat_B[185][1] +
                mat_A[46][0] * mat_B[193][1] +
                mat_A[46][1] * mat_B[201][1] +
                mat_A[46][2] * mat_B[209][1] +
                mat_A[46][3] * mat_B[217][1] +
                mat_A[47][0] * mat_B[225][1] +
                mat_A[47][1] * mat_B[233][1] +
                mat_A[47][2] * mat_B[241][1] +
                mat_A[47][3] * mat_B[249][1];
    mat_C[41][2] <=
                mat_A[40][0] * mat_B[1][2] +
                mat_A[40][1] * mat_B[9][2] +
                mat_A[40][2] * mat_B[17][2] +
                mat_A[40][3] * mat_B[25][2] +
                mat_A[41][0] * mat_B[33][2] +
                mat_A[41][1] * mat_B[41][2] +
                mat_A[41][2] * mat_B[49][2] +
                mat_A[41][3] * mat_B[57][2] +
                mat_A[42][0] * mat_B[65][2] +
                mat_A[42][1] * mat_B[73][2] +
                mat_A[42][2] * mat_B[81][2] +
                mat_A[42][3] * mat_B[89][2] +
                mat_A[43][0] * mat_B[97][2] +
                mat_A[43][1] * mat_B[105][2] +
                mat_A[43][2] * mat_B[113][2] +
                mat_A[43][3] * mat_B[121][2] +
                mat_A[44][0] * mat_B[129][2] +
                mat_A[44][1] * mat_B[137][2] +
                mat_A[44][2] * mat_B[145][2] +
                mat_A[44][3] * mat_B[153][2] +
                mat_A[45][0] * mat_B[161][2] +
                mat_A[45][1] * mat_B[169][2] +
                mat_A[45][2] * mat_B[177][2] +
                mat_A[45][3] * mat_B[185][2] +
                mat_A[46][0] * mat_B[193][2] +
                mat_A[46][1] * mat_B[201][2] +
                mat_A[46][2] * mat_B[209][2] +
                mat_A[46][3] * mat_B[217][2] +
                mat_A[47][0] * mat_B[225][2] +
                mat_A[47][1] * mat_B[233][2] +
                mat_A[47][2] * mat_B[241][2] +
                mat_A[47][3] * mat_B[249][2];
    mat_C[41][3] <=
                mat_A[40][0] * mat_B[1][3] +
                mat_A[40][1] * mat_B[9][3] +
                mat_A[40][2] * mat_B[17][3] +
                mat_A[40][3] * mat_B[25][3] +
                mat_A[41][0] * mat_B[33][3] +
                mat_A[41][1] * mat_B[41][3] +
                mat_A[41][2] * mat_B[49][3] +
                mat_A[41][3] * mat_B[57][3] +
                mat_A[42][0] * mat_B[65][3] +
                mat_A[42][1] * mat_B[73][3] +
                mat_A[42][2] * mat_B[81][3] +
                mat_A[42][3] * mat_B[89][3] +
                mat_A[43][0] * mat_B[97][3] +
                mat_A[43][1] * mat_B[105][3] +
                mat_A[43][2] * mat_B[113][3] +
                mat_A[43][3] * mat_B[121][3] +
                mat_A[44][0] * mat_B[129][3] +
                mat_A[44][1] * mat_B[137][3] +
                mat_A[44][2] * mat_B[145][3] +
                mat_A[44][3] * mat_B[153][3] +
                mat_A[45][0] * mat_B[161][3] +
                mat_A[45][1] * mat_B[169][3] +
                mat_A[45][2] * mat_B[177][3] +
                mat_A[45][3] * mat_B[185][3] +
                mat_A[46][0] * mat_B[193][3] +
                mat_A[46][1] * mat_B[201][3] +
                mat_A[46][2] * mat_B[209][3] +
                mat_A[46][3] * mat_B[217][3] +
                mat_A[47][0] * mat_B[225][3] +
                mat_A[47][1] * mat_B[233][3] +
                mat_A[47][2] * mat_B[241][3] +
                mat_A[47][3] * mat_B[249][3];
    mat_C[42][0] <=
                mat_A[40][0] * mat_B[2][0] +
                mat_A[40][1] * mat_B[10][0] +
                mat_A[40][2] * mat_B[18][0] +
                mat_A[40][3] * mat_B[26][0] +
                mat_A[41][0] * mat_B[34][0] +
                mat_A[41][1] * mat_B[42][0] +
                mat_A[41][2] * mat_B[50][0] +
                mat_A[41][3] * mat_B[58][0] +
                mat_A[42][0] * mat_B[66][0] +
                mat_A[42][1] * mat_B[74][0] +
                mat_A[42][2] * mat_B[82][0] +
                mat_A[42][3] * mat_B[90][0] +
                mat_A[43][0] * mat_B[98][0] +
                mat_A[43][1] * mat_B[106][0] +
                mat_A[43][2] * mat_B[114][0] +
                mat_A[43][3] * mat_B[122][0] +
                mat_A[44][0] * mat_B[130][0] +
                mat_A[44][1] * mat_B[138][0] +
                mat_A[44][2] * mat_B[146][0] +
                mat_A[44][3] * mat_B[154][0] +
                mat_A[45][0] * mat_B[162][0] +
                mat_A[45][1] * mat_B[170][0] +
                mat_A[45][2] * mat_B[178][0] +
                mat_A[45][3] * mat_B[186][0] +
                mat_A[46][0] * mat_B[194][0] +
                mat_A[46][1] * mat_B[202][0] +
                mat_A[46][2] * mat_B[210][0] +
                mat_A[46][3] * mat_B[218][0] +
                mat_A[47][0] * mat_B[226][0] +
                mat_A[47][1] * mat_B[234][0] +
                mat_A[47][2] * mat_B[242][0] +
                mat_A[47][3] * mat_B[250][0];
    mat_C[42][1] <=
                mat_A[40][0] * mat_B[2][1] +
                mat_A[40][1] * mat_B[10][1] +
                mat_A[40][2] * mat_B[18][1] +
                mat_A[40][3] * mat_B[26][1] +
                mat_A[41][0] * mat_B[34][1] +
                mat_A[41][1] * mat_B[42][1] +
                mat_A[41][2] * mat_B[50][1] +
                mat_A[41][3] * mat_B[58][1] +
                mat_A[42][0] * mat_B[66][1] +
                mat_A[42][1] * mat_B[74][1] +
                mat_A[42][2] * mat_B[82][1] +
                mat_A[42][3] * mat_B[90][1] +
                mat_A[43][0] * mat_B[98][1] +
                mat_A[43][1] * mat_B[106][1] +
                mat_A[43][2] * mat_B[114][1] +
                mat_A[43][3] * mat_B[122][1] +
                mat_A[44][0] * mat_B[130][1] +
                mat_A[44][1] * mat_B[138][1] +
                mat_A[44][2] * mat_B[146][1] +
                mat_A[44][3] * mat_B[154][1] +
                mat_A[45][0] * mat_B[162][1] +
                mat_A[45][1] * mat_B[170][1] +
                mat_A[45][2] * mat_B[178][1] +
                mat_A[45][3] * mat_B[186][1] +
                mat_A[46][0] * mat_B[194][1] +
                mat_A[46][1] * mat_B[202][1] +
                mat_A[46][2] * mat_B[210][1] +
                mat_A[46][3] * mat_B[218][1] +
                mat_A[47][0] * mat_B[226][1] +
                mat_A[47][1] * mat_B[234][1] +
                mat_A[47][2] * mat_B[242][1] +
                mat_A[47][3] * mat_B[250][1];
    mat_C[42][2] <=
                mat_A[40][0] * mat_B[2][2] +
                mat_A[40][1] * mat_B[10][2] +
                mat_A[40][2] * mat_B[18][2] +
                mat_A[40][3] * mat_B[26][2] +
                mat_A[41][0] * mat_B[34][2] +
                mat_A[41][1] * mat_B[42][2] +
                mat_A[41][2] * mat_B[50][2] +
                mat_A[41][3] * mat_B[58][2] +
                mat_A[42][0] * mat_B[66][2] +
                mat_A[42][1] * mat_B[74][2] +
                mat_A[42][2] * mat_B[82][2] +
                mat_A[42][3] * mat_B[90][2] +
                mat_A[43][0] * mat_B[98][2] +
                mat_A[43][1] * mat_B[106][2] +
                mat_A[43][2] * mat_B[114][2] +
                mat_A[43][3] * mat_B[122][2] +
                mat_A[44][0] * mat_B[130][2] +
                mat_A[44][1] * mat_B[138][2] +
                mat_A[44][2] * mat_B[146][2] +
                mat_A[44][3] * mat_B[154][2] +
                mat_A[45][0] * mat_B[162][2] +
                mat_A[45][1] * mat_B[170][2] +
                mat_A[45][2] * mat_B[178][2] +
                mat_A[45][3] * mat_B[186][2] +
                mat_A[46][0] * mat_B[194][2] +
                mat_A[46][1] * mat_B[202][2] +
                mat_A[46][2] * mat_B[210][2] +
                mat_A[46][3] * mat_B[218][2] +
                mat_A[47][0] * mat_B[226][2] +
                mat_A[47][1] * mat_B[234][2] +
                mat_A[47][2] * mat_B[242][2] +
                mat_A[47][3] * mat_B[250][2];
    mat_C[42][3] <=
                mat_A[40][0] * mat_B[2][3] +
                mat_A[40][1] * mat_B[10][3] +
                mat_A[40][2] * mat_B[18][3] +
                mat_A[40][3] * mat_B[26][3] +
                mat_A[41][0] * mat_B[34][3] +
                mat_A[41][1] * mat_B[42][3] +
                mat_A[41][2] * mat_B[50][3] +
                mat_A[41][3] * mat_B[58][3] +
                mat_A[42][0] * mat_B[66][3] +
                mat_A[42][1] * mat_B[74][3] +
                mat_A[42][2] * mat_B[82][3] +
                mat_A[42][3] * mat_B[90][3] +
                mat_A[43][0] * mat_B[98][3] +
                mat_A[43][1] * mat_B[106][3] +
                mat_A[43][2] * mat_B[114][3] +
                mat_A[43][3] * mat_B[122][3] +
                mat_A[44][0] * mat_B[130][3] +
                mat_A[44][1] * mat_B[138][3] +
                mat_A[44][2] * mat_B[146][3] +
                mat_A[44][3] * mat_B[154][3] +
                mat_A[45][0] * mat_B[162][3] +
                mat_A[45][1] * mat_B[170][3] +
                mat_A[45][2] * mat_B[178][3] +
                mat_A[45][3] * mat_B[186][3] +
                mat_A[46][0] * mat_B[194][3] +
                mat_A[46][1] * mat_B[202][3] +
                mat_A[46][2] * mat_B[210][3] +
                mat_A[46][3] * mat_B[218][3] +
                mat_A[47][0] * mat_B[226][3] +
                mat_A[47][1] * mat_B[234][3] +
                mat_A[47][2] * mat_B[242][3] +
                mat_A[47][3] * mat_B[250][3];
    mat_C[43][0] <=
                mat_A[40][0] * mat_B[3][0] +
                mat_A[40][1] * mat_B[11][0] +
                mat_A[40][2] * mat_B[19][0] +
                mat_A[40][3] * mat_B[27][0] +
                mat_A[41][0] * mat_B[35][0] +
                mat_A[41][1] * mat_B[43][0] +
                mat_A[41][2] * mat_B[51][0] +
                mat_A[41][3] * mat_B[59][0] +
                mat_A[42][0] * mat_B[67][0] +
                mat_A[42][1] * mat_B[75][0] +
                mat_A[42][2] * mat_B[83][0] +
                mat_A[42][3] * mat_B[91][0] +
                mat_A[43][0] * mat_B[99][0] +
                mat_A[43][1] * mat_B[107][0] +
                mat_A[43][2] * mat_B[115][0] +
                mat_A[43][3] * mat_B[123][0] +
                mat_A[44][0] * mat_B[131][0] +
                mat_A[44][1] * mat_B[139][0] +
                mat_A[44][2] * mat_B[147][0] +
                mat_A[44][3] * mat_B[155][0] +
                mat_A[45][0] * mat_B[163][0] +
                mat_A[45][1] * mat_B[171][0] +
                mat_A[45][2] * mat_B[179][0] +
                mat_A[45][3] * mat_B[187][0] +
                mat_A[46][0] * mat_B[195][0] +
                mat_A[46][1] * mat_B[203][0] +
                mat_A[46][2] * mat_B[211][0] +
                mat_A[46][3] * mat_B[219][0] +
                mat_A[47][0] * mat_B[227][0] +
                mat_A[47][1] * mat_B[235][0] +
                mat_A[47][2] * mat_B[243][0] +
                mat_A[47][3] * mat_B[251][0];
    mat_C[43][1] <=
                mat_A[40][0] * mat_B[3][1] +
                mat_A[40][1] * mat_B[11][1] +
                mat_A[40][2] * mat_B[19][1] +
                mat_A[40][3] * mat_B[27][1] +
                mat_A[41][0] * mat_B[35][1] +
                mat_A[41][1] * mat_B[43][1] +
                mat_A[41][2] * mat_B[51][1] +
                mat_A[41][3] * mat_B[59][1] +
                mat_A[42][0] * mat_B[67][1] +
                mat_A[42][1] * mat_B[75][1] +
                mat_A[42][2] * mat_B[83][1] +
                mat_A[42][3] * mat_B[91][1] +
                mat_A[43][0] * mat_B[99][1] +
                mat_A[43][1] * mat_B[107][1] +
                mat_A[43][2] * mat_B[115][1] +
                mat_A[43][3] * mat_B[123][1] +
                mat_A[44][0] * mat_B[131][1] +
                mat_A[44][1] * mat_B[139][1] +
                mat_A[44][2] * mat_B[147][1] +
                mat_A[44][3] * mat_B[155][1] +
                mat_A[45][0] * mat_B[163][1] +
                mat_A[45][1] * mat_B[171][1] +
                mat_A[45][2] * mat_B[179][1] +
                mat_A[45][3] * mat_B[187][1] +
                mat_A[46][0] * mat_B[195][1] +
                mat_A[46][1] * mat_B[203][1] +
                mat_A[46][2] * mat_B[211][1] +
                mat_A[46][3] * mat_B[219][1] +
                mat_A[47][0] * mat_B[227][1] +
                mat_A[47][1] * mat_B[235][1] +
                mat_A[47][2] * mat_B[243][1] +
                mat_A[47][3] * mat_B[251][1];
    mat_C[43][2] <=
                mat_A[40][0] * mat_B[3][2] +
                mat_A[40][1] * mat_B[11][2] +
                mat_A[40][2] * mat_B[19][2] +
                mat_A[40][3] * mat_B[27][2] +
                mat_A[41][0] * mat_B[35][2] +
                mat_A[41][1] * mat_B[43][2] +
                mat_A[41][2] * mat_B[51][2] +
                mat_A[41][3] * mat_B[59][2] +
                mat_A[42][0] * mat_B[67][2] +
                mat_A[42][1] * mat_B[75][2] +
                mat_A[42][2] * mat_B[83][2] +
                mat_A[42][3] * mat_B[91][2] +
                mat_A[43][0] * mat_B[99][2] +
                mat_A[43][1] * mat_B[107][2] +
                mat_A[43][2] * mat_B[115][2] +
                mat_A[43][3] * mat_B[123][2] +
                mat_A[44][0] * mat_B[131][2] +
                mat_A[44][1] * mat_B[139][2] +
                mat_A[44][2] * mat_B[147][2] +
                mat_A[44][3] * mat_B[155][2] +
                mat_A[45][0] * mat_B[163][2] +
                mat_A[45][1] * mat_B[171][2] +
                mat_A[45][2] * mat_B[179][2] +
                mat_A[45][3] * mat_B[187][2] +
                mat_A[46][0] * mat_B[195][2] +
                mat_A[46][1] * mat_B[203][2] +
                mat_A[46][2] * mat_B[211][2] +
                mat_A[46][3] * mat_B[219][2] +
                mat_A[47][0] * mat_B[227][2] +
                mat_A[47][1] * mat_B[235][2] +
                mat_A[47][2] * mat_B[243][2] +
                mat_A[47][3] * mat_B[251][2];
    mat_C[43][3] <=
                mat_A[40][0] * mat_B[3][3] +
                mat_A[40][1] * mat_B[11][3] +
                mat_A[40][2] * mat_B[19][3] +
                mat_A[40][3] * mat_B[27][3] +
                mat_A[41][0] * mat_B[35][3] +
                mat_A[41][1] * mat_B[43][3] +
                mat_A[41][2] * mat_B[51][3] +
                mat_A[41][3] * mat_B[59][3] +
                mat_A[42][0] * mat_B[67][3] +
                mat_A[42][1] * mat_B[75][3] +
                mat_A[42][2] * mat_B[83][3] +
                mat_A[42][3] * mat_B[91][3] +
                mat_A[43][0] * mat_B[99][3] +
                mat_A[43][1] * mat_B[107][3] +
                mat_A[43][2] * mat_B[115][3] +
                mat_A[43][3] * mat_B[123][3] +
                mat_A[44][0] * mat_B[131][3] +
                mat_A[44][1] * mat_B[139][3] +
                mat_A[44][2] * mat_B[147][3] +
                mat_A[44][3] * mat_B[155][3] +
                mat_A[45][0] * mat_B[163][3] +
                mat_A[45][1] * mat_B[171][3] +
                mat_A[45][2] * mat_B[179][3] +
                mat_A[45][3] * mat_B[187][3] +
                mat_A[46][0] * mat_B[195][3] +
                mat_A[46][1] * mat_B[203][3] +
                mat_A[46][2] * mat_B[211][3] +
                mat_A[46][3] * mat_B[219][3] +
                mat_A[47][0] * mat_B[227][3] +
                mat_A[47][1] * mat_B[235][3] +
                mat_A[47][2] * mat_B[243][3] +
                mat_A[47][3] * mat_B[251][3];
    mat_C[44][0] <=
                mat_A[40][0] * mat_B[4][0] +
                mat_A[40][1] * mat_B[12][0] +
                mat_A[40][2] * mat_B[20][0] +
                mat_A[40][3] * mat_B[28][0] +
                mat_A[41][0] * mat_B[36][0] +
                mat_A[41][1] * mat_B[44][0] +
                mat_A[41][2] * mat_B[52][0] +
                mat_A[41][3] * mat_B[60][0] +
                mat_A[42][0] * mat_B[68][0] +
                mat_A[42][1] * mat_B[76][0] +
                mat_A[42][2] * mat_B[84][0] +
                mat_A[42][3] * mat_B[92][0] +
                mat_A[43][0] * mat_B[100][0] +
                mat_A[43][1] * mat_B[108][0] +
                mat_A[43][2] * mat_B[116][0] +
                mat_A[43][3] * mat_B[124][0] +
                mat_A[44][0] * mat_B[132][0] +
                mat_A[44][1] * mat_B[140][0] +
                mat_A[44][2] * mat_B[148][0] +
                mat_A[44][3] * mat_B[156][0] +
                mat_A[45][0] * mat_B[164][0] +
                mat_A[45][1] * mat_B[172][0] +
                mat_A[45][2] * mat_B[180][0] +
                mat_A[45][3] * mat_B[188][0] +
                mat_A[46][0] * mat_B[196][0] +
                mat_A[46][1] * mat_B[204][0] +
                mat_A[46][2] * mat_B[212][0] +
                mat_A[46][3] * mat_B[220][0] +
                mat_A[47][0] * mat_B[228][0] +
                mat_A[47][1] * mat_B[236][0] +
                mat_A[47][2] * mat_B[244][0] +
                mat_A[47][3] * mat_B[252][0];
    mat_C[44][1] <=
                mat_A[40][0] * mat_B[4][1] +
                mat_A[40][1] * mat_B[12][1] +
                mat_A[40][2] * mat_B[20][1] +
                mat_A[40][3] * mat_B[28][1] +
                mat_A[41][0] * mat_B[36][1] +
                mat_A[41][1] * mat_B[44][1] +
                mat_A[41][2] * mat_B[52][1] +
                mat_A[41][3] * mat_B[60][1] +
                mat_A[42][0] * mat_B[68][1] +
                mat_A[42][1] * mat_B[76][1] +
                mat_A[42][2] * mat_B[84][1] +
                mat_A[42][3] * mat_B[92][1] +
                mat_A[43][0] * mat_B[100][1] +
                mat_A[43][1] * mat_B[108][1] +
                mat_A[43][2] * mat_B[116][1] +
                mat_A[43][3] * mat_B[124][1] +
                mat_A[44][0] * mat_B[132][1] +
                mat_A[44][1] * mat_B[140][1] +
                mat_A[44][2] * mat_B[148][1] +
                mat_A[44][3] * mat_B[156][1] +
                mat_A[45][0] * mat_B[164][1] +
                mat_A[45][1] * mat_B[172][1] +
                mat_A[45][2] * mat_B[180][1] +
                mat_A[45][3] * mat_B[188][1] +
                mat_A[46][0] * mat_B[196][1] +
                mat_A[46][1] * mat_B[204][1] +
                mat_A[46][2] * mat_B[212][1] +
                mat_A[46][3] * mat_B[220][1] +
                mat_A[47][0] * mat_B[228][1] +
                mat_A[47][1] * mat_B[236][1] +
                mat_A[47][2] * mat_B[244][1] +
                mat_A[47][3] * mat_B[252][1];
    mat_C[44][2] <=
                mat_A[40][0] * mat_B[4][2] +
                mat_A[40][1] * mat_B[12][2] +
                mat_A[40][2] * mat_B[20][2] +
                mat_A[40][3] * mat_B[28][2] +
                mat_A[41][0] * mat_B[36][2] +
                mat_A[41][1] * mat_B[44][2] +
                mat_A[41][2] * mat_B[52][2] +
                mat_A[41][3] * mat_B[60][2] +
                mat_A[42][0] * mat_B[68][2] +
                mat_A[42][1] * mat_B[76][2] +
                mat_A[42][2] * mat_B[84][2] +
                mat_A[42][3] * mat_B[92][2] +
                mat_A[43][0] * mat_B[100][2] +
                mat_A[43][1] * mat_B[108][2] +
                mat_A[43][2] * mat_B[116][2] +
                mat_A[43][3] * mat_B[124][2] +
                mat_A[44][0] * mat_B[132][2] +
                mat_A[44][1] * mat_B[140][2] +
                mat_A[44][2] * mat_B[148][2] +
                mat_A[44][3] * mat_B[156][2] +
                mat_A[45][0] * mat_B[164][2] +
                mat_A[45][1] * mat_B[172][2] +
                mat_A[45][2] * mat_B[180][2] +
                mat_A[45][3] * mat_B[188][2] +
                mat_A[46][0] * mat_B[196][2] +
                mat_A[46][1] * mat_B[204][2] +
                mat_A[46][2] * mat_B[212][2] +
                mat_A[46][3] * mat_B[220][2] +
                mat_A[47][0] * mat_B[228][2] +
                mat_A[47][1] * mat_B[236][2] +
                mat_A[47][2] * mat_B[244][2] +
                mat_A[47][3] * mat_B[252][2];
    mat_C[44][3] <=
                mat_A[40][0] * mat_B[4][3] +
                mat_A[40][1] * mat_B[12][3] +
                mat_A[40][2] * mat_B[20][3] +
                mat_A[40][3] * mat_B[28][3] +
                mat_A[41][0] * mat_B[36][3] +
                mat_A[41][1] * mat_B[44][3] +
                mat_A[41][2] * mat_B[52][3] +
                mat_A[41][3] * mat_B[60][3] +
                mat_A[42][0] * mat_B[68][3] +
                mat_A[42][1] * mat_B[76][3] +
                mat_A[42][2] * mat_B[84][3] +
                mat_A[42][3] * mat_B[92][3] +
                mat_A[43][0] * mat_B[100][3] +
                mat_A[43][1] * mat_B[108][3] +
                mat_A[43][2] * mat_B[116][3] +
                mat_A[43][3] * mat_B[124][3] +
                mat_A[44][0] * mat_B[132][3] +
                mat_A[44][1] * mat_B[140][3] +
                mat_A[44][2] * mat_B[148][3] +
                mat_A[44][3] * mat_B[156][3] +
                mat_A[45][0] * mat_B[164][3] +
                mat_A[45][1] * mat_B[172][3] +
                mat_A[45][2] * mat_B[180][3] +
                mat_A[45][3] * mat_B[188][3] +
                mat_A[46][0] * mat_B[196][3] +
                mat_A[46][1] * mat_B[204][3] +
                mat_A[46][2] * mat_B[212][3] +
                mat_A[46][3] * mat_B[220][3] +
                mat_A[47][0] * mat_B[228][3] +
                mat_A[47][1] * mat_B[236][3] +
                mat_A[47][2] * mat_B[244][3] +
                mat_A[47][3] * mat_B[252][3];
    mat_C[45][0] <=
                mat_A[40][0] * mat_B[5][0] +
                mat_A[40][1] * mat_B[13][0] +
                mat_A[40][2] * mat_B[21][0] +
                mat_A[40][3] * mat_B[29][0] +
                mat_A[41][0] * mat_B[37][0] +
                mat_A[41][1] * mat_B[45][0] +
                mat_A[41][2] * mat_B[53][0] +
                mat_A[41][3] * mat_B[61][0] +
                mat_A[42][0] * mat_B[69][0] +
                mat_A[42][1] * mat_B[77][0] +
                mat_A[42][2] * mat_B[85][0] +
                mat_A[42][3] * mat_B[93][0] +
                mat_A[43][0] * mat_B[101][0] +
                mat_A[43][1] * mat_B[109][0] +
                mat_A[43][2] * mat_B[117][0] +
                mat_A[43][3] * mat_B[125][0] +
                mat_A[44][0] * mat_B[133][0] +
                mat_A[44][1] * mat_B[141][0] +
                mat_A[44][2] * mat_B[149][0] +
                mat_A[44][3] * mat_B[157][0] +
                mat_A[45][0] * mat_B[165][0] +
                mat_A[45][1] * mat_B[173][0] +
                mat_A[45][2] * mat_B[181][0] +
                mat_A[45][3] * mat_B[189][0] +
                mat_A[46][0] * mat_B[197][0] +
                mat_A[46][1] * mat_B[205][0] +
                mat_A[46][2] * mat_B[213][0] +
                mat_A[46][3] * mat_B[221][0] +
                mat_A[47][0] * mat_B[229][0] +
                mat_A[47][1] * mat_B[237][0] +
                mat_A[47][2] * mat_B[245][0] +
                mat_A[47][3] * mat_B[253][0];
    mat_C[45][1] <=
                mat_A[40][0] * mat_B[5][1] +
                mat_A[40][1] * mat_B[13][1] +
                mat_A[40][2] * mat_B[21][1] +
                mat_A[40][3] * mat_B[29][1] +
                mat_A[41][0] * mat_B[37][1] +
                mat_A[41][1] * mat_B[45][1] +
                mat_A[41][2] * mat_B[53][1] +
                mat_A[41][3] * mat_B[61][1] +
                mat_A[42][0] * mat_B[69][1] +
                mat_A[42][1] * mat_B[77][1] +
                mat_A[42][2] * mat_B[85][1] +
                mat_A[42][3] * mat_B[93][1] +
                mat_A[43][0] * mat_B[101][1] +
                mat_A[43][1] * mat_B[109][1] +
                mat_A[43][2] * mat_B[117][1] +
                mat_A[43][3] * mat_B[125][1] +
                mat_A[44][0] * mat_B[133][1] +
                mat_A[44][1] * mat_B[141][1] +
                mat_A[44][2] * mat_B[149][1] +
                mat_A[44][3] * mat_B[157][1] +
                mat_A[45][0] * mat_B[165][1] +
                mat_A[45][1] * mat_B[173][1] +
                mat_A[45][2] * mat_B[181][1] +
                mat_A[45][3] * mat_B[189][1] +
                mat_A[46][0] * mat_B[197][1] +
                mat_A[46][1] * mat_B[205][1] +
                mat_A[46][2] * mat_B[213][1] +
                mat_A[46][3] * mat_B[221][1] +
                mat_A[47][0] * mat_B[229][1] +
                mat_A[47][1] * mat_B[237][1] +
                mat_A[47][2] * mat_B[245][1] +
                mat_A[47][3] * mat_B[253][1];
    mat_C[45][2] <=
                mat_A[40][0] * mat_B[5][2] +
                mat_A[40][1] * mat_B[13][2] +
                mat_A[40][2] * mat_B[21][2] +
                mat_A[40][3] * mat_B[29][2] +
                mat_A[41][0] * mat_B[37][2] +
                mat_A[41][1] * mat_B[45][2] +
                mat_A[41][2] * mat_B[53][2] +
                mat_A[41][3] * mat_B[61][2] +
                mat_A[42][0] * mat_B[69][2] +
                mat_A[42][1] * mat_B[77][2] +
                mat_A[42][2] * mat_B[85][2] +
                mat_A[42][3] * mat_B[93][2] +
                mat_A[43][0] * mat_B[101][2] +
                mat_A[43][1] * mat_B[109][2] +
                mat_A[43][2] * mat_B[117][2] +
                mat_A[43][3] * mat_B[125][2] +
                mat_A[44][0] * mat_B[133][2] +
                mat_A[44][1] * mat_B[141][2] +
                mat_A[44][2] * mat_B[149][2] +
                mat_A[44][3] * mat_B[157][2] +
                mat_A[45][0] * mat_B[165][2] +
                mat_A[45][1] * mat_B[173][2] +
                mat_A[45][2] * mat_B[181][2] +
                mat_A[45][3] * mat_B[189][2] +
                mat_A[46][0] * mat_B[197][2] +
                mat_A[46][1] * mat_B[205][2] +
                mat_A[46][2] * mat_B[213][2] +
                mat_A[46][3] * mat_B[221][2] +
                mat_A[47][0] * mat_B[229][2] +
                mat_A[47][1] * mat_B[237][2] +
                mat_A[47][2] * mat_B[245][2] +
                mat_A[47][3] * mat_B[253][2];
    mat_C[45][3] <=
                mat_A[40][0] * mat_B[5][3] +
                mat_A[40][1] * mat_B[13][3] +
                mat_A[40][2] * mat_B[21][3] +
                mat_A[40][3] * mat_B[29][3] +
                mat_A[41][0] * mat_B[37][3] +
                mat_A[41][1] * mat_B[45][3] +
                mat_A[41][2] * mat_B[53][3] +
                mat_A[41][3] * mat_B[61][3] +
                mat_A[42][0] * mat_B[69][3] +
                mat_A[42][1] * mat_B[77][3] +
                mat_A[42][2] * mat_B[85][3] +
                mat_A[42][3] * mat_B[93][3] +
                mat_A[43][0] * mat_B[101][3] +
                mat_A[43][1] * mat_B[109][3] +
                mat_A[43][2] * mat_B[117][3] +
                mat_A[43][3] * mat_B[125][3] +
                mat_A[44][0] * mat_B[133][3] +
                mat_A[44][1] * mat_B[141][3] +
                mat_A[44][2] * mat_B[149][3] +
                mat_A[44][3] * mat_B[157][3] +
                mat_A[45][0] * mat_B[165][3] +
                mat_A[45][1] * mat_B[173][3] +
                mat_A[45][2] * mat_B[181][3] +
                mat_A[45][3] * mat_B[189][3] +
                mat_A[46][0] * mat_B[197][3] +
                mat_A[46][1] * mat_B[205][3] +
                mat_A[46][2] * mat_B[213][3] +
                mat_A[46][3] * mat_B[221][3] +
                mat_A[47][0] * mat_B[229][3] +
                mat_A[47][1] * mat_B[237][3] +
                mat_A[47][2] * mat_B[245][3] +
                mat_A[47][3] * mat_B[253][3];
    mat_C[46][0] <=
                mat_A[40][0] * mat_B[6][0] +
                mat_A[40][1] * mat_B[14][0] +
                mat_A[40][2] * mat_B[22][0] +
                mat_A[40][3] * mat_B[30][0] +
                mat_A[41][0] * mat_B[38][0] +
                mat_A[41][1] * mat_B[46][0] +
                mat_A[41][2] * mat_B[54][0] +
                mat_A[41][3] * mat_B[62][0] +
                mat_A[42][0] * mat_B[70][0] +
                mat_A[42][1] * mat_B[78][0] +
                mat_A[42][2] * mat_B[86][0] +
                mat_A[42][3] * mat_B[94][0] +
                mat_A[43][0] * mat_B[102][0] +
                mat_A[43][1] * mat_B[110][0] +
                mat_A[43][2] * mat_B[118][0] +
                mat_A[43][3] * mat_B[126][0] +
                mat_A[44][0] * mat_B[134][0] +
                mat_A[44][1] * mat_B[142][0] +
                mat_A[44][2] * mat_B[150][0] +
                mat_A[44][3] * mat_B[158][0] +
                mat_A[45][0] * mat_B[166][0] +
                mat_A[45][1] * mat_B[174][0] +
                mat_A[45][2] * mat_B[182][0] +
                mat_A[45][3] * mat_B[190][0] +
                mat_A[46][0] * mat_B[198][0] +
                mat_A[46][1] * mat_B[206][0] +
                mat_A[46][2] * mat_B[214][0] +
                mat_A[46][3] * mat_B[222][0] +
                mat_A[47][0] * mat_B[230][0] +
                mat_A[47][1] * mat_B[238][0] +
                mat_A[47][2] * mat_B[246][0] +
                mat_A[47][3] * mat_B[254][0];
    mat_C[46][1] <=
                mat_A[40][0] * mat_B[6][1] +
                mat_A[40][1] * mat_B[14][1] +
                mat_A[40][2] * mat_B[22][1] +
                mat_A[40][3] * mat_B[30][1] +
                mat_A[41][0] * mat_B[38][1] +
                mat_A[41][1] * mat_B[46][1] +
                mat_A[41][2] * mat_B[54][1] +
                mat_A[41][3] * mat_B[62][1] +
                mat_A[42][0] * mat_B[70][1] +
                mat_A[42][1] * mat_B[78][1] +
                mat_A[42][2] * mat_B[86][1] +
                mat_A[42][3] * mat_B[94][1] +
                mat_A[43][0] * mat_B[102][1] +
                mat_A[43][1] * mat_B[110][1] +
                mat_A[43][2] * mat_B[118][1] +
                mat_A[43][3] * mat_B[126][1] +
                mat_A[44][0] * mat_B[134][1] +
                mat_A[44][1] * mat_B[142][1] +
                mat_A[44][2] * mat_B[150][1] +
                mat_A[44][3] * mat_B[158][1] +
                mat_A[45][0] * mat_B[166][1] +
                mat_A[45][1] * mat_B[174][1] +
                mat_A[45][2] * mat_B[182][1] +
                mat_A[45][3] * mat_B[190][1] +
                mat_A[46][0] * mat_B[198][1] +
                mat_A[46][1] * mat_B[206][1] +
                mat_A[46][2] * mat_B[214][1] +
                mat_A[46][3] * mat_B[222][1] +
                mat_A[47][0] * mat_B[230][1] +
                mat_A[47][1] * mat_B[238][1] +
                mat_A[47][2] * mat_B[246][1] +
                mat_A[47][3] * mat_B[254][1];
    mat_C[46][2] <=
                mat_A[40][0] * mat_B[6][2] +
                mat_A[40][1] * mat_B[14][2] +
                mat_A[40][2] * mat_B[22][2] +
                mat_A[40][3] * mat_B[30][2] +
                mat_A[41][0] * mat_B[38][2] +
                mat_A[41][1] * mat_B[46][2] +
                mat_A[41][2] * mat_B[54][2] +
                mat_A[41][3] * mat_B[62][2] +
                mat_A[42][0] * mat_B[70][2] +
                mat_A[42][1] * mat_B[78][2] +
                mat_A[42][2] * mat_B[86][2] +
                mat_A[42][3] * mat_B[94][2] +
                mat_A[43][0] * mat_B[102][2] +
                mat_A[43][1] * mat_B[110][2] +
                mat_A[43][2] * mat_B[118][2] +
                mat_A[43][3] * mat_B[126][2] +
                mat_A[44][0] * mat_B[134][2] +
                mat_A[44][1] * mat_B[142][2] +
                mat_A[44][2] * mat_B[150][2] +
                mat_A[44][3] * mat_B[158][2] +
                mat_A[45][0] * mat_B[166][2] +
                mat_A[45][1] * mat_B[174][2] +
                mat_A[45][2] * mat_B[182][2] +
                mat_A[45][3] * mat_B[190][2] +
                mat_A[46][0] * mat_B[198][2] +
                mat_A[46][1] * mat_B[206][2] +
                mat_A[46][2] * mat_B[214][2] +
                mat_A[46][3] * mat_B[222][2] +
                mat_A[47][0] * mat_B[230][2] +
                mat_A[47][1] * mat_B[238][2] +
                mat_A[47][2] * mat_B[246][2] +
                mat_A[47][3] * mat_B[254][2];
    mat_C[46][3] <=
                mat_A[40][0] * mat_B[6][3] +
                mat_A[40][1] * mat_B[14][3] +
                mat_A[40][2] * mat_B[22][3] +
                mat_A[40][3] * mat_B[30][3] +
                mat_A[41][0] * mat_B[38][3] +
                mat_A[41][1] * mat_B[46][3] +
                mat_A[41][2] * mat_B[54][3] +
                mat_A[41][3] * mat_B[62][3] +
                mat_A[42][0] * mat_B[70][3] +
                mat_A[42][1] * mat_B[78][3] +
                mat_A[42][2] * mat_B[86][3] +
                mat_A[42][3] * mat_B[94][3] +
                mat_A[43][0] * mat_B[102][3] +
                mat_A[43][1] * mat_B[110][3] +
                mat_A[43][2] * mat_B[118][3] +
                mat_A[43][3] * mat_B[126][3] +
                mat_A[44][0] * mat_B[134][3] +
                mat_A[44][1] * mat_B[142][3] +
                mat_A[44][2] * mat_B[150][3] +
                mat_A[44][3] * mat_B[158][3] +
                mat_A[45][0] * mat_B[166][3] +
                mat_A[45][1] * mat_B[174][3] +
                mat_A[45][2] * mat_B[182][3] +
                mat_A[45][3] * mat_B[190][3] +
                mat_A[46][0] * mat_B[198][3] +
                mat_A[46][1] * mat_B[206][3] +
                mat_A[46][2] * mat_B[214][3] +
                mat_A[46][3] * mat_B[222][3] +
                mat_A[47][0] * mat_B[230][3] +
                mat_A[47][1] * mat_B[238][3] +
                mat_A[47][2] * mat_B[246][3] +
                mat_A[47][3] * mat_B[254][3];
    mat_C[47][0] <=
                mat_A[40][0] * mat_B[7][0] +
                mat_A[40][1] * mat_B[15][0] +
                mat_A[40][2] * mat_B[23][0] +
                mat_A[40][3] * mat_B[31][0] +
                mat_A[41][0] * mat_B[39][0] +
                mat_A[41][1] * mat_B[47][0] +
                mat_A[41][2] * mat_B[55][0] +
                mat_A[41][3] * mat_B[63][0] +
                mat_A[42][0] * mat_B[71][0] +
                mat_A[42][1] * mat_B[79][0] +
                mat_A[42][2] * mat_B[87][0] +
                mat_A[42][3] * mat_B[95][0] +
                mat_A[43][0] * mat_B[103][0] +
                mat_A[43][1] * mat_B[111][0] +
                mat_A[43][2] * mat_B[119][0] +
                mat_A[43][3] * mat_B[127][0] +
                mat_A[44][0] * mat_B[135][0] +
                mat_A[44][1] * mat_B[143][0] +
                mat_A[44][2] * mat_B[151][0] +
                mat_A[44][3] * mat_B[159][0] +
                mat_A[45][0] * mat_B[167][0] +
                mat_A[45][1] * mat_B[175][0] +
                mat_A[45][2] * mat_B[183][0] +
                mat_A[45][3] * mat_B[191][0] +
                mat_A[46][0] * mat_B[199][0] +
                mat_A[46][1] * mat_B[207][0] +
                mat_A[46][2] * mat_B[215][0] +
                mat_A[46][3] * mat_B[223][0] +
                mat_A[47][0] * mat_B[231][0] +
                mat_A[47][1] * mat_B[239][0] +
                mat_A[47][2] * mat_B[247][0] +
                mat_A[47][3] * mat_B[255][0];
    mat_C[47][1] <=
                mat_A[40][0] * mat_B[7][1] +
                mat_A[40][1] * mat_B[15][1] +
                mat_A[40][2] * mat_B[23][1] +
                mat_A[40][3] * mat_B[31][1] +
                mat_A[41][0] * mat_B[39][1] +
                mat_A[41][1] * mat_B[47][1] +
                mat_A[41][2] * mat_B[55][1] +
                mat_A[41][3] * mat_B[63][1] +
                mat_A[42][0] * mat_B[71][1] +
                mat_A[42][1] * mat_B[79][1] +
                mat_A[42][2] * mat_B[87][1] +
                mat_A[42][3] * mat_B[95][1] +
                mat_A[43][0] * mat_B[103][1] +
                mat_A[43][1] * mat_B[111][1] +
                mat_A[43][2] * mat_B[119][1] +
                mat_A[43][3] * mat_B[127][1] +
                mat_A[44][0] * mat_B[135][1] +
                mat_A[44][1] * mat_B[143][1] +
                mat_A[44][2] * mat_B[151][1] +
                mat_A[44][3] * mat_B[159][1] +
                mat_A[45][0] * mat_B[167][1] +
                mat_A[45][1] * mat_B[175][1] +
                mat_A[45][2] * mat_B[183][1] +
                mat_A[45][3] * mat_B[191][1] +
                mat_A[46][0] * mat_B[199][1] +
                mat_A[46][1] * mat_B[207][1] +
                mat_A[46][2] * mat_B[215][1] +
                mat_A[46][3] * mat_B[223][1] +
                mat_A[47][0] * mat_B[231][1] +
                mat_A[47][1] * mat_B[239][1] +
                mat_A[47][2] * mat_B[247][1] +
                mat_A[47][3] * mat_B[255][1];
    mat_C[47][2] <=
                mat_A[40][0] * mat_B[7][2] +
                mat_A[40][1] * mat_B[15][2] +
                mat_A[40][2] * mat_B[23][2] +
                mat_A[40][3] * mat_B[31][2] +
                mat_A[41][0] * mat_B[39][2] +
                mat_A[41][1] * mat_B[47][2] +
                mat_A[41][2] * mat_B[55][2] +
                mat_A[41][3] * mat_B[63][2] +
                mat_A[42][0] * mat_B[71][2] +
                mat_A[42][1] * mat_B[79][2] +
                mat_A[42][2] * mat_B[87][2] +
                mat_A[42][3] * mat_B[95][2] +
                mat_A[43][0] * mat_B[103][2] +
                mat_A[43][1] * mat_B[111][2] +
                mat_A[43][2] * mat_B[119][2] +
                mat_A[43][3] * mat_B[127][2] +
                mat_A[44][0] * mat_B[135][2] +
                mat_A[44][1] * mat_B[143][2] +
                mat_A[44][2] * mat_B[151][2] +
                mat_A[44][3] * mat_B[159][2] +
                mat_A[45][0] * mat_B[167][2] +
                mat_A[45][1] * mat_B[175][2] +
                mat_A[45][2] * mat_B[183][2] +
                mat_A[45][3] * mat_B[191][2] +
                mat_A[46][0] * mat_B[199][2] +
                mat_A[46][1] * mat_B[207][2] +
                mat_A[46][2] * mat_B[215][2] +
                mat_A[46][3] * mat_B[223][2] +
                mat_A[47][0] * mat_B[231][2] +
                mat_A[47][1] * mat_B[239][2] +
                mat_A[47][2] * mat_B[247][2] +
                mat_A[47][3] * mat_B[255][2];
    mat_C[47][3] <=
                mat_A[40][0] * mat_B[7][3] +
                mat_A[40][1] * mat_B[15][3] +
                mat_A[40][2] * mat_B[23][3] +
                mat_A[40][3] * mat_B[31][3] +
                mat_A[41][0] * mat_B[39][3] +
                mat_A[41][1] * mat_B[47][3] +
                mat_A[41][2] * mat_B[55][3] +
                mat_A[41][3] * mat_B[63][3] +
                mat_A[42][0] * mat_B[71][3] +
                mat_A[42][1] * mat_B[79][3] +
                mat_A[42][2] * mat_B[87][3] +
                mat_A[42][3] * mat_B[95][3] +
                mat_A[43][0] * mat_B[103][3] +
                mat_A[43][1] * mat_B[111][3] +
                mat_A[43][2] * mat_B[119][3] +
                mat_A[43][3] * mat_B[127][3] +
                mat_A[44][0] * mat_B[135][3] +
                mat_A[44][1] * mat_B[143][3] +
                mat_A[44][2] * mat_B[151][3] +
                mat_A[44][3] * mat_B[159][3] +
                mat_A[45][0] * mat_B[167][3] +
                mat_A[45][1] * mat_B[175][3] +
                mat_A[45][2] * mat_B[183][3] +
                mat_A[45][3] * mat_B[191][3] +
                mat_A[46][0] * mat_B[199][3] +
                mat_A[46][1] * mat_B[207][3] +
                mat_A[46][2] * mat_B[215][3] +
                mat_A[46][3] * mat_B[223][3] +
                mat_A[47][0] * mat_B[231][3] +
                mat_A[47][1] * mat_B[239][3] +
                mat_A[47][2] * mat_B[247][3] +
                mat_A[47][3] * mat_B[255][3];
    mat_C[48][0] <=
                mat_A[48][0] * mat_B[0][0] +
                mat_A[48][1] * mat_B[8][0] +
                mat_A[48][2] * mat_B[16][0] +
                mat_A[48][3] * mat_B[24][0] +
                mat_A[49][0] * mat_B[32][0] +
                mat_A[49][1] * mat_B[40][0] +
                mat_A[49][2] * mat_B[48][0] +
                mat_A[49][3] * mat_B[56][0] +
                mat_A[50][0] * mat_B[64][0] +
                mat_A[50][1] * mat_B[72][0] +
                mat_A[50][2] * mat_B[80][0] +
                mat_A[50][3] * mat_B[88][0] +
                mat_A[51][0] * mat_B[96][0] +
                mat_A[51][1] * mat_B[104][0] +
                mat_A[51][2] * mat_B[112][0] +
                mat_A[51][3] * mat_B[120][0] +
                mat_A[52][0] * mat_B[128][0] +
                mat_A[52][1] * mat_B[136][0] +
                mat_A[52][2] * mat_B[144][0] +
                mat_A[52][3] * mat_B[152][0] +
                mat_A[53][0] * mat_B[160][0] +
                mat_A[53][1] * mat_B[168][0] +
                mat_A[53][2] * mat_B[176][0] +
                mat_A[53][3] * mat_B[184][0] +
                mat_A[54][0] * mat_B[192][0] +
                mat_A[54][1] * mat_B[200][0] +
                mat_A[54][2] * mat_B[208][0] +
                mat_A[54][3] * mat_B[216][0] +
                mat_A[55][0] * mat_B[224][0] +
                mat_A[55][1] * mat_B[232][0] +
                mat_A[55][2] * mat_B[240][0] +
                mat_A[55][3] * mat_B[248][0];
    mat_C[48][1] <=
                mat_A[48][0] * mat_B[0][1] +
                mat_A[48][1] * mat_B[8][1] +
                mat_A[48][2] * mat_B[16][1] +
                mat_A[48][3] * mat_B[24][1] +
                mat_A[49][0] * mat_B[32][1] +
                mat_A[49][1] * mat_B[40][1] +
                mat_A[49][2] * mat_B[48][1] +
                mat_A[49][3] * mat_B[56][1] +
                mat_A[50][0] * mat_B[64][1] +
                mat_A[50][1] * mat_B[72][1] +
                mat_A[50][2] * mat_B[80][1] +
                mat_A[50][3] * mat_B[88][1] +
                mat_A[51][0] * mat_B[96][1] +
                mat_A[51][1] * mat_B[104][1] +
                mat_A[51][2] * mat_B[112][1] +
                mat_A[51][3] * mat_B[120][1] +
                mat_A[52][0] * mat_B[128][1] +
                mat_A[52][1] * mat_B[136][1] +
                mat_A[52][2] * mat_B[144][1] +
                mat_A[52][3] * mat_B[152][1] +
                mat_A[53][0] * mat_B[160][1] +
                mat_A[53][1] * mat_B[168][1] +
                mat_A[53][2] * mat_B[176][1] +
                mat_A[53][3] * mat_B[184][1] +
                mat_A[54][0] * mat_B[192][1] +
                mat_A[54][1] * mat_B[200][1] +
                mat_A[54][2] * mat_B[208][1] +
                mat_A[54][3] * mat_B[216][1] +
                mat_A[55][0] * mat_B[224][1] +
                mat_A[55][1] * mat_B[232][1] +
                mat_A[55][2] * mat_B[240][1] +
                mat_A[55][3] * mat_B[248][1];
    mat_C[48][2] <=
                mat_A[48][0] * mat_B[0][2] +
                mat_A[48][1] * mat_B[8][2] +
                mat_A[48][2] * mat_B[16][2] +
                mat_A[48][3] * mat_B[24][2] +
                mat_A[49][0] * mat_B[32][2] +
                mat_A[49][1] * mat_B[40][2] +
                mat_A[49][2] * mat_B[48][2] +
                mat_A[49][3] * mat_B[56][2] +
                mat_A[50][0] * mat_B[64][2] +
                mat_A[50][1] * mat_B[72][2] +
                mat_A[50][2] * mat_B[80][2] +
                mat_A[50][3] * mat_B[88][2] +
                mat_A[51][0] * mat_B[96][2] +
                mat_A[51][1] * mat_B[104][2] +
                mat_A[51][2] * mat_B[112][2] +
                mat_A[51][3] * mat_B[120][2] +
                mat_A[52][0] * mat_B[128][2] +
                mat_A[52][1] * mat_B[136][2] +
                mat_A[52][2] * mat_B[144][2] +
                mat_A[52][3] * mat_B[152][2] +
                mat_A[53][0] * mat_B[160][2] +
                mat_A[53][1] * mat_B[168][2] +
                mat_A[53][2] * mat_B[176][2] +
                mat_A[53][3] * mat_B[184][2] +
                mat_A[54][0] * mat_B[192][2] +
                mat_A[54][1] * mat_B[200][2] +
                mat_A[54][2] * mat_B[208][2] +
                mat_A[54][3] * mat_B[216][2] +
                mat_A[55][0] * mat_B[224][2] +
                mat_A[55][1] * mat_B[232][2] +
                mat_A[55][2] * mat_B[240][2] +
                mat_A[55][3] * mat_B[248][2];
    mat_C[48][3] <=
                mat_A[48][0] * mat_B[0][3] +
                mat_A[48][1] * mat_B[8][3] +
                mat_A[48][2] * mat_B[16][3] +
                mat_A[48][3] * mat_B[24][3] +
                mat_A[49][0] * mat_B[32][3] +
                mat_A[49][1] * mat_B[40][3] +
                mat_A[49][2] * mat_B[48][3] +
                mat_A[49][3] * mat_B[56][3] +
                mat_A[50][0] * mat_B[64][3] +
                mat_A[50][1] * mat_B[72][3] +
                mat_A[50][2] * mat_B[80][3] +
                mat_A[50][3] * mat_B[88][3] +
                mat_A[51][0] * mat_B[96][3] +
                mat_A[51][1] * mat_B[104][3] +
                mat_A[51][2] * mat_B[112][3] +
                mat_A[51][3] * mat_B[120][3] +
                mat_A[52][0] * mat_B[128][3] +
                mat_A[52][1] * mat_B[136][3] +
                mat_A[52][2] * mat_B[144][3] +
                mat_A[52][3] * mat_B[152][3] +
                mat_A[53][0] * mat_B[160][3] +
                mat_A[53][1] * mat_B[168][3] +
                mat_A[53][2] * mat_B[176][3] +
                mat_A[53][3] * mat_B[184][3] +
                mat_A[54][0] * mat_B[192][3] +
                mat_A[54][1] * mat_B[200][3] +
                mat_A[54][2] * mat_B[208][3] +
                mat_A[54][3] * mat_B[216][3] +
                mat_A[55][0] * mat_B[224][3] +
                mat_A[55][1] * mat_B[232][3] +
                mat_A[55][2] * mat_B[240][3] +
                mat_A[55][3] * mat_B[248][3];
    mat_C[49][0] <=
                mat_A[48][0] * mat_B[1][0] +
                mat_A[48][1] * mat_B[9][0] +
                mat_A[48][2] * mat_B[17][0] +
                mat_A[48][3] * mat_B[25][0] +
                mat_A[49][0] * mat_B[33][0] +
                mat_A[49][1] * mat_B[41][0] +
                mat_A[49][2] * mat_B[49][0] +
                mat_A[49][3] * mat_B[57][0] +
                mat_A[50][0] * mat_B[65][0] +
                mat_A[50][1] * mat_B[73][0] +
                mat_A[50][2] * mat_B[81][0] +
                mat_A[50][3] * mat_B[89][0] +
                mat_A[51][0] * mat_B[97][0] +
                mat_A[51][1] * mat_B[105][0] +
                mat_A[51][2] * mat_B[113][0] +
                mat_A[51][3] * mat_B[121][0] +
                mat_A[52][0] * mat_B[129][0] +
                mat_A[52][1] * mat_B[137][0] +
                mat_A[52][2] * mat_B[145][0] +
                mat_A[52][3] * mat_B[153][0] +
                mat_A[53][0] * mat_B[161][0] +
                mat_A[53][1] * mat_B[169][0] +
                mat_A[53][2] * mat_B[177][0] +
                mat_A[53][3] * mat_B[185][0] +
                mat_A[54][0] * mat_B[193][0] +
                mat_A[54][1] * mat_B[201][0] +
                mat_A[54][2] * mat_B[209][0] +
                mat_A[54][3] * mat_B[217][0] +
                mat_A[55][0] * mat_B[225][0] +
                mat_A[55][1] * mat_B[233][0] +
                mat_A[55][2] * mat_B[241][0] +
                mat_A[55][3] * mat_B[249][0];
    mat_C[49][1] <=
                mat_A[48][0] * mat_B[1][1] +
                mat_A[48][1] * mat_B[9][1] +
                mat_A[48][2] * mat_B[17][1] +
                mat_A[48][3] * mat_B[25][1] +
                mat_A[49][0] * mat_B[33][1] +
                mat_A[49][1] * mat_B[41][1] +
                mat_A[49][2] * mat_B[49][1] +
                mat_A[49][3] * mat_B[57][1] +
                mat_A[50][0] * mat_B[65][1] +
                mat_A[50][1] * mat_B[73][1] +
                mat_A[50][2] * mat_B[81][1] +
                mat_A[50][3] * mat_B[89][1] +
                mat_A[51][0] * mat_B[97][1] +
                mat_A[51][1] * mat_B[105][1] +
                mat_A[51][2] * mat_B[113][1] +
                mat_A[51][3] * mat_B[121][1] +
                mat_A[52][0] * mat_B[129][1] +
                mat_A[52][1] * mat_B[137][1] +
                mat_A[52][2] * mat_B[145][1] +
                mat_A[52][3] * mat_B[153][1] +
                mat_A[53][0] * mat_B[161][1] +
                mat_A[53][1] * mat_B[169][1] +
                mat_A[53][2] * mat_B[177][1] +
                mat_A[53][3] * mat_B[185][1] +
                mat_A[54][0] * mat_B[193][1] +
                mat_A[54][1] * mat_B[201][1] +
                mat_A[54][2] * mat_B[209][1] +
                mat_A[54][3] * mat_B[217][1] +
                mat_A[55][0] * mat_B[225][1] +
                mat_A[55][1] * mat_B[233][1] +
                mat_A[55][2] * mat_B[241][1] +
                mat_A[55][3] * mat_B[249][1];
    mat_C[49][2] <=
                mat_A[48][0] * mat_B[1][2] +
                mat_A[48][1] * mat_B[9][2] +
                mat_A[48][2] * mat_B[17][2] +
                mat_A[48][3] * mat_B[25][2] +
                mat_A[49][0] * mat_B[33][2] +
                mat_A[49][1] * mat_B[41][2] +
                mat_A[49][2] * mat_B[49][2] +
                mat_A[49][3] * mat_B[57][2] +
                mat_A[50][0] * mat_B[65][2] +
                mat_A[50][1] * mat_B[73][2] +
                mat_A[50][2] * mat_B[81][2] +
                mat_A[50][3] * mat_B[89][2] +
                mat_A[51][0] * mat_B[97][2] +
                mat_A[51][1] * mat_B[105][2] +
                mat_A[51][2] * mat_B[113][2] +
                mat_A[51][3] * mat_B[121][2] +
                mat_A[52][0] * mat_B[129][2] +
                mat_A[52][1] * mat_B[137][2] +
                mat_A[52][2] * mat_B[145][2] +
                mat_A[52][3] * mat_B[153][2] +
                mat_A[53][0] * mat_B[161][2] +
                mat_A[53][1] * mat_B[169][2] +
                mat_A[53][2] * mat_B[177][2] +
                mat_A[53][3] * mat_B[185][2] +
                mat_A[54][0] * mat_B[193][2] +
                mat_A[54][1] * mat_B[201][2] +
                mat_A[54][2] * mat_B[209][2] +
                mat_A[54][3] * mat_B[217][2] +
                mat_A[55][0] * mat_B[225][2] +
                mat_A[55][1] * mat_B[233][2] +
                mat_A[55][2] * mat_B[241][2] +
                mat_A[55][3] * mat_B[249][2];
    mat_C[49][3] <=
                mat_A[48][0] * mat_B[1][3] +
                mat_A[48][1] * mat_B[9][3] +
                mat_A[48][2] * mat_B[17][3] +
                mat_A[48][3] * mat_B[25][3] +
                mat_A[49][0] * mat_B[33][3] +
                mat_A[49][1] * mat_B[41][3] +
                mat_A[49][2] * mat_B[49][3] +
                mat_A[49][3] * mat_B[57][3] +
                mat_A[50][0] * mat_B[65][3] +
                mat_A[50][1] * mat_B[73][3] +
                mat_A[50][2] * mat_B[81][3] +
                mat_A[50][3] * mat_B[89][3] +
                mat_A[51][0] * mat_B[97][3] +
                mat_A[51][1] * mat_B[105][3] +
                mat_A[51][2] * mat_B[113][3] +
                mat_A[51][3] * mat_B[121][3] +
                mat_A[52][0] * mat_B[129][3] +
                mat_A[52][1] * mat_B[137][3] +
                mat_A[52][2] * mat_B[145][3] +
                mat_A[52][3] * mat_B[153][3] +
                mat_A[53][0] * mat_B[161][3] +
                mat_A[53][1] * mat_B[169][3] +
                mat_A[53][2] * mat_B[177][3] +
                mat_A[53][3] * mat_B[185][3] +
                mat_A[54][0] * mat_B[193][3] +
                mat_A[54][1] * mat_B[201][3] +
                mat_A[54][2] * mat_B[209][3] +
                mat_A[54][3] * mat_B[217][3] +
                mat_A[55][0] * mat_B[225][3] +
                mat_A[55][1] * mat_B[233][3] +
                mat_A[55][2] * mat_B[241][3] +
                mat_A[55][3] * mat_B[249][3];
    mat_C[50][0] <=
                mat_A[48][0] * mat_B[2][0] +
                mat_A[48][1] * mat_B[10][0] +
                mat_A[48][2] * mat_B[18][0] +
                mat_A[48][3] * mat_B[26][0] +
                mat_A[49][0] * mat_B[34][0] +
                mat_A[49][1] * mat_B[42][0] +
                mat_A[49][2] * mat_B[50][0] +
                mat_A[49][3] * mat_B[58][0] +
                mat_A[50][0] * mat_B[66][0] +
                mat_A[50][1] * mat_B[74][0] +
                mat_A[50][2] * mat_B[82][0] +
                mat_A[50][3] * mat_B[90][0] +
                mat_A[51][0] * mat_B[98][0] +
                mat_A[51][1] * mat_B[106][0] +
                mat_A[51][2] * mat_B[114][0] +
                mat_A[51][3] * mat_B[122][0] +
                mat_A[52][0] * mat_B[130][0] +
                mat_A[52][1] * mat_B[138][0] +
                mat_A[52][2] * mat_B[146][0] +
                mat_A[52][3] * mat_B[154][0] +
                mat_A[53][0] * mat_B[162][0] +
                mat_A[53][1] * mat_B[170][0] +
                mat_A[53][2] * mat_B[178][0] +
                mat_A[53][3] * mat_B[186][0] +
                mat_A[54][0] * mat_B[194][0] +
                mat_A[54][1] * mat_B[202][0] +
                mat_A[54][2] * mat_B[210][0] +
                mat_A[54][3] * mat_B[218][0] +
                mat_A[55][0] * mat_B[226][0] +
                mat_A[55][1] * mat_B[234][0] +
                mat_A[55][2] * mat_B[242][0] +
                mat_A[55][3] * mat_B[250][0];
    mat_C[50][1] <=
                mat_A[48][0] * mat_B[2][1] +
                mat_A[48][1] * mat_B[10][1] +
                mat_A[48][2] * mat_B[18][1] +
                mat_A[48][3] * mat_B[26][1] +
                mat_A[49][0] * mat_B[34][1] +
                mat_A[49][1] * mat_B[42][1] +
                mat_A[49][2] * mat_B[50][1] +
                mat_A[49][3] * mat_B[58][1] +
                mat_A[50][0] * mat_B[66][1] +
                mat_A[50][1] * mat_B[74][1] +
                mat_A[50][2] * mat_B[82][1] +
                mat_A[50][3] * mat_B[90][1] +
                mat_A[51][0] * mat_B[98][1] +
                mat_A[51][1] * mat_B[106][1] +
                mat_A[51][2] * mat_B[114][1] +
                mat_A[51][3] * mat_B[122][1] +
                mat_A[52][0] * mat_B[130][1] +
                mat_A[52][1] * mat_B[138][1] +
                mat_A[52][2] * mat_B[146][1] +
                mat_A[52][3] * mat_B[154][1] +
                mat_A[53][0] * mat_B[162][1] +
                mat_A[53][1] * mat_B[170][1] +
                mat_A[53][2] * mat_B[178][1] +
                mat_A[53][3] * mat_B[186][1] +
                mat_A[54][0] * mat_B[194][1] +
                mat_A[54][1] * mat_B[202][1] +
                mat_A[54][2] * mat_B[210][1] +
                mat_A[54][3] * mat_B[218][1] +
                mat_A[55][0] * mat_B[226][1] +
                mat_A[55][1] * mat_B[234][1] +
                mat_A[55][2] * mat_B[242][1] +
                mat_A[55][3] * mat_B[250][1];
    mat_C[50][2] <=
                mat_A[48][0] * mat_B[2][2] +
                mat_A[48][1] * mat_B[10][2] +
                mat_A[48][2] * mat_B[18][2] +
                mat_A[48][3] * mat_B[26][2] +
                mat_A[49][0] * mat_B[34][2] +
                mat_A[49][1] * mat_B[42][2] +
                mat_A[49][2] * mat_B[50][2] +
                mat_A[49][3] * mat_B[58][2] +
                mat_A[50][0] * mat_B[66][2] +
                mat_A[50][1] * mat_B[74][2] +
                mat_A[50][2] * mat_B[82][2] +
                mat_A[50][3] * mat_B[90][2] +
                mat_A[51][0] * mat_B[98][2] +
                mat_A[51][1] * mat_B[106][2] +
                mat_A[51][2] * mat_B[114][2] +
                mat_A[51][3] * mat_B[122][2] +
                mat_A[52][0] * mat_B[130][2] +
                mat_A[52][1] * mat_B[138][2] +
                mat_A[52][2] * mat_B[146][2] +
                mat_A[52][3] * mat_B[154][2] +
                mat_A[53][0] * mat_B[162][2] +
                mat_A[53][1] * mat_B[170][2] +
                mat_A[53][2] * mat_B[178][2] +
                mat_A[53][3] * mat_B[186][2] +
                mat_A[54][0] * mat_B[194][2] +
                mat_A[54][1] * mat_B[202][2] +
                mat_A[54][2] * mat_B[210][2] +
                mat_A[54][3] * mat_B[218][2] +
                mat_A[55][0] * mat_B[226][2] +
                mat_A[55][1] * mat_B[234][2] +
                mat_A[55][2] * mat_B[242][2] +
                mat_A[55][3] * mat_B[250][2];
    mat_C[50][3] <=
                mat_A[48][0] * mat_B[2][3] +
                mat_A[48][1] * mat_B[10][3] +
                mat_A[48][2] * mat_B[18][3] +
                mat_A[48][3] * mat_B[26][3] +
                mat_A[49][0] * mat_B[34][3] +
                mat_A[49][1] * mat_B[42][3] +
                mat_A[49][2] * mat_B[50][3] +
                mat_A[49][3] * mat_B[58][3] +
                mat_A[50][0] * mat_B[66][3] +
                mat_A[50][1] * mat_B[74][3] +
                mat_A[50][2] * mat_B[82][3] +
                mat_A[50][3] * mat_B[90][3] +
                mat_A[51][0] * mat_B[98][3] +
                mat_A[51][1] * mat_B[106][3] +
                mat_A[51][2] * mat_B[114][3] +
                mat_A[51][3] * mat_B[122][3] +
                mat_A[52][0] * mat_B[130][3] +
                mat_A[52][1] * mat_B[138][3] +
                mat_A[52][2] * mat_B[146][3] +
                mat_A[52][3] * mat_B[154][3] +
                mat_A[53][0] * mat_B[162][3] +
                mat_A[53][1] * mat_B[170][3] +
                mat_A[53][2] * mat_B[178][3] +
                mat_A[53][3] * mat_B[186][3] +
                mat_A[54][0] * mat_B[194][3] +
                mat_A[54][1] * mat_B[202][3] +
                mat_A[54][2] * mat_B[210][3] +
                mat_A[54][3] * mat_B[218][3] +
                mat_A[55][0] * mat_B[226][3] +
                mat_A[55][1] * mat_B[234][3] +
                mat_A[55][2] * mat_B[242][3] +
                mat_A[55][3] * mat_B[250][3];
    mat_C[51][0] <=
                mat_A[48][0] * mat_B[3][0] +
                mat_A[48][1] * mat_B[11][0] +
                mat_A[48][2] * mat_B[19][0] +
                mat_A[48][3] * mat_B[27][0] +
                mat_A[49][0] * mat_B[35][0] +
                mat_A[49][1] * mat_B[43][0] +
                mat_A[49][2] * mat_B[51][0] +
                mat_A[49][3] * mat_B[59][0] +
                mat_A[50][0] * mat_B[67][0] +
                mat_A[50][1] * mat_B[75][0] +
                mat_A[50][2] * mat_B[83][0] +
                mat_A[50][3] * mat_B[91][0] +
                mat_A[51][0] * mat_B[99][0] +
                mat_A[51][1] * mat_B[107][0] +
                mat_A[51][2] * mat_B[115][0] +
                mat_A[51][3] * mat_B[123][0] +
                mat_A[52][0] * mat_B[131][0] +
                mat_A[52][1] * mat_B[139][0] +
                mat_A[52][2] * mat_B[147][0] +
                mat_A[52][3] * mat_B[155][0] +
                mat_A[53][0] * mat_B[163][0] +
                mat_A[53][1] * mat_B[171][0] +
                mat_A[53][2] * mat_B[179][0] +
                mat_A[53][3] * mat_B[187][0] +
                mat_A[54][0] * mat_B[195][0] +
                mat_A[54][1] * mat_B[203][0] +
                mat_A[54][2] * mat_B[211][0] +
                mat_A[54][3] * mat_B[219][0] +
                mat_A[55][0] * mat_B[227][0] +
                mat_A[55][1] * mat_B[235][0] +
                mat_A[55][2] * mat_B[243][0] +
                mat_A[55][3] * mat_B[251][0];
    mat_C[51][1] <=
                mat_A[48][0] * mat_B[3][1] +
                mat_A[48][1] * mat_B[11][1] +
                mat_A[48][2] * mat_B[19][1] +
                mat_A[48][3] * mat_B[27][1] +
                mat_A[49][0] * mat_B[35][1] +
                mat_A[49][1] * mat_B[43][1] +
                mat_A[49][2] * mat_B[51][1] +
                mat_A[49][3] * mat_B[59][1] +
                mat_A[50][0] * mat_B[67][1] +
                mat_A[50][1] * mat_B[75][1] +
                mat_A[50][2] * mat_B[83][1] +
                mat_A[50][3] * mat_B[91][1] +
                mat_A[51][0] * mat_B[99][1] +
                mat_A[51][1] * mat_B[107][1] +
                mat_A[51][2] * mat_B[115][1] +
                mat_A[51][3] * mat_B[123][1] +
                mat_A[52][0] * mat_B[131][1] +
                mat_A[52][1] * mat_B[139][1] +
                mat_A[52][2] * mat_B[147][1] +
                mat_A[52][3] * mat_B[155][1] +
                mat_A[53][0] * mat_B[163][1] +
                mat_A[53][1] * mat_B[171][1] +
                mat_A[53][2] * mat_B[179][1] +
                mat_A[53][3] * mat_B[187][1] +
                mat_A[54][0] * mat_B[195][1] +
                mat_A[54][1] * mat_B[203][1] +
                mat_A[54][2] * mat_B[211][1] +
                mat_A[54][3] * mat_B[219][1] +
                mat_A[55][0] * mat_B[227][1] +
                mat_A[55][1] * mat_B[235][1] +
                mat_A[55][2] * mat_B[243][1] +
                mat_A[55][3] * mat_B[251][1];
    mat_C[51][2] <=
                mat_A[48][0] * mat_B[3][2] +
                mat_A[48][1] * mat_B[11][2] +
                mat_A[48][2] * mat_B[19][2] +
                mat_A[48][3] * mat_B[27][2] +
                mat_A[49][0] * mat_B[35][2] +
                mat_A[49][1] * mat_B[43][2] +
                mat_A[49][2] * mat_B[51][2] +
                mat_A[49][3] * mat_B[59][2] +
                mat_A[50][0] * mat_B[67][2] +
                mat_A[50][1] * mat_B[75][2] +
                mat_A[50][2] * mat_B[83][2] +
                mat_A[50][3] * mat_B[91][2] +
                mat_A[51][0] * mat_B[99][2] +
                mat_A[51][1] * mat_B[107][2] +
                mat_A[51][2] * mat_B[115][2] +
                mat_A[51][3] * mat_B[123][2] +
                mat_A[52][0] * mat_B[131][2] +
                mat_A[52][1] * mat_B[139][2] +
                mat_A[52][2] * mat_B[147][2] +
                mat_A[52][3] * mat_B[155][2] +
                mat_A[53][0] * mat_B[163][2] +
                mat_A[53][1] * mat_B[171][2] +
                mat_A[53][2] * mat_B[179][2] +
                mat_A[53][3] * mat_B[187][2] +
                mat_A[54][0] * mat_B[195][2] +
                mat_A[54][1] * mat_B[203][2] +
                mat_A[54][2] * mat_B[211][2] +
                mat_A[54][3] * mat_B[219][2] +
                mat_A[55][0] * mat_B[227][2] +
                mat_A[55][1] * mat_B[235][2] +
                mat_A[55][2] * mat_B[243][2] +
                mat_A[55][3] * mat_B[251][2];
    mat_C[51][3] <=
                mat_A[48][0] * mat_B[3][3] +
                mat_A[48][1] * mat_B[11][3] +
                mat_A[48][2] * mat_B[19][3] +
                mat_A[48][3] * mat_B[27][3] +
                mat_A[49][0] * mat_B[35][3] +
                mat_A[49][1] * mat_B[43][3] +
                mat_A[49][2] * mat_B[51][3] +
                mat_A[49][3] * mat_B[59][3] +
                mat_A[50][0] * mat_B[67][3] +
                mat_A[50][1] * mat_B[75][3] +
                mat_A[50][2] * mat_B[83][3] +
                mat_A[50][3] * mat_B[91][3] +
                mat_A[51][0] * mat_B[99][3] +
                mat_A[51][1] * mat_B[107][3] +
                mat_A[51][2] * mat_B[115][3] +
                mat_A[51][3] * mat_B[123][3] +
                mat_A[52][0] * mat_B[131][3] +
                mat_A[52][1] * mat_B[139][3] +
                mat_A[52][2] * mat_B[147][3] +
                mat_A[52][3] * mat_B[155][3] +
                mat_A[53][0] * mat_B[163][3] +
                mat_A[53][1] * mat_B[171][3] +
                mat_A[53][2] * mat_B[179][3] +
                mat_A[53][3] * mat_B[187][3] +
                mat_A[54][0] * mat_B[195][3] +
                mat_A[54][1] * mat_B[203][3] +
                mat_A[54][2] * mat_B[211][3] +
                mat_A[54][3] * mat_B[219][3] +
                mat_A[55][0] * mat_B[227][3] +
                mat_A[55][1] * mat_B[235][3] +
                mat_A[55][2] * mat_B[243][3] +
                mat_A[55][3] * mat_B[251][3];
    mat_C[52][0] <=
                mat_A[48][0] * mat_B[4][0] +
                mat_A[48][1] * mat_B[12][0] +
                mat_A[48][2] * mat_B[20][0] +
                mat_A[48][3] * mat_B[28][0] +
                mat_A[49][0] * mat_B[36][0] +
                mat_A[49][1] * mat_B[44][0] +
                mat_A[49][2] * mat_B[52][0] +
                mat_A[49][3] * mat_B[60][0] +
                mat_A[50][0] * mat_B[68][0] +
                mat_A[50][1] * mat_B[76][0] +
                mat_A[50][2] * mat_B[84][0] +
                mat_A[50][3] * mat_B[92][0] +
                mat_A[51][0] * mat_B[100][0] +
                mat_A[51][1] * mat_B[108][0] +
                mat_A[51][2] * mat_B[116][0] +
                mat_A[51][3] * mat_B[124][0] +
                mat_A[52][0] * mat_B[132][0] +
                mat_A[52][1] * mat_B[140][0] +
                mat_A[52][2] * mat_B[148][0] +
                mat_A[52][3] * mat_B[156][0] +
                mat_A[53][0] * mat_B[164][0] +
                mat_A[53][1] * mat_B[172][0] +
                mat_A[53][2] * mat_B[180][0] +
                mat_A[53][3] * mat_B[188][0] +
                mat_A[54][0] * mat_B[196][0] +
                mat_A[54][1] * mat_B[204][0] +
                mat_A[54][2] * mat_B[212][0] +
                mat_A[54][3] * mat_B[220][0] +
                mat_A[55][0] * mat_B[228][0] +
                mat_A[55][1] * mat_B[236][0] +
                mat_A[55][2] * mat_B[244][0] +
                mat_A[55][3] * mat_B[252][0];
    mat_C[52][1] <=
                mat_A[48][0] * mat_B[4][1] +
                mat_A[48][1] * mat_B[12][1] +
                mat_A[48][2] * mat_B[20][1] +
                mat_A[48][3] * mat_B[28][1] +
                mat_A[49][0] * mat_B[36][1] +
                mat_A[49][1] * mat_B[44][1] +
                mat_A[49][2] * mat_B[52][1] +
                mat_A[49][3] * mat_B[60][1] +
                mat_A[50][0] * mat_B[68][1] +
                mat_A[50][1] * mat_B[76][1] +
                mat_A[50][2] * mat_B[84][1] +
                mat_A[50][3] * mat_B[92][1] +
                mat_A[51][0] * mat_B[100][1] +
                mat_A[51][1] * mat_B[108][1] +
                mat_A[51][2] * mat_B[116][1] +
                mat_A[51][3] * mat_B[124][1] +
                mat_A[52][0] * mat_B[132][1] +
                mat_A[52][1] * mat_B[140][1] +
                mat_A[52][2] * mat_B[148][1] +
                mat_A[52][3] * mat_B[156][1] +
                mat_A[53][0] * mat_B[164][1] +
                mat_A[53][1] * mat_B[172][1] +
                mat_A[53][2] * mat_B[180][1] +
                mat_A[53][3] * mat_B[188][1] +
                mat_A[54][0] * mat_B[196][1] +
                mat_A[54][1] * mat_B[204][1] +
                mat_A[54][2] * mat_B[212][1] +
                mat_A[54][3] * mat_B[220][1] +
                mat_A[55][0] * mat_B[228][1] +
                mat_A[55][1] * mat_B[236][1] +
                mat_A[55][2] * mat_B[244][1] +
                mat_A[55][3] * mat_B[252][1];
    mat_C[52][2] <=
                mat_A[48][0] * mat_B[4][2] +
                mat_A[48][1] * mat_B[12][2] +
                mat_A[48][2] * mat_B[20][2] +
                mat_A[48][3] * mat_B[28][2] +
                mat_A[49][0] * mat_B[36][2] +
                mat_A[49][1] * mat_B[44][2] +
                mat_A[49][2] * mat_B[52][2] +
                mat_A[49][3] * mat_B[60][2] +
                mat_A[50][0] * mat_B[68][2] +
                mat_A[50][1] * mat_B[76][2] +
                mat_A[50][2] * mat_B[84][2] +
                mat_A[50][3] * mat_B[92][2] +
                mat_A[51][0] * mat_B[100][2] +
                mat_A[51][1] * mat_B[108][2] +
                mat_A[51][2] * mat_B[116][2] +
                mat_A[51][3] * mat_B[124][2] +
                mat_A[52][0] * mat_B[132][2] +
                mat_A[52][1] * mat_B[140][2] +
                mat_A[52][2] * mat_B[148][2] +
                mat_A[52][3] * mat_B[156][2] +
                mat_A[53][0] * mat_B[164][2] +
                mat_A[53][1] * mat_B[172][2] +
                mat_A[53][2] * mat_B[180][2] +
                mat_A[53][3] * mat_B[188][2] +
                mat_A[54][0] * mat_B[196][2] +
                mat_A[54][1] * mat_B[204][2] +
                mat_A[54][2] * mat_B[212][2] +
                mat_A[54][3] * mat_B[220][2] +
                mat_A[55][0] * mat_B[228][2] +
                mat_A[55][1] * mat_B[236][2] +
                mat_A[55][2] * mat_B[244][2] +
                mat_A[55][3] * mat_B[252][2];
    mat_C[52][3] <=
                mat_A[48][0] * mat_B[4][3] +
                mat_A[48][1] * mat_B[12][3] +
                mat_A[48][2] * mat_B[20][3] +
                mat_A[48][3] * mat_B[28][3] +
                mat_A[49][0] * mat_B[36][3] +
                mat_A[49][1] * mat_B[44][3] +
                mat_A[49][2] * mat_B[52][3] +
                mat_A[49][3] * mat_B[60][3] +
                mat_A[50][0] * mat_B[68][3] +
                mat_A[50][1] * mat_B[76][3] +
                mat_A[50][2] * mat_B[84][3] +
                mat_A[50][3] * mat_B[92][3] +
                mat_A[51][0] * mat_B[100][3] +
                mat_A[51][1] * mat_B[108][3] +
                mat_A[51][2] * mat_B[116][3] +
                mat_A[51][3] * mat_B[124][3] +
                mat_A[52][0] * mat_B[132][3] +
                mat_A[52][1] * mat_B[140][3] +
                mat_A[52][2] * mat_B[148][3] +
                mat_A[52][3] * mat_B[156][3] +
                mat_A[53][0] * mat_B[164][3] +
                mat_A[53][1] * mat_B[172][3] +
                mat_A[53][2] * mat_B[180][3] +
                mat_A[53][3] * mat_B[188][3] +
                mat_A[54][0] * mat_B[196][3] +
                mat_A[54][1] * mat_B[204][3] +
                mat_A[54][2] * mat_B[212][3] +
                mat_A[54][3] * mat_B[220][3] +
                mat_A[55][0] * mat_B[228][3] +
                mat_A[55][1] * mat_B[236][3] +
                mat_A[55][2] * mat_B[244][3] +
                mat_A[55][3] * mat_B[252][3];
    mat_C[53][0] <=
                mat_A[48][0] * mat_B[5][0] +
                mat_A[48][1] * mat_B[13][0] +
                mat_A[48][2] * mat_B[21][0] +
                mat_A[48][3] * mat_B[29][0] +
                mat_A[49][0] * mat_B[37][0] +
                mat_A[49][1] * mat_B[45][0] +
                mat_A[49][2] * mat_B[53][0] +
                mat_A[49][3] * mat_B[61][0] +
                mat_A[50][0] * mat_B[69][0] +
                mat_A[50][1] * mat_B[77][0] +
                mat_A[50][2] * mat_B[85][0] +
                mat_A[50][3] * mat_B[93][0] +
                mat_A[51][0] * mat_B[101][0] +
                mat_A[51][1] * mat_B[109][0] +
                mat_A[51][2] * mat_B[117][0] +
                mat_A[51][3] * mat_B[125][0] +
                mat_A[52][0] * mat_B[133][0] +
                mat_A[52][1] * mat_B[141][0] +
                mat_A[52][2] * mat_B[149][0] +
                mat_A[52][3] * mat_B[157][0] +
                mat_A[53][0] * mat_B[165][0] +
                mat_A[53][1] * mat_B[173][0] +
                mat_A[53][2] * mat_B[181][0] +
                mat_A[53][3] * mat_B[189][0] +
                mat_A[54][0] * mat_B[197][0] +
                mat_A[54][1] * mat_B[205][0] +
                mat_A[54][2] * mat_B[213][0] +
                mat_A[54][3] * mat_B[221][0] +
                mat_A[55][0] * mat_B[229][0] +
                mat_A[55][1] * mat_B[237][0] +
                mat_A[55][2] * mat_B[245][0] +
                mat_A[55][3] * mat_B[253][0];
    mat_C[53][1] <=
                mat_A[48][0] * mat_B[5][1] +
                mat_A[48][1] * mat_B[13][1] +
                mat_A[48][2] * mat_B[21][1] +
                mat_A[48][3] * mat_B[29][1] +
                mat_A[49][0] * mat_B[37][1] +
                mat_A[49][1] * mat_B[45][1] +
                mat_A[49][2] * mat_B[53][1] +
                mat_A[49][3] * mat_B[61][1] +
                mat_A[50][0] * mat_B[69][1] +
                mat_A[50][1] * mat_B[77][1] +
                mat_A[50][2] * mat_B[85][1] +
                mat_A[50][3] * mat_B[93][1] +
                mat_A[51][0] * mat_B[101][1] +
                mat_A[51][1] * mat_B[109][1] +
                mat_A[51][2] * mat_B[117][1] +
                mat_A[51][3] * mat_B[125][1] +
                mat_A[52][0] * mat_B[133][1] +
                mat_A[52][1] * mat_B[141][1] +
                mat_A[52][2] * mat_B[149][1] +
                mat_A[52][3] * mat_B[157][1] +
                mat_A[53][0] * mat_B[165][1] +
                mat_A[53][1] * mat_B[173][1] +
                mat_A[53][2] * mat_B[181][1] +
                mat_A[53][3] * mat_B[189][1] +
                mat_A[54][0] * mat_B[197][1] +
                mat_A[54][1] * mat_B[205][1] +
                mat_A[54][2] * mat_B[213][1] +
                mat_A[54][3] * mat_B[221][1] +
                mat_A[55][0] * mat_B[229][1] +
                mat_A[55][1] * mat_B[237][1] +
                mat_A[55][2] * mat_B[245][1] +
                mat_A[55][3] * mat_B[253][1];
    mat_C[53][2] <=
                mat_A[48][0] * mat_B[5][2] +
                mat_A[48][1] * mat_B[13][2] +
                mat_A[48][2] * mat_B[21][2] +
                mat_A[48][3] * mat_B[29][2] +
                mat_A[49][0] * mat_B[37][2] +
                mat_A[49][1] * mat_B[45][2] +
                mat_A[49][2] * mat_B[53][2] +
                mat_A[49][3] * mat_B[61][2] +
                mat_A[50][0] * mat_B[69][2] +
                mat_A[50][1] * mat_B[77][2] +
                mat_A[50][2] * mat_B[85][2] +
                mat_A[50][3] * mat_B[93][2] +
                mat_A[51][0] * mat_B[101][2] +
                mat_A[51][1] * mat_B[109][2] +
                mat_A[51][2] * mat_B[117][2] +
                mat_A[51][3] * mat_B[125][2] +
                mat_A[52][0] * mat_B[133][2] +
                mat_A[52][1] * mat_B[141][2] +
                mat_A[52][2] * mat_B[149][2] +
                mat_A[52][3] * mat_B[157][2] +
                mat_A[53][0] * mat_B[165][2] +
                mat_A[53][1] * mat_B[173][2] +
                mat_A[53][2] * mat_B[181][2] +
                mat_A[53][3] * mat_B[189][2] +
                mat_A[54][0] * mat_B[197][2] +
                mat_A[54][1] * mat_B[205][2] +
                mat_A[54][2] * mat_B[213][2] +
                mat_A[54][3] * mat_B[221][2] +
                mat_A[55][0] * mat_B[229][2] +
                mat_A[55][1] * mat_B[237][2] +
                mat_A[55][2] * mat_B[245][2] +
                mat_A[55][3] * mat_B[253][2];
    mat_C[53][3] <=
                mat_A[48][0] * mat_B[5][3] +
                mat_A[48][1] * mat_B[13][3] +
                mat_A[48][2] * mat_B[21][3] +
                mat_A[48][3] * mat_B[29][3] +
                mat_A[49][0] * mat_B[37][3] +
                mat_A[49][1] * mat_B[45][3] +
                mat_A[49][2] * mat_B[53][3] +
                mat_A[49][3] * mat_B[61][3] +
                mat_A[50][0] * mat_B[69][3] +
                mat_A[50][1] * mat_B[77][3] +
                mat_A[50][2] * mat_B[85][3] +
                mat_A[50][3] * mat_B[93][3] +
                mat_A[51][0] * mat_B[101][3] +
                mat_A[51][1] * mat_B[109][3] +
                mat_A[51][2] * mat_B[117][3] +
                mat_A[51][3] * mat_B[125][3] +
                mat_A[52][0] * mat_B[133][3] +
                mat_A[52][1] * mat_B[141][3] +
                mat_A[52][2] * mat_B[149][3] +
                mat_A[52][3] * mat_B[157][3] +
                mat_A[53][0] * mat_B[165][3] +
                mat_A[53][1] * mat_B[173][3] +
                mat_A[53][2] * mat_B[181][3] +
                mat_A[53][3] * mat_B[189][3] +
                mat_A[54][0] * mat_B[197][3] +
                mat_A[54][1] * mat_B[205][3] +
                mat_A[54][2] * mat_B[213][3] +
                mat_A[54][3] * mat_B[221][3] +
                mat_A[55][0] * mat_B[229][3] +
                mat_A[55][1] * mat_B[237][3] +
                mat_A[55][2] * mat_B[245][3] +
                mat_A[55][3] * mat_B[253][3];
    mat_C[54][0] <=
                mat_A[48][0] * mat_B[6][0] +
                mat_A[48][1] * mat_B[14][0] +
                mat_A[48][2] * mat_B[22][0] +
                mat_A[48][3] * mat_B[30][0] +
                mat_A[49][0] * mat_B[38][0] +
                mat_A[49][1] * mat_B[46][0] +
                mat_A[49][2] * mat_B[54][0] +
                mat_A[49][3] * mat_B[62][0] +
                mat_A[50][0] * mat_B[70][0] +
                mat_A[50][1] * mat_B[78][0] +
                mat_A[50][2] * mat_B[86][0] +
                mat_A[50][3] * mat_B[94][0] +
                mat_A[51][0] * mat_B[102][0] +
                mat_A[51][1] * mat_B[110][0] +
                mat_A[51][2] * mat_B[118][0] +
                mat_A[51][3] * mat_B[126][0] +
                mat_A[52][0] * mat_B[134][0] +
                mat_A[52][1] * mat_B[142][0] +
                mat_A[52][2] * mat_B[150][0] +
                mat_A[52][3] * mat_B[158][0] +
                mat_A[53][0] * mat_B[166][0] +
                mat_A[53][1] * mat_B[174][0] +
                mat_A[53][2] * mat_B[182][0] +
                mat_A[53][3] * mat_B[190][0] +
                mat_A[54][0] * mat_B[198][0] +
                mat_A[54][1] * mat_B[206][0] +
                mat_A[54][2] * mat_B[214][0] +
                mat_A[54][3] * mat_B[222][0] +
                mat_A[55][0] * mat_B[230][0] +
                mat_A[55][1] * mat_B[238][0] +
                mat_A[55][2] * mat_B[246][0] +
                mat_A[55][3] * mat_B[254][0];
    mat_C[54][1] <=
                mat_A[48][0] * mat_B[6][1] +
                mat_A[48][1] * mat_B[14][1] +
                mat_A[48][2] * mat_B[22][1] +
                mat_A[48][3] * mat_B[30][1] +
                mat_A[49][0] * mat_B[38][1] +
                mat_A[49][1] * mat_B[46][1] +
                mat_A[49][2] * mat_B[54][1] +
                mat_A[49][3] * mat_B[62][1] +
                mat_A[50][0] * mat_B[70][1] +
                mat_A[50][1] * mat_B[78][1] +
                mat_A[50][2] * mat_B[86][1] +
                mat_A[50][3] * mat_B[94][1] +
                mat_A[51][0] * mat_B[102][1] +
                mat_A[51][1] * mat_B[110][1] +
                mat_A[51][2] * mat_B[118][1] +
                mat_A[51][3] * mat_B[126][1] +
                mat_A[52][0] * mat_B[134][1] +
                mat_A[52][1] * mat_B[142][1] +
                mat_A[52][2] * mat_B[150][1] +
                mat_A[52][3] * mat_B[158][1] +
                mat_A[53][0] * mat_B[166][1] +
                mat_A[53][1] * mat_B[174][1] +
                mat_A[53][2] * mat_B[182][1] +
                mat_A[53][3] * mat_B[190][1] +
                mat_A[54][0] * mat_B[198][1] +
                mat_A[54][1] * mat_B[206][1] +
                mat_A[54][2] * mat_B[214][1] +
                mat_A[54][3] * mat_B[222][1] +
                mat_A[55][0] * mat_B[230][1] +
                mat_A[55][1] * mat_B[238][1] +
                mat_A[55][2] * mat_B[246][1] +
                mat_A[55][3] * mat_B[254][1];
    mat_C[54][2] <=
                mat_A[48][0] * mat_B[6][2] +
                mat_A[48][1] * mat_B[14][2] +
                mat_A[48][2] * mat_B[22][2] +
                mat_A[48][3] * mat_B[30][2] +
                mat_A[49][0] * mat_B[38][2] +
                mat_A[49][1] * mat_B[46][2] +
                mat_A[49][2] * mat_B[54][2] +
                mat_A[49][3] * mat_B[62][2] +
                mat_A[50][0] * mat_B[70][2] +
                mat_A[50][1] * mat_B[78][2] +
                mat_A[50][2] * mat_B[86][2] +
                mat_A[50][3] * mat_B[94][2] +
                mat_A[51][0] * mat_B[102][2] +
                mat_A[51][1] * mat_B[110][2] +
                mat_A[51][2] * mat_B[118][2] +
                mat_A[51][3] * mat_B[126][2] +
                mat_A[52][0] * mat_B[134][2] +
                mat_A[52][1] * mat_B[142][2] +
                mat_A[52][2] * mat_B[150][2] +
                mat_A[52][3] * mat_B[158][2] +
                mat_A[53][0] * mat_B[166][2] +
                mat_A[53][1] * mat_B[174][2] +
                mat_A[53][2] * mat_B[182][2] +
                mat_A[53][3] * mat_B[190][2] +
                mat_A[54][0] * mat_B[198][2] +
                mat_A[54][1] * mat_B[206][2] +
                mat_A[54][2] * mat_B[214][2] +
                mat_A[54][3] * mat_B[222][2] +
                mat_A[55][0] * mat_B[230][2] +
                mat_A[55][1] * mat_B[238][2] +
                mat_A[55][2] * mat_B[246][2] +
                mat_A[55][3] * mat_B[254][2];
    mat_C[54][3] <=
                mat_A[48][0] * mat_B[6][3] +
                mat_A[48][1] * mat_B[14][3] +
                mat_A[48][2] * mat_B[22][3] +
                mat_A[48][3] * mat_B[30][3] +
                mat_A[49][0] * mat_B[38][3] +
                mat_A[49][1] * mat_B[46][3] +
                mat_A[49][2] * mat_B[54][3] +
                mat_A[49][3] * mat_B[62][3] +
                mat_A[50][0] * mat_B[70][3] +
                mat_A[50][1] * mat_B[78][3] +
                mat_A[50][2] * mat_B[86][3] +
                mat_A[50][3] * mat_B[94][3] +
                mat_A[51][0] * mat_B[102][3] +
                mat_A[51][1] * mat_B[110][3] +
                mat_A[51][2] * mat_B[118][3] +
                mat_A[51][3] * mat_B[126][3] +
                mat_A[52][0] * mat_B[134][3] +
                mat_A[52][1] * mat_B[142][3] +
                mat_A[52][2] * mat_B[150][3] +
                mat_A[52][3] * mat_B[158][3] +
                mat_A[53][0] * mat_B[166][3] +
                mat_A[53][1] * mat_B[174][3] +
                mat_A[53][2] * mat_B[182][3] +
                mat_A[53][3] * mat_B[190][3] +
                mat_A[54][0] * mat_B[198][3] +
                mat_A[54][1] * mat_B[206][3] +
                mat_A[54][2] * mat_B[214][3] +
                mat_A[54][3] * mat_B[222][3] +
                mat_A[55][0] * mat_B[230][3] +
                mat_A[55][1] * mat_B[238][3] +
                mat_A[55][2] * mat_B[246][3] +
                mat_A[55][3] * mat_B[254][3];
    mat_C[55][0] <=
                mat_A[48][0] * mat_B[7][0] +
                mat_A[48][1] * mat_B[15][0] +
                mat_A[48][2] * mat_B[23][0] +
                mat_A[48][3] * mat_B[31][0] +
                mat_A[49][0] * mat_B[39][0] +
                mat_A[49][1] * mat_B[47][0] +
                mat_A[49][2] * mat_B[55][0] +
                mat_A[49][3] * mat_B[63][0] +
                mat_A[50][0] * mat_B[71][0] +
                mat_A[50][1] * mat_B[79][0] +
                mat_A[50][2] * mat_B[87][0] +
                mat_A[50][3] * mat_B[95][0] +
                mat_A[51][0] * mat_B[103][0] +
                mat_A[51][1] * mat_B[111][0] +
                mat_A[51][2] * mat_B[119][0] +
                mat_A[51][3] * mat_B[127][0] +
                mat_A[52][0] * mat_B[135][0] +
                mat_A[52][1] * mat_B[143][0] +
                mat_A[52][2] * mat_B[151][0] +
                mat_A[52][3] * mat_B[159][0] +
                mat_A[53][0] * mat_B[167][0] +
                mat_A[53][1] * mat_B[175][0] +
                mat_A[53][2] * mat_B[183][0] +
                mat_A[53][3] * mat_B[191][0] +
                mat_A[54][0] * mat_B[199][0] +
                mat_A[54][1] * mat_B[207][0] +
                mat_A[54][2] * mat_B[215][0] +
                mat_A[54][3] * mat_B[223][0] +
                mat_A[55][0] * mat_B[231][0] +
                mat_A[55][1] * mat_B[239][0] +
                mat_A[55][2] * mat_B[247][0] +
                mat_A[55][3] * mat_B[255][0];
    mat_C[55][1] <=
                mat_A[48][0] * mat_B[7][1] +
                mat_A[48][1] * mat_B[15][1] +
                mat_A[48][2] * mat_B[23][1] +
                mat_A[48][3] * mat_B[31][1] +
                mat_A[49][0] * mat_B[39][1] +
                mat_A[49][1] * mat_B[47][1] +
                mat_A[49][2] * mat_B[55][1] +
                mat_A[49][3] * mat_B[63][1] +
                mat_A[50][0] * mat_B[71][1] +
                mat_A[50][1] * mat_B[79][1] +
                mat_A[50][2] * mat_B[87][1] +
                mat_A[50][3] * mat_B[95][1] +
                mat_A[51][0] * mat_B[103][1] +
                mat_A[51][1] * mat_B[111][1] +
                mat_A[51][2] * mat_B[119][1] +
                mat_A[51][3] * mat_B[127][1] +
                mat_A[52][0] * mat_B[135][1] +
                mat_A[52][1] * mat_B[143][1] +
                mat_A[52][2] * mat_B[151][1] +
                mat_A[52][3] * mat_B[159][1] +
                mat_A[53][0] * mat_B[167][1] +
                mat_A[53][1] * mat_B[175][1] +
                mat_A[53][2] * mat_B[183][1] +
                mat_A[53][3] * mat_B[191][1] +
                mat_A[54][0] * mat_B[199][1] +
                mat_A[54][1] * mat_B[207][1] +
                mat_A[54][2] * mat_B[215][1] +
                mat_A[54][3] * mat_B[223][1] +
                mat_A[55][0] * mat_B[231][1] +
                mat_A[55][1] * mat_B[239][1] +
                mat_A[55][2] * mat_B[247][1] +
                mat_A[55][3] * mat_B[255][1];
    mat_C[55][2] <=
                mat_A[48][0] * mat_B[7][2] +
                mat_A[48][1] * mat_B[15][2] +
                mat_A[48][2] * mat_B[23][2] +
                mat_A[48][3] * mat_B[31][2] +
                mat_A[49][0] * mat_B[39][2] +
                mat_A[49][1] * mat_B[47][2] +
                mat_A[49][2] * mat_B[55][2] +
                mat_A[49][3] * mat_B[63][2] +
                mat_A[50][0] * mat_B[71][2] +
                mat_A[50][1] * mat_B[79][2] +
                mat_A[50][2] * mat_B[87][2] +
                mat_A[50][3] * mat_B[95][2] +
                mat_A[51][0] * mat_B[103][2] +
                mat_A[51][1] * mat_B[111][2] +
                mat_A[51][2] * mat_B[119][2] +
                mat_A[51][3] * mat_B[127][2] +
                mat_A[52][0] * mat_B[135][2] +
                mat_A[52][1] * mat_B[143][2] +
                mat_A[52][2] * mat_B[151][2] +
                mat_A[52][3] * mat_B[159][2] +
                mat_A[53][0] * mat_B[167][2] +
                mat_A[53][1] * mat_B[175][2] +
                mat_A[53][2] * mat_B[183][2] +
                mat_A[53][3] * mat_B[191][2] +
                mat_A[54][0] * mat_B[199][2] +
                mat_A[54][1] * mat_B[207][2] +
                mat_A[54][2] * mat_B[215][2] +
                mat_A[54][3] * mat_B[223][2] +
                mat_A[55][0] * mat_B[231][2] +
                mat_A[55][1] * mat_B[239][2] +
                mat_A[55][2] * mat_B[247][2] +
                mat_A[55][3] * mat_B[255][2];
    mat_C[55][3] <=
                mat_A[48][0] * mat_B[7][3] +
                mat_A[48][1] * mat_B[15][3] +
                mat_A[48][2] * mat_B[23][3] +
                mat_A[48][3] * mat_B[31][3] +
                mat_A[49][0] * mat_B[39][3] +
                mat_A[49][1] * mat_B[47][3] +
                mat_A[49][2] * mat_B[55][3] +
                mat_A[49][3] * mat_B[63][3] +
                mat_A[50][0] * mat_B[71][3] +
                mat_A[50][1] * mat_B[79][3] +
                mat_A[50][2] * mat_B[87][3] +
                mat_A[50][3] * mat_B[95][3] +
                mat_A[51][0] * mat_B[103][3] +
                mat_A[51][1] * mat_B[111][3] +
                mat_A[51][2] * mat_B[119][3] +
                mat_A[51][3] * mat_B[127][3] +
                mat_A[52][0] * mat_B[135][3] +
                mat_A[52][1] * mat_B[143][3] +
                mat_A[52][2] * mat_B[151][3] +
                mat_A[52][3] * mat_B[159][3] +
                mat_A[53][0] * mat_B[167][3] +
                mat_A[53][1] * mat_B[175][3] +
                mat_A[53][2] * mat_B[183][3] +
                mat_A[53][3] * mat_B[191][3] +
                mat_A[54][0] * mat_B[199][3] +
                mat_A[54][1] * mat_B[207][3] +
                mat_A[54][2] * mat_B[215][3] +
                mat_A[54][3] * mat_B[223][3] +
                mat_A[55][0] * mat_B[231][3] +
                mat_A[55][1] * mat_B[239][3] +
                mat_A[55][2] * mat_B[247][3] +
                mat_A[55][3] * mat_B[255][3];
    mat_C[56][0] <=
                mat_A[56][0] * mat_B[0][0] +
                mat_A[56][1] * mat_B[8][0] +
                mat_A[56][2] * mat_B[16][0] +
                mat_A[56][3] * mat_B[24][0] +
                mat_A[57][0] * mat_B[32][0] +
                mat_A[57][1] * mat_B[40][0] +
                mat_A[57][2] * mat_B[48][0] +
                mat_A[57][3] * mat_B[56][0] +
                mat_A[58][0] * mat_B[64][0] +
                mat_A[58][1] * mat_B[72][0] +
                mat_A[58][2] * mat_B[80][0] +
                mat_A[58][3] * mat_B[88][0] +
                mat_A[59][0] * mat_B[96][0] +
                mat_A[59][1] * mat_B[104][0] +
                mat_A[59][2] * mat_B[112][0] +
                mat_A[59][3] * mat_B[120][0] +
                mat_A[60][0] * mat_B[128][0] +
                mat_A[60][1] * mat_B[136][0] +
                mat_A[60][2] * mat_B[144][0] +
                mat_A[60][3] * mat_B[152][0] +
                mat_A[61][0] * mat_B[160][0] +
                mat_A[61][1] * mat_B[168][0] +
                mat_A[61][2] * mat_B[176][0] +
                mat_A[61][3] * mat_B[184][0] +
                mat_A[62][0] * mat_B[192][0] +
                mat_A[62][1] * mat_B[200][0] +
                mat_A[62][2] * mat_B[208][0] +
                mat_A[62][3] * mat_B[216][0] +
                mat_A[63][0] * mat_B[224][0] +
                mat_A[63][1] * mat_B[232][0] +
                mat_A[63][2] * mat_B[240][0] +
                mat_A[63][3] * mat_B[248][0];
    mat_C[56][1] <=
                mat_A[56][0] * mat_B[0][1] +
                mat_A[56][1] * mat_B[8][1] +
                mat_A[56][2] * mat_B[16][1] +
                mat_A[56][3] * mat_B[24][1] +
                mat_A[57][0] * mat_B[32][1] +
                mat_A[57][1] * mat_B[40][1] +
                mat_A[57][2] * mat_B[48][1] +
                mat_A[57][3] * mat_B[56][1] +
                mat_A[58][0] * mat_B[64][1] +
                mat_A[58][1] * mat_B[72][1] +
                mat_A[58][2] * mat_B[80][1] +
                mat_A[58][3] * mat_B[88][1] +
                mat_A[59][0] * mat_B[96][1] +
                mat_A[59][1] * mat_B[104][1] +
                mat_A[59][2] * mat_B[112][1] +
                mat_A[59][3] * mat_B[120][1] +
                mat_A[60][0] * mat_B[128][1] +
                mat_A[60][1] * mat_B[136][1] +
                mat_A[60][2] * mat_B[144][1] +
                mat_A[60][3] * mat_B[152][1] +
                mat_A[61][0] * mat_B[160][1] +
                mat_A[61][1] * mat_B[168][1] +
                mat_A[61][2] * mat_B[176][1] +
                mat_A[61][3] * mat_B[184][1] +
                mat_A[62][0] * mat_B[192][1] +
                mat_A[62][1] * mat_B[200][1] +
                mat_A[62][2] * mat_B[208][1] +
                mat_A[62][3] * mat_B[216][1] +
                mat_A[63][0] * mat_B[224][1] +
                mat_A[63][1] * mat_B[232][1] +
                mat_A[63][2] * mat_B[240][1] +
                mat_A[63][3] * mat_B[248][1];
    mat_C[56][2] <=
                mat_A[56][0] * mat_B[0][2] +
                mat_A[56][1] * mat_B[8][2] +
                mat_A[56][2] * mat_B[16][2] +
                mat_A[56][3] * mat_B[24][2] +
                mat_A[57][0] * mat_B[32][2] +
                mat_A[57][1] * mat_B[40][2] +
                mat_A[57][2] * mat_B[48][2] +
                mat_A[57][3] * mat_B[56][2] +
                mat_A[58][0] * mat_B[64][2] +
                mat_A[58][1] * mat_B[72][2] +
                mat_A[58][2] * mat_B[80][2] +
                mat_A[58][3] * mat_B[88][2] +
                mat_A[59][0] * mat_B[96][2] +
                mat_A[59][1] * mat_B[104][2] +
                mat_A[59][2] * mat_B[112][2] +
                mat_A[59][3] * mat_B[120][2] +
                mat_A[60][0] * mat_B[128][2] +
                mat_A[60][1] * mat_B[136][2] +
                mat_A[60][2] * mat_B[144][2] +
                mat_A[60][3] * mat_B[152][2] +
                mat_A[61][0] * mat_B[160][2] +
                mat_A[61][1] * mat_B[168][2] +
                mat_A[61][2] * mat_B[176][2] +
                mat_A[61][3] * mat_B[184][2] +
                mat_A[62][0] * mat_B[192][2] +
                mat_A[62][1] * mat_B[200][2] +
                mat_A[62][2] * mat_B[208][2] +
                mat_A[62][3] * mat_B[216][2] +
                mat_A[63][0] * mat_B[224][2] +
                mat_A[63][1] * mat_B[232][2] +
                mat_A[63][2] * mat_B[240][2] +
                mat_A[63][3] * mat_B[248][2];
    mat_C[56][3] <=
                mat_A[56][0] * mat_B[0][3] +
                mat_A[56][1] * mat_B[8][3] +
                mat_A[56][2] * mat_B[16][3] +
                mat_A[56][3] * mat_B[24][3] +
                mat_A[57][0] * mat_B[32][3] +
                mat_A[57][1] * mat_B[40][3] +
                mat_A[57][2] * mat_B[48][3] +
                mat_A[57][3] * mat_B[56][3] +
                mat_A[58][0] * mat_B[64][3] +
                mat_A[58][1] * mat_B[72][3] +
                mat_A[58][2] * mat_B[80][3] +
                mat_A[58][3] * mat_B[88][3] +
                mat_A[59][0] * mat_B[96][3] +
                mat_A[59][1] * mat_B[104][3] +
                mat_A[59][2] * mat_B[112][3] +
                mat_A[59][3] * mat_B[120][3] +
                mat_A[60][0] * mat_B[128][3] +
                mat_A[60][1] * mat_B[136][3] +
                mat_A[60][2] * mat_B[144][3] +
                mat_A[60][3] * mat_B[152][3] +
                mat_A[61][0] * mat_B[160][3] +
                mat_A[61][1] * mat_B[168][3] +
                mat_A[61][2] * mat_B[176][3] +
                mat_A[61][3] * mat_B[184][3] +
                mat_A[62][0] * mat_B[192][3] +
                mat_A[62][1] * mat_B[200][3] +
                mat_A[62][2] * mat_B[208][3] +
                mat_A[62][3] * mat_B[216][3] +
                mat_A[63][0] * mat_B[224][3] +
                mat_A[63][1] * mat_B[232][3] +
                mat_A[63][2] * mat_B[240][3] +
                mat_A[63][3] * mat_B[248][3];
    mat_C[57][0] <=
                mat_A[56][0] * mat_B[1][0] +
                mat_A[56][1] * mat_B[9][0] +
                mat_A[56][2] * mat_B[17][0] +
                mat_A[56][3] * mat_B[25][0] +
                mat_A[57][0] * mat_B[33][0] +
                mat_A[57][1] * mat_B[41][0] +
                mat_A[57][2] * mat_B[49][0] +
                mat_A[57][3] * mat_B[57][0] +
                mat_A[58][0] * mat_B[65][0] +
                mat_A[58][1] * mat_B[73][0] +
                mat_A[58][2] * mat_B[81][0] +
                mat_A[58][3] * mat_B[89][0] +
                mat_A[59][0] * mat_B[97][0] +
                mat_A[59][1] * mat_B[105][0] +
                mat_A[59][2] * mat_B[113][0] +
                mat_A[59][3] * mat_B[121][0] +
                mat_A[60][0] * mat_B[129][0] +
                mat_A[60][1] * mat_B[137][0] +
                mat_A[60][2] * mat_B[145][0] +
                mat_A[60][3] * mat_B[153][0] +
                mat_A[61][0] * mat_B[161][0] +
                mat_A[61][1] * mat_B[169][0] +
                mat_A[61][2] * mat_B[177][0] +
                mat_A[61][3] * mat_B[185][0] +
                mat_A[62][0] * mat_B[193][0] +
                mat_A[62][1] * mat_B[201][0] +
                mat_A[62][2] * mat_B[209][0] +
                mat_A[62][3] * mat_B[217][0] +
                mat_A[63][0] * mat_B[225][0] +
                mat_A[63][1] * mat_B[233][0] +
                mat_A[63][2] * mat_B[241][0] +
                mat_A[63][3] * mat_B[249][0];
    mat_C[57][1] <=
                mat_A[56][0] * mat_B[1][1] +
                mat_A[56][1] * mat_B[9][1] +
                mat_A[56][2] * mat_B[17][1] +
                mat_A[56][3] * mat_B[25][1] +
                mat_A[57][0] * mat_B[33][1] +
                mat_A[57][1] * mat_B[41][1] +
                mat_A[57][2] * mat_B[49][1] +
                mat_A[57][3] * mat_B[57][1] +
                mat_A[58][0] * mat_B[65][1] +
                mat_A[58][1] * mat_B[73][1] +
                mat_A[58][2] * mat_B[81][1] +
                mat_A[58][3] * mat_B[89][1] +
                mat_A[59][0] * mat_B[97][1] +
                mat_A[59][1] * mat_B[105][1] +
                mat_A[59][2] * mat_B[113][1] +
                mat_A[59][3] * mat_B[121][1] +
                mat_A[60][0] * mat_B[129][1] +
                mat_A[60][1] * mat_B[137][1] +
                mat_A[60][2] * mat_B[145][1] +
                mat_A[60][3] * mat_B[153][1] +
                mat_A[61][0] * mat_B[161][1] +
                mat_A[61][1] * mat_B[169][1] +
                mat_A[61][2] * mat_B[177][1] +
                mat_A[61][3] * mat_B[185][1] +
                mat_A[62][0] * mat_B[193][1] +
                mat_A[62][1] * mat_B[201][1] +
                mat_A[62][2] * mat_B[209][1] +
                mat_A[62][3] * mat_B[217][1] +
                mat_A[63][0] * mat_B[225][1] +
                mat_A[63][1] * mat_B[233][1] +
                mat_A[63][2] * mat_B[241][1] +
                mat_A[63][3] * mat_B[249][1];
    mat_C[57][2] <=
                mat_A[56][0] * mat_B[1][2] +
                mat_A[56][1] * mat_B[9][2] +
                mat_A[56][2] * mat_B[17][2] +
                mat_A[56][3] * mat_B[25][2] +
                mat_A[57][0] * mat_B[33][2] +
                mat_A[57][1] * mat_B[41][2] +
                mat_A[57][2] * mat_B[49][2] +
                mat_A[57][3] * mat_B[57][2] +
                mat_A[58][0] * mat_B[65][2] +
                mat_A[58][1] * mat_B[73][2] +
                mat_A[58][2] * mat_B[81][2] +
                mat_A[58][3] * mat_B[89][2] +
                mat_A[59][0] * mat_B[97][2] +
                mat_A[59][1] * mat_B[105][2] +
                mat_A[59][2] * mat_B[113][2] +
                mat_A[59][3] * mat_B[121][2] +
                mat_A[60][0] * mat_B[129][2] +
                mat_A[60][1] * mat_B[137][2] +
                mat_A[60][2] * mat_B[145][2] +
                mat_A[60][3] * mat_B[153][2] +
                mat_A[61][0] * mat_B[161][2] +
                mat_A[61][1] * mat_B[169][2] +
                mat_A[61][2] * mat_B[177][2] +
                mat_A[61][3] * mat_B[185][2] +
                mat_A[62][0] * mat_B[193][2] +
                mat_A[62][1] * mat_B[201][2] +
                mat_A[62][2] * mat_B[209][2] +
                mat_A[62][3] * mat_B[217][2] +
                mat_A[63][0] * mat_B[225][2] +
                mat_A[63][1] * mat_B[233][2] +
                mat_A[63][2] * mat_B[241][2] +
                mat_A[63][3] * mat_B[249][2];
    mat_C[57][3] <=
                mat_A[56][0] * mat_B[1][3] +
                mat_A[56][1] * mat_B[9][3] +
                mat_A[56][2] * mat_B[17][3] +
                mat_A[56][3] * mat_B[25][3] +
                mat_A[57][0] * mat_B[33][3] +
                mat_A[57][1] * mat_B[41][3] +
                mat_A[57][2] * mat_B[49][3] +
                mat_A[57][3] * mat_B[57][3] +
                mat_A[58][0] * mat_B[65][3] +
                mat_A[58][1] * mat_B[73][3] +
                mat_A[58][2] * mat_B[81][3] +
                mat_A[58][3] * mat_B[89][3] +
                mat_A[59][0] * mat_B[97][3] +
                mat_A[59][1] * mat_B[105][3] +
                mat_A[59][2] * mat_B[113][3] +
                mat_A[59][3] * mat_B[121][3] +
                mat_A[60][0] * mat_B[129][3] +
                mat_A[60][1] * mat_B[137][3] +
                mat_A[60][2] * mat_B[145][3] +
                mat_A[60][3] * mat_B[153][3] +
                mat_A[61][0] * mat_B[161][3] +
                mat_A[61][1] * mat_B[169][3] +
                mat_A[61][2] * mat_B[177][3] +
                mat_A[61][3] * mat_B[185][3] +
                mat_A[62][0] * mat_B[193][3] +
                mat_A[62][1] * mat_B[201][3] +
                mat_A[62][2] * mat_B[209][3] +
                mat_A[62][3] * mat_B[217][3] +
                mat_A[63][0] * mat_B[225][3] +
                mat_A[63][1] * mat_B[233][3] +
                mat_A[63][2] * mat_B[241][3] +
                mat_A[63][3] * mat_B[249][3];
    mat_C[58][0] <=
                mat_A[56][0] * mat_B[2][0] +
                mat_A[56][1] * mat_B[10][0] +
                mat_A[56][2] * mat_B[18][0] +
                mat_A[56][3] * mat_B[26][0] +
                mat_A[57][0] * mat_B[34][0] +
                mat_A[57][1] * mat_B[42][0] +
                mat_A[57][2] * mat_B[50][0] +
                mat_A[57][3] * mat_B[58][0] +
                mat_A[58][0] * mat_B[66][0] +
                mat_A[58][1] * mat_B[74][0] +
                mat_A[58][2] * mat_B[82][0] +
                mat_A[58][3] * mat_B[90][0] +
                mat_A[59][0] * mat_B[98][0] +
                mat_A[59][1] * mat_B[106][0] +
                mat_A[59][2] * mat_B[114][0] +
                mat_A[59][3] * mat_B[122][0] +
                mat_A[60][0] * mat_B[130][0] +
                mat_A[60][1] * mat_B[138][0] +
                mat_A[60][2] * mat_B[146][0] +
                mat_A[60][3] * mat_B[154][0] +
                mat_A[61][0] * mat_B[162][0] +
                mat_A[61][1] * mat_B[170][0] +
                mat_A[61][2] * mat_B[178][0] +
                mat_A[61][3] * mat_B[186][0] +
                mat_A[62][0] * mat_B[194][0] +
                mat_A[62][1] * mat_B[202][0] +
                mat_A[62][2] * mat_B[210][0] +
                mat_A[62][3] * mat_B[218][0] +
                mat_A[63][0] * mat_B[226][0] +
                mat_A[63][1] * mat_B[234][0] +
                mat_A[63][2] * mat_B[242][0] +
                mat_A[63][3] * mat_B[250][0];
    mat_C[58][1] <=
                mat_A[56][0] * mat_B[2][1] +
                mat_A[56][1] * mat_B[10][1] +
                mat_A[56][2] * mat_B[18][1] +
                mat_A[56][3] * mat_B[26][1] +
                mat_A[57][0] * mat_B[34][1] +
                mat_A[57][1] * mat_B[42][1] +
                mat_A[57][2] * mat_B[50][1] +
                mat_A[57][3] * mat_B[58][1] +
                mat_A[58][0] * mat_B[66][1] +
                mat_A[58][1] * mat_B[74][1] +
                mat_A[58][2] * mat_B[82][1] +
                mat_A[58][3] * mat_B[90][1] +
                mat_A[59][0] * mat_B[98][1] +
                mat_A[59][1] * mat_B[106][1] +
                mat_A[59][2] * mat_B[114][1] +
                mat_A[59][3] * mat_B[122][1] +
                mat_A[60][0] * mat_B[130][1] +
                mat_A[60][1] * mat_B[138][1] +
                mat_A[60][2] * mat_B[146][1] +
                mat_A[60][3] * mat_B[154][1] +
                mat_A[61][0] * mat_B[162][1] +
                mat_A[61][1] * mat_B[170][1] +
                mat_A[61][2] * mat_B[178][1] +
                mat_A[61][3] * mat_B[186][1] +
                mat_A[62][0] * mat_B[194][1] +
                mat_A[62][1] * mat_B[202][1] +
                mat_A[62][2] * mat_B[210][1] +
                mat_A[62][3] * mat_B[218][1] +
                mat_A[63][0] * mat_B[226][1] +
                mat_A[63][1] * mat_B[234][1] +
                mat_A[63][2] * mat_B[242][1] +
                mat_A[63][3] * mat_B[250][1];
    mat_C[58][2] <=
                mat_A[56][0] * mat_B[2][2] +
                mat_A[56][1] * mat_B[10][2] +
                mat_A[56][2] * mat_B[18][2] +
                mat_A[56][3] * mat_B[26][2] +
                mat_A[57][0] * mat_B[34][2] +
                mat_A[57][1] * mat_B[42][2] +
                mat_A[57][2] * mat_B[50][2] +
                mat_A[57][3] * mat_B[58][2] +
                mat_A[58][0] * mat_B[66][2] +
                mat_A[58][1] * mat_B[74][2] +
                mat_A[58][2] * mat_B[82][2] +
                mat_A[58][3] * mat_B[90][2] +
                mat_A[59][0] * mat_B[98][2] +
                mat_A[59][1] * mat_B[106][2] +
                mat_A[59][2] * mat_B[114][2] +
                mat_A[59][3] * mat_B[122][2] +
                mat_A[60][0] * mat_B[130][2] +
                mat_A[60][1] * mat_B[138][2] +
                mat_A[60][2] * mat_B[146][2] +
                mat_A[60][3] * mat_B[154][2] +
                mat_A[61][0] * mat_B[162][2] +
                mat_A[61][1] * mat_B[170][2] +
                mat_A[61][2] * mat_B[178][2] +
                mat_A[61][3] * mat_B[186][2] +
                mat_A[62][0] * mat_B[194][2] +
                mat_A[62][1] * mat_B[202][2] +
                mat_A[62][2] * mat_B[210][2] +
                mat_A[62][3] * mat_B[218][2] +
                mat_A[63][0] * mat_B[226][2] +
                mat_A[63][1] * mat_B[234][2] +
                mat_A[63][2] * mat_B[242][2] +
                mat_A[63][3] * mat_B[250][2];
    mat_C[58][3] <=
                mat_A[56][0] * mat_B[2][3] +
                mat_A[56][1] * mat_B[10][3] +
                mat_A[56][2] * mat_B[18][3] +
                mat_A[56][3] * mat_B[26][3] +
                mat_A[57][0] * mat_B[34][3] +
                mat_A[57][1] * mat_B[42][3] +
                mat_A[57][2] * mat_B[50][3] +
                mat_A[57][3] * mat_B[58][3] +
                mat_A[58][0] * mat_B[66][3] +
                mat_A[58][1] * mat_B[74][3] +
                mat_A[58][2] * mat_B[82][3] +
                mat_A[58][3] * mat_B[90][3] +
                mat_A[59][0] * mat_B[98][3] +
                mat_A[59][1] * mat_B[106][3] +
                mat_A[59][2] * mat_B[114][3] +
                mat_A[59][3] * mat_B[122][3] +
                mat_A[60][0] * mat_B[130][3] +
                mat_A[60][1] * mat_B[138][3] +
                mat_A[60][2] * mat_B[146][3] +
                mat_A[60][3] * mat_B[154][3] +
                mat_A[61][0] * mat_B[162][3] +
                mat_A[61][1] * mat_B[170][3] +
                mat_A[61][2] * mat_B[178][3] +
                mat_A[61][3] * mat_B[186][3] +
                mat_A[62][0] * mat_B[194][3] +
                mat_A[62][1] * mat_B[202][3] +
                mat_A[62][2] * mat_B[210][3] +
                mat_A[62][3] * mat_B[218][3] +
                mat_A[63][0] * mat_B[226][3] +
                mat_A[63][1] * mat_B[234][3] +
                mat_A[63][2] * mat_B[242][3] +
                mat_A[63][3] * mat_B[250][3];
    mat_C[59][0] <=
                mat_A[56][0] * mat_B[3][0] +
                mat_A[56][1] * mat_B[11][0] +
                mat_A[56][2] * mat_B[19][0] +
                mat_A[56][3] * mat_B[27][0] +
                mat_A[57][0] * mat_B[35][0] +
                mat_A[57][1] * mat_B[43][0] +
                mat_A[57][2] * mat_B[51][0] +
                mat_A[57][3] * mat_B[59][0] +
                mat_A[58][0] * mat_B[67][0] +
                mat_A[58][1] * mat_B[75][0] +
                mat_A[58][2] * mat_B[83][0] +
                mat_A[58][3] * mat_B[91][0] +
                mat_A[59][0] * mat_B[99][0] +
                mat_A[59][1] * mat_B[107][0] +
                mat_A[59][2] * mat_B[115][0] +
                mat_A[59][3] * mat_B[123][0] +
                mat_A[60][0] * mat_B[131][0] +
                mat_A[60][1] * mat_B[139][0] +
                mat_A[60][2] * mat_B[147][0] +
                mat_A[60][3] * mat_B[155][0] +
                mat_A[61][0] * mat_B[163][0] +
                mat_A[61][1] * mat_B[171][0] +
                mat_A[61][2] * mat_B[179][0] +
                mat_A[61][3] * mat_B[187][0] +
                mat_A[62][0] * mat_B[195][0] +
                mat_A[62][1] * mat_B[203][0] +
                mat_A[62][2] * mat_B[211][0] +
                mat_A[62][3] * mat_B[219][0] +
                mat_A[63][0] * mat_B[227][0] +
                mat_A[63][1] * mat_B[235][0] +
                mat_A[63][2] * mat_B[243][0] +
                mat_A[63][3] * mat_B[251][0];
    mat_C[59][1] <=
                mat_A[56][0] * mat_B[3][1] +
                mat_A[56][1] * mat_B[11][1] +
                mat_A[56][2] * mat_B[19][1] +
                mat_A[56][3] * mat_B[27][1] +
                mat_A[57][0] * mat_B[35][1] +
                mat_A[57][1] * mat_B[43][1] +
                mat_A[57][2] * mat_B[51][1] +
                mat_A[57][3] * mat_B[59][1] +
                mat_A[58][0] * mat_B[67][1] +
                mat_A[58][1] * mat_B[75][1] +
                mat_A[58][2] * mat_B[83][1] +
                mat_A[58][3] * mat_B[91][1] +
                mat_A[59][0] * mat_B[99][1] +
                mat_A[59][1] * mat_B[107][1] +
                mat_A[59][2] * mat_B[115][1] +
                mat_A[59][3] * mat_B[123][1] +
                mat_A[60][0] * mat_B[131][1] +
                mat_A[60][1] * mat_B[139][1] +
                mat_A[60][2] * mat_B[147][1] +
                mat_A[60][3] * mat_B[155][1] +
                mat_A[61][0] * mat_B[163][1] +
                mat_A[61][1] * mat_B[171][1] +
                mat_A[61][2] * mat_B[179][1] +
                mat_A[61][3] * mat_B[187][1] +
                mat_A[62][0] * mat_B[195][1] +
                mat_A[62][1] * mat_B[203][1] +
                mat_A[62][2] * mat_B[211][1] +
                mat_A[62][3] * mat_B[219][1] +
                mat_A[63][0] * mat_B[227][1] +
                mat_A[63][1] * mat_B[235][1] +
                mat_A[63][2] * mat_B[243][1] +
                mat_A[63][3] * mat_B[251][1];
    mat_C[59][2] <=
                mat_A[56][0] * mat_B[3][2] +
                mat_A[56][1] * mat_B[11][2] +
                mat_A[56][2] * mat_B[19][2] +
                mat_A[56][3] * mat_B[27][2] +
                mat_A[57][0] * mat_B[35][2] +
                mat_A[57][1] * mat_B[43][2] +
                mat_A[57][2] * mat_B[51][2] +
                mat_A[57][3] * mat_B[59][2] +
                mat_A[58][0] * mat_B[67][2] +
                mat_A[58][1] * mat_B[75][2] +
                mat_A[58][2] * mat_B[83][2] +
                mat_A[58][3] * mat_B[91][2] +
                mat_A[59][0] * mat_B[99][2] +
                mat_A[59][1] * mat_B[107][2] +
                mat_A[59][2] * mat_B[115][2] +
                mat_A[59][3] * mat_B[123][2] +
                mat_A[60][0] * mat_B[131][2] +
                mat_A[60][1] * mat_B[139][2] +
                mat_A[60][2] * mat_B[147][2] +
                mat_A[60][3] * mat_B[155][2] +
                mat_A[61][0] * mat_B[163][2] +
                mat_A[61][1] * mat_B[171][2] +
                mat_A[61][2] * mat_B[179][2] +
                mat_A[61][3] * mat_B[187][2] +
                mat_A[62][0] * mat_B[195][2] +
                mat_A[62][1] * mat_B[203][2] +
                mat_A[62][2] * mat_B[211][2] +
                mat_A[62][3] * mat_B[219][2] +
                mat_A[63][0] * mat_B[227][2] +
                mat_A[63][1] * mat_B[235][2] +
                mat_A[63][2] * mat_B[243][2] +
                mat_A[63][3] * mat_B[251][2];
    mat_C[59][3] <=
                mat_A[56][0] * mat_B[3][3] +
                mat_A[56][1] * mat_B[11][3] +
                mat_A[56][2] * mat_B[19][3] +
                mat_A[56][3] * mat_B[27][3] +
                mat_A[57][0] * mat_B[35][3] +
                mat_A[57][1] * mat_B[43][3] +
                mat_A[57][2] * mat_B[51][3] +
                mat_A[57][3] * mat_B[59][3] +
                mat_A[58][0] * mat_B[67][3] +
                mat_A[58][1] * mat_B[75][3] +
                mat_A[58][2] * mat_B[83][3] +
                mat_A[58][3] * mat_B[91][3] +
                mat_A[59][0] * mat_B[99][3] +
                mat_A[59][1] * mat_B[107][3] +
                mat_A[59][2] * mat_B[115][3] +
                mat_A[59][3] * mat_B[123][3] +
                mat_A[60][0] * mat_B[131][3] +
                mat_A[60][1] * mat_B[139][3] +
                mat_A[60][2] * mat_B[147][3] +
                mat_A[60][3] * mat_B[155][3] +
                mat_A[61][0] * mat_B[163][3] +
                mat_A[61][1] * mat_B[171][3] +
                mat_A[61][2] * mat_B[179][3] +
                mat_A[61][3] * mat_B[187][3] +
                mat_A[62][0] * mat_B[195][3] +
                mat_A[62][1] * mat_B[203][3] +
                mat_A[62][2] * mat_B[211][3] +
                mat_A[62][3] * mat_B[219][3] +
                mat_A[63][0] * mat_B[227][3] +
                mat_A[63][1] * mat_B[235][3] +
                mat_A[63][2] * mat_B[243][3] +
                mat_A[63][3] * mat_B[251][3];
    mat_C[60][0] <=
                mat_A[56][0] * mat_B[4][0] +
                mat_A[56][1] * mat_B[12][0] +
                mat_A[56][2] * mat_B[20][0] +
                mat_A[56][3] * mat_B[28][0] +
                mat_A[57][0] * mat_B[36][0] +
                mat_A[57][1] * mat_B[44][0] +
                mat_A[57][2] * mat_B[52][0] +
                mat_A[57][3] * mat_B[60][0] +
                mat_A[58][0] * mat_B[68][0] +
                mat_A[58][1] * mat_B[76][0] +
                mat_A[58][2] * mat_B[84][0] +
                mat_A[58][3] * mat_B[92][0] +
                mat_A[59][0] * mat_B[100][0] +
                mat_A[59][1] * mat_B[108][0] +
                mat_A[59][2] * mat_B[116][0] +
                mat_A[59][3] * mat_B[124][0] +
                mat_A[60][0] * mat_B[132][0] +
                mat_A[60][1] * mat_B[140][0] +
                mat_A[60][2] * mat_B[148][0] +
                mat_A[60][3] * mat_B[156][0] +
                mat_A[61][0] * mat_B[164][0] +
                mat_A[61][1] * mat_B[172][0] +
                mat_A[61][2] * mat_B[180][0] +
                mat_A[61][3] * mat_B[188][0] +
                mat_A[62][0] * mat_B[196][0] +
                mat_A[62][1] * mat_B[204][0] +
                mat_A[62][2] * mat_B[212][0] +
                mat_A[62][3] * mat_B[220][0] +
                mat_A[63][0] * mat_B[228][0] +
                mat_A[63][1] * mat_B[236][0] +
                mat_A[63][2] * mat_B[244][0] +
                mat_A[63][3] * mat_B[252][0];
    mat_C[60][1] <=
                mat_A[56][0] * mat_B[4][1] +
                mat_A[56][1] * mat_B[12][1] +
                mat_A[56][2] * mat_B[20][1] +
                mat_A[56][3] * mat_B[28][1] +
                mat_A[57][0] * mat_B[36][1] +
                mat_A[57][1] * mat_B[44][1] +
                mat_A[57][2] * mat_B[52][1] +
                mat_A[57][3] * mat_B[60][1] +
                mat_A[58][0] * mat_B[68][1] +
                mat_A[58][1] * mat_B[76][1] +
                mat_A[58][2] * mat_B[84][1] +
                mat_A[58][3] * mat_B[92][1] +
                mat_A[59][0] * mat_B[100][1] +
                mat_A[59][1] * mat_B[108][1] +
                mat_A[59][2] * mat_B[116][1] +
                mat_A[59][3] * mat_B[124][1] +
                mat_A[60][0] * mat_B[132][1] +
                mat_A[60][1] * mat_B[140][1] +
                mat_A[60][2] * mat_B[148][1] +
                mat_A[60][3] * mat_B[156][1] +
                mat_A[61][0] * mat_B[164][1] +
                mat_A[61][1] * mat_B[172][1] +
                mat_A[61][2] * mat_B[180][1] +
                mat_A[61][3] * mat_B[188][1] +
                mat_A[62][0] * mat_B[196][1] +
                mat_A[62][1] * mat_B[204][1] +
                mat_A[62][2] * mat_B[212][1] +
                mat_A[62][3] * mat_B[220][1] +
                mat_A[63][0] * mat_B[228][1] +
                mat_A[63][1] * mat_B[236][1] +
                mat_A[63][2] * mat_B[244][1] +
                mat_A[63][3] * mat_B[252][1];
    mat_C[60][2] <=
                mat_A[56][0] * mat_B[4][2] +
                mat_A[56][1] * mat_B[12][2] +
                mat_A[56][2] * mat_B[20][2] +
                mat_A[56][3] * mat_B[28][2] +
                mat_A[57][0] * mat_B[36][2] +
                mat_A[57][1] * mat_B[44][2] +
                mat_A[57][2] * mat_B[52][2] +
                mat_A[57][3] * mat_B[60][2] +
                mat_A[58][0] * mat_B[68][2] +
                mat_A[58][1] * mat_B[76][2] +
                mat_A[58][2] * mat_B[84][2] +
                mat_A[58][3] * mat_B[92][2] +
                mat_A[59][0] * mat_B[100][2] +
                mat_A[59][1] * mat_B[108][2] +
                mat_A[59][2] * mat_B[116][2] +
                mat_A[59][3] * mat_B[124][2] +
                mat_A[60][0] * mat_B[132][2] +
                mat_A[60][1] * mat_B[140][2] +
                mat_A[60][2] * mat_B[148][2] +
                mat_A[60][3] * mat_B[156][2] +
                mat_A[61][0] * mat_B[164][2] +
                mat_A[61][1] * mat_B[172][2] +
                mat_A[61][2] * mat_B[180][2] +
                mat_A[61][3] * mat_B[188][2] +
                mat_A[62][0] * mat_B[196][2] +
                mat_A[62][1] * mat_B[204][2] +
                mat_A[62][2] * mat_B[212][2] +
                mat_A[62][3] * mat_B[220][2] +
                mat_A[63][0] * mat_B[228][2] +
                mat_A[63][1] * mat_B[236][2] +
                mat_A[63][2] * mat_B[244][2] +
                mat_A[63][3] * mat_B[252][2];
    mat_C[60][3] <=
                mat_A[56][0] * mat_B[4][3] +
                mat_A[56][1] * mat_B[12][3] +
                mat_A[56][2] * mat_B[20][3] +
                mat_A[56][3] * mat_B[28][3] +
                mat_A[57][0] * mat_B[36][3] +
                mat_A[57][1] * mat_B[44][3] +
                mat_A[57][2] * mat_B[52][3] +
                mat_A[57][3] * mat_B[60][3] +
                mat_A[58][0] * mat_B[68][3] +
                mat_A[58][1] * mat_B[76][3] +
                mat_A[58][2] * mat_B[84][3] +
                mat_A[58][3] * mat_B[92][3] +
                mat_A[59][0] * mat_B[100][3] +
                mat_A[59][1] * mat_B[108][3] +
                mat_A[59][2] * mat_B[116][3] +
                mat_A[59][3] * mat_B[124][3] +
                mat_A[60][0] * mat_B[132][3] +
                mat_A[60][1] * mat_B[140][3] +
                mat_A[60][2] * mat_B[148][3] +
                mat_A[60][3] * mat_B[156][3] +
                mat_A[61][0] * mat_B[164][3] +
                mat_A[61][1] * mat_B[172][3] +
                mat_A[61][2] * mat_B[180][3] +
                mat_A[61][3] * mat_B[188][3] +
                mat_A[62][0] * mat_B[196][3] +
                mat_A[62][1] * mat_B[204][3] +
                mat_A[62][2] * mat_B[212][3] +
                mat_A[62][3] * mat_B[220][3] +
                mat_A[63][0] * mat_B[228][3] +
                mat_A[63][1] * mat_B[236][3] +
                mat_A[63][2] * mat_B[244][3] +
                mat_A[63][3] * mat_B[252][3];
    mat_C[61][0] <=
                mat_A[56][0] * mat_B[5][0] +
                mat_A[56][1] * mat_B[13][0] +
                mat_A[56][2] * mat_B[21][0] +
                mat_A[56][3] * mat_B[29][0] +
                mat_A[57][0] * mat_B[37][0] +
                mat_A[57][1] * mat_B[45][0] +
                mat_A[57][2] * mat_B[53][0] +
                mat_A[57][3] * mat_B[61][0] +
                mat_A[58][0] * mat_B[69][0] +
                mat_A[58][1] * mat_B[77][0] +
                mat_A[58][2] * mat_B[85][0] +
                mat_A[58][3] * mat_B[93][0] +
                mat_A[59][0] * mat_B[101][0] +
                mat_A[59][1] * mat_B[109][0] +
                mat_A[59][2] * mat_B[117][0] +
                mat_A[59][3] * mat_B[125][0] +
                mat_A[60][0] * mat_B[133][0] +
                mat_A[60][1] * mat_B[141][0] +
                mat_A[60][2] * mat_B[149][0] +
                mat_A[60][3] * mat_B[157][0] +
                mat_A[61][0] * mat_B[165][0] +
                mat_A[61][1] * mat_B[173][0] +
                mat_A[61][2] * mat_B[181][0] +
                mat_A[61][3] * mat_B[189][0] +
                mat_A[62][0] * mat_B[197][0] +
                mat_A[62][1] * mat_B[205][0] +
                mat_A[62][2] * mat_B[213][0] +
                mat_A[62][3] * mat_B[221][0] +
                mat_A[63][0] * mat_B[229][0] +
                mat_A[63][1] * mat_B[237][0] +
                mat_A[63][2] * mat_B[245][0] +
                mat_A[63][3] * mat_B[253][0];
    mat_C[61][1] <=
                mat_A[56][0] * mat_B[5][1] +
                mat_A[56][1] * mat_B[13][1] +
                mat_A[56][2] * mat_B[21][1] +
                mat_A[56][3] * mat_B[29][1] +
                mat_A[57][0] * mat_B[37][1] +
                mat_A[57][1] * mat_B[45][1] +
                mat_A[57][2] * mat_B[53][1] +
                mat_A[57][3] * mat_B[61][1] +
                mat_A[58][0] * mat_B[69][1] +
                mat_A[58][1] * mat_B[77][1] +
                mat_A[58][2] * mat_B[85][1] +
                mat_A[58][3] * mat_B[93][1] +
                mat_A[59][0] * mat_B[101][1] +
                mat_A[59][1] * mat_B[109][1] +
                mat_A[59][2] * mat_B[117][1] +
                mat_A[59][3] * mat_B[125][1] +
                mat_A[60][0] * mat_B[133][1] +
                mat_A[60][1] * mat_B[141][1] +
                mat_A[60][2] * mat_B[149][1] +
                mat_A[60][3] * mat_B[157][1] +
                mat_A[61][0] * mat_B[165][1] +
                mat_A[61][1] * mat_B[173][1] +
                mat_A[61][2] * mat_B[181][1] +
                mat_A[61][3] * mat_B[189][1] +
                mat_A[62][0] * mat_B[197][1] +
                mat_A[62][1] * mat_B[205][1] +
                mat_A[62][2] * mat_B[213][1] +
                mat_A[62][3] * mat_B[221][1] +
                mat_A[63][0] * mat_B[229][1] +
                mat_A[63][1] * mat_B[237][1] +
                mat_A[63][2] * mat_B[245][1] +
                mat_A[63][3] * mat_B[253][1];
    mat_C[61][2] <=
                mat_A[56][0] * mat_B[5][2] +
                mat_A[56][1] * mat_B[13][2] +
                mat_A[56][2] * mat_B[21][2] +
                mat_A[56][3] * mat_B[29][2] +
                mat_A[57][0] * mat_B[37][2] +
                mat_A[57][1] * mat_B[45][2] +
                mat_A[57][2] * mat_B[53][2] +
                mat_A[57][3] * mat_B[61][2] +
                mat_A[58][0] * mat_B[69][2] +
                mat_A[58][1] * mat_B[77][2] +
                mat_A[58][2] * mat_B[85][2] +
                mat_A[58][3] * mat_B[93][2] +
                mat_A[59][0] * mat_B[101][2] +
                mat_A[59][1] * mat_B[109][2] +
                mat_A[59][2] * mat_B[117][2] +
                mat_A[59][3] * mat_B[125][2] +
                mat_A[60][0] * mat_B[133][2] +
                mat_A[60][1] * mat_B[141][2] +
                mat_A[60][2] * mat_B[149][2] +
                mat_A[60][3] * mat_B[157][2] +
                mat_A[61][0] * mat_B[165][2] +
                mat_A[61][1] * mat_B[173][2] +
                mat_A[61][2] * mat_B[181][2] +
                mat_A[61][3] * mat_B[189][2] +
                mat_A[62][0] * mat_B[197][2] +
                mat_A[62][1] * mat_B[205][2] +
                mat_A[62][2] * mat_B[213][2] +
                mat_A[62][3] * mat_B[221][2] +
                mat_A[63][0] * mat_B[229][2] +
                mat_A[63][1] * mat_B[237][2] +
                mat_A[63][2] * mat_B[245][2] +
                mat_A[63][3] * mat_B[253][2];
    mat_C[61][3] <=
                mat_A[56][0] * mat_B[5][3] +
                mat_A[56][1] * mat_B[13][3] +
                mat_A[56][2] * mat_B[21][3] +
                mat_A[56][3] * mat_B[29][3] +
                mat_A[57][0] * mat_B[37][3] +
                mat_A[57][1] * mat_B[45][3] +
                mat_A[57][2] * mat_B[53][3] +
                mat_A[57][3] * mat_B[61][3] +
                mat_A[58][0] * mat_B[69][3] +
                mat_A[58][1] * mat_B[77][3] +
                mat_A[58][2] * mat_B[85][3] +
                mat_A[58][3] * mat_B[93][3] +
                mat_A[59][0] * mat_B[101][3] +
                mat_A[59][1] * mat_B[109][3] +
                mat_A[59][2] * mat_B[117][3] +
                mat_A[59][3] * mat_B[125][3] +
                mat_A[60][0] * mat_B[133][3] +
                mat_A[60][1] * mat_B[141][3] +
                mat_A[60][2] * mat_B[149][3] +
                mat_A[60][3] * mat_B[157][3] +
                mat_A[61][0] * mat_B[165][3] +
                mat_A[61][1] * mat_B[173][3] +
                mat_A[61][2] * mat_B[181][3] +
                mat_A[61][3] * mat_B[189][3] +
                mat_A[62][0] * mat_B[197][3] +
                mat_A[62][1] * mat_B[205][3] +
                mat_A[62][2] * mat_B[213][3] +
                mat_A[62][3] * mat_B[221][3] +
                mat_A[63][0] * mat_B[229][3] +
                mat_A[63][1] * mat_B[237][3] +
                mat_A[63][2] * mat_B[245][3] +
                mat_A[63][3] * mat_B[253][3];
    mat_C[62][0] <=
                mat_A[56][0] * mat_B[6][0] +
                mat_A[56][1] * mat_B[14][0] +
                mat_A[56][2] * mat_B[22][0] +
                mat_A[56][3] * mat_B[30][0] +
                mat_A[57][0] * mat_B[38][0] +
                mat_A[57][1] * mat_B[46][0] +
                mat_A[57][2] * mat_B[54][0] +
                mat_A[57][3] * mat_B[62][0] +
                mat_A[58][0] * mat_B[70][0] +
                mat_A[58][1] * mat_B[78][0] +
                mat_A[58][2] * mat_B[86][0] +
                mat_A[58][3] * mat_B[94][0] +
                mat_A[59][0] * mat_B[102][0] +
                mat_A[59][1] * mat_B[110][0] +
                mat_A[59][2] * mat_B[118][0] +
                mat_A[59][3] * mat_B[126][0] +
                mat_A[60][0] * mat_B[134][0] +
                mat_A[60][1] * mat_B[142][0] +
                mat_A[60][2] * mat_B[150][0] +
                mat_A[60][3] * mat_B[158][0] +
                mat_A[61][0] * mat_B[166][0] +
                mat_A[61][1] * mat_B[174][0] +
                mat_A[61][2] * mat_B[182][0] +
                mat_A[61][3] * mat_B[190][0] +
                mat_A[62][0] * mat_B[198][0] +
                mat_A[62][1] * mat_B[206][0] +
                mat_A[62][2] * mat_B[214][0] +
                mat_A[62][3] * mat_B[222][0] +
                mat_A[63][0] * mat_B[230][0] +
                mat_A[63][1] * mat_B[238][0] +
                mat_A[63][2] * mat_B[246][0] +
                mat_A[63][3] * mat_B[254][0];
    mat_C[62][1] <=
                mat_A[56][0] * mat_B[6][1] +
                mat_A[56][1] * mat_B[14][1] +
                mat_A[56][2] * mat_B[22][1] +
                mat_A[56][3] * mat_B[30][1] +
                mat_A[57][0] * mat_B[38][1] +
                mat_A[57][1] * mat_B[46][1] +
                mat_A[57][2] * mat_B[54][1] +
                mat_A[57][3] * mat_B[62][1] +
                mat_A[58][0] * mat_B[70][1] +
                mat_A[58][1] * mat_B[78][1] +
                mat_A[58][2] * mat_B[86][1] +
                mat_A[58][3] * mat_B[94][1] +
                mat_A[59][0] * mat_B[102][1] +
                mat_A[59][1] * mat_B[110][1] +
                mat_A[59][2] * mat_B[118][1] +
                mat_A[59][3] * mat_B[126][1] +
                mat_A[60][0] * mat_B[134][1] +
                mat_A[60][1] * mat_B[142][1] +
                mat_A[60][2] * mat_B[150][1] +
                mat_A[60][3] * mat_B[158][1] +
                mat_A[61][0] * mat_B[166][1] +
                mat_A[61][1] * mat_B[174][1] +
                mat_A[61][2] * mat_B[182][1] +
                mat_A[61][3] * mat_B[190][1] +
                mat_A[62][0] * mat_B[198][1] +
                mat_A[62][1] * mat_B[206][1] +
                mat_A[62][2] * mat_B[214][1] +
                mat_A[62][3] * mat_B[222][1] +
                mat_A[63][0] * mat_B[230][1] +
                mat_A[63][1] * mat_B[238][1] +
                mat_A[63][2] * mat_B[246][1] +
                mat_A[63][3] * mat_B[254][1];
    mat_C[62][2] <=
                mat_A[56][0] * mat_B[6][2] +
                mat_A[56][1] * mat_B[14][2] +
                mat_A[56][2] * mat_B[22][2] +
                mat_A[56][3] * mat_B[30][2] +
                mat_A[57][0] * mat_B[38][2] +
                mat_A[57][1] * mat_B[46][2] +
                mat_A[57][2] * mat_B[54][2] +
                mat_A[57][3] * mat_B[62][2] +
                mat_A[58][0] * mat_B[70][2] +
                mat_A[58][1] * mat_B[78][2] +
                mat_A[58][2] * mat_B[86][2] +
                mat_A[58][3] * mat_B[94][2] +
                mat_A[59][0] * mat_B[102][2] +
                mat_A[59][1] * mat_B[110][2] +
                mat_A[59][2] * mat_B[118][2] +
                mat_A[59][3] * mat_B[126][2] +
                mat_A[60][0] * mat_B[134][2] +
                mat_A[60][1] * mat_B[142][2] +
                mat_A[60][2] * mat_B[150][2] +
                mat_A[60][3] * mat_B[158][2] +
                mat_A[61][0] * mat_B[166][2] +
                mat_A[61][1] * mat_B[174][2] +
                mat_A[61][2] * mat_B[182][2] +
                mat_A[61][3] * mat_B[190][2] +
                mat_A[62][0] * mat_B[198][2] +
                mat_A[62][1] * mat_B[206][2] +
                mat_A[62][2] * mat_B[214][2] +
                mat_A[62][3] * mat_B[222][2] +
                mat_A[63][0] * mat_B[230][2] +
                mat_A[63][1] * mat_B[238][2] +
                mat_A[63][2] * mat_B[246][2] +
                mat_A[63][3] * mat_B[254][2];
    mat_C[62][3] <=
                mat_A[56][0] * mat_B[6][3] +
                mat_A[56][1] * mat_B[14][3] +
                mat_A[56][2] * mat_B[22][3] +
                mat_A[56][3] * mat_B[30][3] +
                mat_A[57][0] * mat_B[38][3] +
                mat_A[57][1] * mat_B[46][3] +
                mat_A[57][2] * mat_B[54][3] +
                mat_A[57][3] * mat_B[62][3] +
                mat_A[58][0] * mat_B[70][3] +
                mat_A[58][1] * mat_B[78][3] +
                mat_A[58][2] * mat_B[86][3] +
                mat_A[58][3] * mat_B[94][3] +
                mat_A[59][0] * mat_B[102][3] +
                mat_A[59][1] * mat_B[110][3] +
                mat_A[59][2] * mat_B[118][3] +
                mat_A[59][3] * mat_B[126][3] +
                mat_A[60][0] * mat_B[134][3] +
                mat_A[60][1] * mat_B[142][3] +
                mat_A[60][2] * mat_B[150][3] +
                mat_A[60][3] * mat_B[158][3] +
                mat_A[61][0] * mat_B[166][3] +
                mat_A[61][1] * mat_B[174][3] +
                mat_A[61][2] * mat_B[182][3] +
                mat_A[61][3] * mat_B[190][3] +
                mat_A[62][0] * mat_B[198][3] +
                mat_A[62][1] * mat_B[206][3] +
                mat_A[62][2] * mat_B[214][3] +
                mat_A[62][3] * mat_B[222][3] +
                mat_A[63][0] * mat_B[230][3] +
                mat_A[63][1] * mat_B[238][3] +
                mat_A[63][2] * mat_B[246][3] +
                mat_A[63][3] * mat_B[254][3];
    mat_C[63][0] <=
                mat_A[56][0] * mat_B[7][0] +
                mat_A[56][1] * mat_B[15][0] +
                mat_A[56][2] * mat_B[23][0] +
                mat_A[56][3] * mat_B[31][0] +
                mat_A[57][0] * mat_B[39][0] +
                mat_A[57][1] * mat_B[47][0] +
                mat_A[57][2] * mat_B[55][0] +
                mat_A[57][3] * mat_B[63][0] +
                mat_A[58][0] * mat_B[71][0] +
                mat_A[58][1] * mat_B[79][0] +
                mat_A[58][2] * mat_B[87][0] +
                mat_A[58][3] * mat_B[95][0] +
                mat_A[59][0] * mat_B[103][0] +
                mat_A[59][1] * mat_B[111][0] +
                mat_A[59][2] * mat_B[119][0] +
                mat_A[59][3] * mat_B[127][0] +
                mat_A[60][0] * mat_B[135][0] +
                mat_A[60][1] * mat_B[143][0] +
                mat_A[60][2] * mat_B[151][0] +
                mat_A[60][3] * mat_B[159][0] +
                mat_A[61][0] * mat_B[167][0] +
                mat_A[61][1] * mat_B[175][0] +
                mat_A[61][2] * mat_B[183][0] +
                mat_A[61][3] * mat_B[191][0] +
                mat_A[62][0] * mat_B[199][0] +
                mat_A[62][1] * mat_B[207][0] +
                mat_A[62][2] * mat_B[215][0] +
                mat_A[62][3] * mat_B[223][0] +
                mat_A[63][0] * mat_B[231][0] +
                mat_A[63][1] * mat_B[239][0] +
                mat_A[63][2] * mat_B[247][0] +
                mat_A[63][3] * mat_B[255][0];
    mat_C[63][1] <=
                mat_A[56][0] * mat_B[7][1] +
                mat_A[56][1] * mat_B[15][1] +
                mat_A[56][2] * mat_B[23][1] +
                mat_A[56][3] * mat_B[31][1] +
                mat_A[57][0] * mat_B[39][1] +
                mat_A[57][1] * mat_B[47][1] +
                mat_A[57][2] * mat_B[55][1] +
                mat_A[57][3] * mat_B[63][1] +
                mat_A[58][0] * mat_B[71][1] +
                mat_A[58][1] * mat_B[79][1] +
                mat_A[58][2] * mat_B[87][1] +
                mat_A[58][3] * mat_B[95][1] +
                mat_A[59][0] * mat_B[103][1] +
                mat_A[59][1] * mat_B[111][1] +
                mat_A[59][2] * mat_B[119][1] +
                mat_A[59][3] * mat_B[127][1] +
                mat_A[60][0] * mat_B[135][1] +
                mat_A[60][1] * mat_B[143][1] +
                mat_A[60][2] * mat_B[151][1] +
                mat_A[60][3] * mat_B[159][1] +
                mat_A[61][0] * mat_B[167][1] +
                mat_A[61][1] * mat_B[175][1] +
                mat_A[61][2] * mat_B[183][1] +
                mat_A[61][3] * mat_B[191][1] +
                mat_A[62][0] * mat_B[199][1] +
                mat_A[62][1] * mat_B[207][1] +
                mat_A[62][2] * mat_B[215][1] +
                mat_A[62][3] * mat_B[223][1] +
                mat_A[63][0] * mat_B[231][1] +
                mat_A[63][1] * mat_B[239][1] +
                mat_A[63][2] * mat_B[247][1] +
                mat_A[63][3] * mat_B[255][1];
    mat_C[63][2] <=
                mat_A[56][0] * mat_B[7][2] +
                mat_A[56][1] * mat_B[15][2] +
                mat_A[56][2] * mat_B[23][2] +
                mat_A[56][3] * mat_B[31][2] +
                mat_A[57][0] * mat_B[39][2] +
                mat_A[57][1] * mat_B[47][2] +
                mat_A[57][2] * mat_B[55][2] +
                mat_A[57][3] * mat_B[63][2] +
                mat_A[58][0] * mat_B[71][2] +
                mat_A[58][1] * mat_B[79][2] +
                mat_A[58][2] * mat_B[87][2] +
                mat_A[58][3] * mat_B[95][2] +
                mat_A[59][0] * mat_B[103][2] +
                mat_A[59][1] * mat_B[111][2] +
                mat_A[59][2] * mat_B[119][2] +
                mat_A[59][3] * mat_B[127][2] +
                mat_A[60][0] * mat_B[135][2] +
                mat_A[60][1] * mat_B[143][2] +
                mat_A[60][2] * mat_B[151][2] +
                mat_A[60][3] * mat_B[159][2] +
                mat_A[61][0] * mat_B[167][2] +
                mat_A[61][1] * mat_B[175][2] +
                mat_A[61][2] * mat_B[183][2] +
                mat_A[61][3] * mat_B[191][2] +
                mat_A[62][0] * mat_B[199][2] +
                mat_A[62][1] * mat_B[207][2] +
                mat_A[62][2] * mat_B[215][2] +
                mat_A[62][3] * mat_B[223][2] +
                mat_A[63][0] * mat_B[231][2] +
                mat_A[63][1] * mat_B[239][2] +
                mat_A[63][2] * mat_B[247][2] +
                mat_A[63][3] * mat_B[255][2];
    mat_C[63][3] <=
                mat_A[56][0] * mat_B[7][3] +
                mat_A[56][1] * mat_B[15][3] +
                mat_A[56][2] * mat_B[23][3] +
                mat_A[56][3] * mat_B[31][3] +
                mat_A[57][0] * mat_B[39][3] +
                mat_A[57][1] * mat_B[47][3] +
                mat_A[57][2] * mat_B[55][3] +
                mat_A[57][3] * mat_B[63][3] +
                mat_A[58][0] * mat_B[71][3] +
                mat_A[58][1] * mat_B[79][3] +
                mat_A[58][2] * mat_B[87][3] +
                mat_A[58][3] * mat_B[95][3] +
                mat_A[59][0] * mat_B[103][3] +
                mat_A[59][1] * mat_B[111][3] +
                mat_A[59][2] * mat_B[119][3] +
                mat_A[59][3] * mat_B[127][3] +
                mat_A[60][0] * mat_B[135][3] +
                mat_A[60][1] * mat_B[143][3] +
                mat_A[60][2] * mat_B[151][3] +
                mat_A[60][3] * mat_B[159][3] +
                mat_A[61][0] * mat_B[167][3] +
                mat_A[61][1] * mat_B[175][3] +
                mat_A[61][2] * mat_B[183][3] +
                mat_A[61][3] * mat_B[191][3] +
                mat_A[62][0] * mat_B[199][3] +
                mat_A[62][1] * mat_B[207][3] +
                mat_A[62][2] * mat_B[215][3] +
                mat_A[62][3] * mat_B[223][3] +
                mat_A[63][0] * mat_B[231][3] +
                mat_A[63][1] * mat_B[239][3] +
                mat_A[63][2] * mat_B[247][3] +
                mat_A[63][3] * mat_B[255][3];
    mat_C[64][0] <=
                mat_A[64][0] * mat_B[0][0] +
                mat_A[64][1] * mat_B[8][0] +
                mat_A[64][2] * mat_B[16][0] +
                mat_A[64][3] * mat_B[24][0] +
                mat_A[65][0] * mat_B[32][0] +
                mat_A[65][1] * mat_B[40][0] +
                mat_A[65][2] * mat_B[48][0] +
                mat_A[65][3] * mat_B[56][0] +
                mat_A[66][0] * mat_B[64][0] +
                mat_A[66][1] * mat_B[72][0] +
                mat_A[66][2] * mat_B[80][0] +
                mat_A[66][3] * mat_B[88][0] +
                mat_A[67][0] * mat_B[96][0] +
                mat_A[67][1] * mat_B[104][0] +
                mat_A[67][2] * mat_B[112][0] +
                mat_A[67][3] * mat_B[120][0] +
                mat_A[68][0] * mat_B[128][0] +
                mat_A[68][1] * mat_B[136][0] +
                mat_A[68][2] * mat_B[144][0] +
                mat_A[68][3] * mat_B[152][0] +
                mat_A[69][0] * mat_B[160][0] +
                mat_A[69][1] * mat_B[168][0] +
                mat_A[69][2] * mat_B[176][0] +
                mat_A[69][3] * mat_B[184][0] +
                mat_A[70][0] * mat_B[192][0] +
                mat_A[70][1] * mat_B[200][0] +
                mat_A[70][2] * mat_B[208][0] +
                mat_A[70][3] * mat_B[216][0] +
                mat_A[71][0] * mat_B[224][0] +
                mat_A[71][1] * mat_B[232][0] +
                mat_A[71][2] * mat_B[240][0] +
                mat_A[71][3] * mat_B[248][0];
    mat_C[64][1] <=
                mat_A[64][0] * mat_B[0][1] +
                mat_A[64][1] * mat_B[8][1] +
                mat_A[64][2] * mat_B[16][1] +
                mat_A[64][3] * mat_B[24][1] +
                mat_A[65][0] * mat_B[32][1] +
                mat_A[65][1] * mat_B[40][1] +
                mat_A[65][2] * mat_B[48][1] +
                mat_A[65][3] * mat_B[56][1] +
                mat_A[66][0] * mat_B[64][1] +
                mat_A[66][1] * mat_B[72][1] +
                mat_A[66][2] * mat_B[80][1] +
                mat_A[66][3] * mat_B[88][1] +
                mat_A[67][0] * mat_B[96][1] +
                mat_A[67][1] * mat_B[104][1] +
                mat_A[67][2] * mat_B[112][1] +
                mat_A[67][3] * mat_B[120][1] +
                mat_A[68][0] * mat_B[128][1] +
                mat_A[68][1] * mat_B[136][1] +
                mat_A[68][2] * mat_B[144][1] +
                mat_A[68][3] * mat_B[152][1] +
                mat_A[69][0] * mat_B[160][1] +
                mat_A[69][1] * mat_B[168][1] +
                mat_A[69][2] * mat_B[176][1] +
                mat_A[69][3] * mat_B[184][1] +
                mat_A[70][0] * mat_B[192][1] +
                mat_A[70][1] * mat_B[200][1] +
                mat_A[70][2] * mat_B[208][1] +
                mat_A[70][3] * mat_B[216][1] +
                mat_A[71][0] * mat_B[224][1] +
                mat_A[71][1] * mat_B[232][1] +
                mat_A[71][2] * mat_B[240][1] +
                mat_A[71][3] * mat_B[248][1];
    mat_C[64][2] <=
                mat_A[64][0] * mat_B[0][2] +
                mat_A[64][1] * mat_B[8][2] +
                mat_A[64][2] * mat_B[16][2] +
                mat_A[64][3] * mat_B[24][2] +
                mat_A[65][0] * mat_B[32][2] +
                mat_A[65][1] * mat_B[40][2] +
                mat_A[65][2] * mat_B[48][2] +
                mat_A[65][3] * mat_B[56][2] +
                mat_A[66][0] * mat_B[64][2] +
                mat_A[66][1] * mat_B[72][2] +
                mat_A[66][2] * mat_B[80][2] +
                mat_A[66][3] * mat_B[88][2] +
                mat_A[67][0] * mat_B[96][2] +
                mat_A[67][1] * mat_B[104][2] +
                mat_A[67][2] * mat_B[112][2] +
                mat_A[67][3] * mat_B[120][2] +
                mat_A[68][0] * mat_B[128][2] +
                mat_A[68][1] * mat_B[136][2] +
                mat_A[68][2] * mat_B[144][2] +
                mat_A[68][3] * mat_B[152][2] +
                mat_A[69][0] * mat_B[160][2] +
                mat_A[69][1] * mat_B[168][2] +
                mat_A[69][2] * mat_B[176][2] +
                mat_A[69][3] * mat_B[184][2] +
                mat_A[70][0] * mat_B[192][2] +
                mat_A[70][1] * mat_B[200][2] +
                mat_A[70][2] * mat_B[208][2] +
                mat_A[70][3] * mat_B[216][2] +
                mat_A[71][0] * mat_B[224][2] +
                mat_A[71][1] * mat_B[232][2] +
                mat_A[71][2] * mat_B[240][2] +
                mat_A[71][3] * mat_B[248][2];
    mat_C[64][3] <=
                mat_A[64][0] * mat_B[0][3] +
                mat_A[64][1] * mat_B[8][3] +
                mat_A[64][2] * mat_B[16][3] +
                mat_A[64][3] * mat_B[24][3] +
                mat_A[65][0] * mat_B[32][3] +
                mat_A[65][1] * mat_B[40][3] +
                mat_A[65][2] * mat_B[48][3] +
                mat_A[65][3] * mat_B[56][3] +
                mat_A[66][0] * mat_B[64][3] +
                mat_A[66][1] * mat_B[72][3] +
                mat_A[66][2] * mat_B[80][3] +
                mat_A[66][3] * mat_B[88][3] +
                mat_A[67][0] * mat_B[96][3] +
                mat_A[67][1] * mat_B[104][3] +
                mat_A[67][2] * mat_B[112][3] +
                mat_A[67][3] * mat_B[120][3] +
                mat_A[68][0] * mat_B[128][3] +
                mat_A[68][1] * mat_B[136][3] +
                mat_A[68][2] * mat_B[144][3] +
                mat_A[68][3] * mat_B[152][3] +
                mat_A[69][0] * mat_B[160][3] +
                mat_A[69][1] * mat_B[168][3] +
                mat_A[69][2] * mat_B[176][3] +
                mat_A[69][3] * mat_B[184][3] +
                mat_A[70][0] * mat_B[192][3] +
                mat_A[70][1] * mat_B[200][3] +
                mat_A[70][2] * mat_B[208][3] +
                mat_A[70][3] * mat_B[216][3] +
                mat_A[71][0] * mat_B[224][3] +
                mat_A[71][1] * mat_B[232][3] +
                mat_A[71][2] * mat_B[240][3] +
                mat_A[71][3] * mat_B[248][3];
    mat_C[65][0] <=
                mat_A[64][0] * mat_B[1][0] +
                mat_A[64][1] * mat_B[9][0] +
                mat_A[64][2] * mat_B[17][0] +
                mat_A[64][3] * mat_B[25][0] +
                mat_A[65][0] * mat_B[33][0] +
                mat_A[65][1] * mat_B[41][0] +
                mat_A[65][2] * mat_B[49][0] +
                mat_A[65][3] * mat_B[57][0] +
                mat_A[66][0] * mat_B[65][0] +
                mat_A[66][1] * mat_B[73][0] +
                mat_A[66][2] * mat_B[81][0] +
                mat_A[66][3] * mat_B[89][0] +
                mat_A[67][0] * mat_B[97][0] +
                mat_A[67][1] * mat_B[105][0] +
                mat_A[67][2] * mat_B[113][0] +
                mat_A[67][3] * mat_B[121][0] +
                mat_A[68][0] * mat_B[129][0] +
                mat_A[68][1] * mat_B[137][0] +
                mat_A[68][2] * mat_B[145][0] +
                mat_A[68][3] * mat_B[153][0] +
                mat_A[69][0] * mat_B[161][0] +
                mat_A[69][1] * mat_B[169][0] +
                mat_A[69][2] * mat_B[177][0] +
                mat_A[69][3] * mat_B[185][0] +
                mat_A[70][0] * mat_B[193][0] +
                mat_A[70][1] * mat_B[201][0] +
                mat_A[70][2] * mat_B[209][0] +
                mat_A[70][3] * mat_B[217][0] +
                mat_A[71][0] * mat_B[225][0] +
                mat_A[71][1] * mat_B[233][0] +
                mat_A[71][2] * mat_B[241][0] +
                mat_A[71][3] * mat_B[249][0];
    mat_C[65][1] <=
                mat_A[64][0] * mat_B[1][1] +
                mat_A[64][1] * mat_B[9][1] +
                mat_A[64][2] * mat_B[17][1] +
                mat_A[64][3] * mat_B[25][1] +
                mat_A[65][0] * mat_B[33][1] +
                mat_A[65][1] * mat_B[41][1] +
                mat_A[65][2] * mat_B[49][1] +
                mat_A[65][3] * mat_B[57][1] +
                mat_A[66][0] * mat_B[65][1] +
                mat_A[66][1] * mat_B[73][1] +
                mat_A[66][2] * mat_B[81][1] +
                mat_A[66][3] * mat_B[89][1] +
                mat_A[67][0] * mat_B[97][1] +
                mat_A[67][1] * mat_B[105][1] +
                mat_A[67][2] * mat_B[113][1] +
                mat_A[67][3] * mat_B[121][1] +
                mat_A[68][0] * mat_B[129][1] +
                mat_A[68][1] * mat_B[137][1] +
                mat_A[68][2] * mat_B[145][1] +
                mat_A[68][3] * mat_B[153][1] +
                mat_A[69][0] * mat_B[161][1] +
                mat_A[69][1] * mat_B[169][1] +
                mat_A[69][2] * mat_B[177][1] +
                mat_A[69][3] * mat_B[185][1] +
                mat_A[70][0] * mat_B[193][1] +
                mat_A[70][1] * mat_B[201][1] +
                mat_A[70][2] * mat_B[209][1] +
                mat_A[70][3] * mat_B[217][1] +
                mat_A[71][0] * mat_B[225][1] +
                mat_A[71][1] * mat_B[233][1] +
                mat_A[71][2] * mat_B[241][1] +
                mat_A[71][3] * mat_B[249][1];
    mat_C[65][2] <=
                mat_A[64][0] * mat_B[1][2] +
                mat_A[64][1] * mat_B[9][2] +
                mat_A[64][2] * mat_B[17][2] +
                mat_A[64][3] * mat_B[25][2] +
                mat_A[65][0] * mat_B[33][2] +
                mat_A[65][1] * mat_B[41][2] +
                mat_A[65][2] * mat_B[49][2] +
                mat_A[65][3] * mat_B[57][2] +
                mat_A[66][0] * mat_B[65][2] +
                mat_A[66][1] * mat_B[73][2] +
                mat_A[66][2] * mat_B[81][2] +
                mat_A[66][3] * mat_B[89][2] +
                mat_A[67][0] * mat_B[97][2] +
                mat_A[67][1] * mat_B[105][2] +
                mat_A[67][2] * mat_B[113][2] +
                mat_A[67][3] * mat_B[121][2] +
                mat_A[68][0] * mat_B[129][2] +
                mat_A[68][1] * mat_B[137][2] +
                mat_A[68][2] * mat_B[145][2] +
                mat_A[68][3] * mat_B[153][2] +
                mat_A[69][0] * mat_B[161][2] +
                mat_A[69][1] * mat_B[169][2] +
                mat_A[69][2] * mat_B[177][2] +
                mat_A[69][3] * mat_B[185][2] +
                mat_A[70][0] * mat_B[193][2] +
                mat_A[70][1] * mat_B[201][2] +
                mat_A[70][2] * mat_B[209][2] +
                mat_A[70][3] * mat_B[217][2] +
                mat_A[71][0] * mat_B[225][2] +
                mat_A[71][1] * mat_B[233][2] +
                mat_A[71][2] * mat_B[241][2] +
                mat_A[71][3] * mat_B[249][2];
    mat_C[65][3] <=
                mat_A[64][0] * mat_B[1][3] +
                mat_A[64][1] * mat_B[9][3] +
                mat_A[64][2] * mat_B[17][3] +
                mat_A[64][3] * mat_B[25][3] +
                mat_A[65][0] * mat_B[33][3] +
                mat_A[65][1] * mat_B[41][3] +
                mat_A[65][2] * mat_B[49][3] +
                mat_A[65][3] * mat_B[57][3] +
                mat_A[66][0] * mat_B[65][3] +
                mat_A[66][1] * mat_B[73][3] +
                mat_A[66][2] * mat_B[81][3] +
                mat_A[66][3] * mat_B[89][3] +
                mat_A[67][0] * mat_B[97][3] +
                mat_A[67][1] * mat_B[105][3] +
                mat_A[67][2] * mat_B[113][3] +
                mat_A[67][3] * mat_B[121][3] +
                mat_A[68][0] * mat_B[129][3] +
                mat_A[68][1] * mat_B[137][3] +
                mat_A[68][2] * mat_B[145][3] +
                mat_A[68][3] * mat_B[153][3] +
                mat_A[69][0] * mat_B[161][3] +
                mat_A[69][1] * mat_B[169][3] +
                mat_A[69][2] * mat_B[177][3] +
                mat_A[69][3] * mat_B[185][3] +
                mat_A[70][0] * mat_B[193][3] +
                mat_A[70][1] * mat_B[201][3] +
                mat_A[70][2] * mat_B[209][3] +
                mat_A[70][3] * mat_B[217][3] +
                mat_A[71][0] * mat_B[225][3] +
                mat_A[71][1] * mat_B[233][3] +
                mat_A[71][2] * mat_B[241][3] +
                mat_A[71][3] * mat_B[249][3];
    mat_C[66][0] <=
                mat_A[64][0] * mat_B[2][0] +
                mat_A[64][1] * mat_B[10][0] +
                mat_A[64][2] * mat_B[18][0] +
                mat_A[64][3] * mat_B[26][0] +
                mat_A[65][0] * mat_B[34][0] +
                mat_A[65][1] * mat_B[42][0] +
                mat_A[65][2] * mat_B[50][0] +
                mat_A[65][3] * mat_B[58][0] +
                mat_A[66][0] * mat_B[66][0] +
                mat_A[66][1] * mat_B[74][0] +
                mat_A[66][2] * mat_B[82][0] +
                mat_A[66][3] * mat_B[90][0] +
                mat_A[67][0] * mat_B[98][0] +
                mat_A[67][1] * mat_B[106][0] +
                mat_A[67][2] * mat_B[114][0] +
                mat_A[67][3] * mat_B[122][0] +
                mat_A[68][0] * mat_B[130][0] +
                mat_A[68][1] * mat_B[138][0] +
                mat_A[68][2] * mat_B[146][0] +
                mat_A[68][3] * mat_B[154][0] +
                mat_A[69][0] * mat_B[162][0] +
                mat_A[69][1] * mat_B[170][0] +
                mat_A[69][2] * mat_B[178][0] +
                mat_A[69][3] * mat_B[186][0] +
                mat_A[70][0] * mat_B[194][0] +
                mat_A[70][1] * mat_B[202][0] +
                mat_A[70][2] * mat_B[210][0] +
                mat_A[70][3] * mat_B[218][0] +
                mat_A[71][0] * mat_B[226][0] +
                mat_A[71][1] * mat_B[234][0] +
                mat_A[71][2] * mat_B[242][0] +
                mat_A[71][3] * mat_B[250][0];
    mat_C[66][1] <=
                mat_A[64][0] * mat_B[2][1] +
                mat_A[64][1] * mat_B[10][1] +
                mat_A[64][2] * mat_B[18][1] +
                mat_A[64][3] * mat_B[26][1] +
                mat_A[65][0] * mat_B[34][1] +
                mat_A[65][1] * mat_B[42][1] +
                mat_A[65][2] * mat_B[50][1] +
                mat_A[65][3] * mat_B[58][1] +
                mat_A[66][0] * mat_B[66][1] +
                mat_A[66][1] * mat_B[74][1] +
                mat_A[66][2] * mat_B[82][1] +
                mat_A[66][3] * mat_B[90][1] +
                mat_A[67][0] * mat_B[98][1] +
                mat_A[67][1] * mat_B[106][1] +
                mat_A[67][2] * mat_B[114][1] +
                mat_A[67][3] * mat_B[122][1] +
                mat_A[68][0] * mat_B[130][1] +
                mat_A[68][1] * mat_B[138][1] +
                mat_A[68][2] * mat_B[146][1] +
                mat_A[68][3] * mat_B[154][1] +
                mat_A[69][0] * mat_B[162][1] +
                mat_A[69][1] * mat_B[170][1] +
                mat_A[69][2] * mat_B[178][1] +
                mat_A[69][3] * mat_B[186][1] +
                mat_A[70][0] * mat_B[194][1] +
                mat_A[70][1] * mat_B[202][1] +
                mat_A[70][2] * mat_B[210][1] +
                mat_A[70][3] * mat_B[218][1] +
                mat_A[71][0] * mat_B[226][1] +
                mat_A[71][1] * mat_B[234][1] +
                mat_A[71][2] * mat_B[242][1] +
                mat_A[71][3] * mat_B[250][1];
    mat_C[66][2] <=
                mat_A[64][0] * mat_B[2][2] +
                mat_A[64][1] * mat_B[10][2] +
                mat_A[64][2] * mat_B[18][2] +
                mat_A[64][3] * mat_B[26][2] +
                mat_A[65][0] * mat_B[34][2] +
                mat_A[65][1] * mat_B[42][2] +
                mat_A[65][2] * mat_B[50][2] +
                mat_A[65][3] * mat_B[58][2] +
                mat_A[66][0] * mat_B[66][2] +
                mat_A[66][1] * mat_B[74][2] +
                mat_A[66][2] * mat_B[82][2] +
                mat_A[66][3] * mat_B[90][2] +
                mat_A[67][0] * mat_B[98][2] +
                mat_A[67][1] * mat_B[106][2] +
                mat_A[67][2] * mat_B[114][2] +
                mat_A[67][3] * mat_B[122][2] +
                mat_A[68][0] * mat_B[130][2] +
                mat_A[68][1] * mat_B[138][2] +
                mat_A[68][2] * mat_B[146][2] +
                mat_A[68][3] * mat_B[154][2] +
                mat_A[69][0] * mat_B[162][2] +
                mat_A[69][1] * mat_B[170][2] +
                mat_A[69][2] * mat_B[178][2] +
                mat_A[69][3] * mat_B[186][2] +
                mat_A[70][0] * mat_B[194][2] +
                mat_A[70][1] * mat_B[202][2] +
                mat_A[70][2] * mat_B[210][2] +
                mat_A[70][3] * mat_B[218][2] +
                mat_A[71][0] * mat_B[226][2] +
                mat_A[71][1] * mat_B[234][2] +
                mat_A[71][2] * mat_B[242][2] +
                mat_A[71][3] * mat_B[250][2];
    mat_C[66][3] <=
                mat_A[64][0] * mat_B[2][3] +
                mat_A[64][1] * mat_B[10][3] +
                mat_A[64][2] * mat_B[18][3] +
                mat_A[64][3] * mat_B[26][3] +
                mat_A[65][0] * mat_B[34][3] +
                mat_A[65][1] * mat_B[42][3] +
                mat_A[65][2] * mat_B[50][3] +
                mat_A[65][3] * mat_B[58][3] +
                mat_A[66][0] * mat_B[66][3] +
                mat_A[66][1] * mat_B[74][3] +
                mat_A[66][2] * mat_B[82][3] +
                mat_A[66][3] * mat_B[90][3] +
                mat_A[67][0] * mat_B[98][3] +
                mat_A[67][1] * mat_B[106][3] +
                mat_A[67][2] * mat_B[114][3] +
                mat_A[67][3] * mat_B[122][3] +
                mat_A[68][0] * mat_B[130][3] +
                mat_A[68][1] * mat_B[138][3] +
                mat_A[68][2] * mat_B[146][3] +
                mat_A[68][3] * mat_B[154][3] +
                mat_A[69][0] * mat_B[162][3] +
                mat_A[69][1] * mat_B[170][3] +
                mat_A[69][2] * mat_B[178][3] +
                mat_A[69][3] * mat_B[186][3] +
                mat_A[70][0] * mat_B[194][3] +
                mat_A[70][1] * mat_B[202][3] +
                mat_A[70][2] * mat_B[210][3] +
                mat_A[70][3] * mat_B[218][3] +
                mat_A[71][0] * mat_B[226][3] +
                mat_A[71][1] * mat_B[234][3] +
                mat_A[71][2] * mat_B[242][3] +
                mat_A[71][3] * mat_B[250][3];
    mat_C[67][0] <=
                mat_A[64][0] * mat_B[3][0] +
                mat_A[64][1] * mat_B[11][0] +
                mat_A[64][2] * mat_B[19][0] +
                mat_A[64][3] * mat_B[27][0] +
                mat_A[65][0] * mat_B[35][0] +
                mat_A[65][1] * mat_B[43][0] +
                mat_A[65][2] * mat_B[51][0] +
                mat_A[65][3] * mat_B[59][0] +
                mat_A[66][0] * mat_B[67][0] +
                mat_A[66][1] * mat_B[75][0] +
                mat_A[66][2] * mat_B[83][0] +
                mat_A[66][3] * mat_B[91][0] +
                mat_A[67][0] * mat_B[99][0] +
                mat_A[67][1] * mat_B[107][0] +
                mat_A[67][2] * mat_B[115][0] +
                mat_A[67][3] * mat_B[123][0] +
                mat_A[68][0] * mat_B[131][0] +
                mat_A[68][1] * mat_B[139][0] +
                mat_A[68][2] * mat_B[147][0] +
                mat_A[68][3] * mat_B[155][0] +
                mat_A[69][0] * mat_B[163][0] +
                mat_A[69][1] * mat_B[171][0] +
                mat_A[69][2] * mat_B[179][0] +
                mat_A[69][3] * mat_B[187][0] +
                mat_A[70][0] * mat_B[195][0] +
                mat_A[70][1] * mat_B[203][0] +
                mat_A[70][2] * mat_B[211][0] +
                mat_A[70][3] * mat_B[219][0] +
                mat_A[71][0] * mat_B[227][0] +
                mat_A[71][1] * mat_B[235][0] +
                mat_A[71][2] * mat_B[243][0] +
                mat_A[71][3] * mat_B[251][0];
    mat_C[67][1] <=
                mat_A[64][0] * mat_B[3][1] +
                mat_A[64][1] * mat_B[11][1] +
                mat_A[64][2] * mat_B[19][1] +
                mat_A[64][3] * mat_B[27][1] +
                mat_A[65][0] * mat_B[35][1] +
                mat_A[65][1] * mat_B[43][1] +
                mat_A[65][2] * mat_B[51][1] +
                mat_A[65][3] * mat_B[59][1] +
                mat_A[66][0] * mat_B[67][1] +
                mat_A[66][1] * mat_B[75][1] +
                mat_A[66][2] * mat_B[83][1] +
                mat_A[66][3] * mat_B[91][1] +
                mat_A[67][0] * mat_B[99][1] +
                mat_A[67][1] * mat_B[107][1] +
                mat_A[67][2] * mat_B[115][1] +
                mat_A[67][3] * mat_B[123][1] +
                mat_A[68][0] * mat_B[131][1] +
                mat_A[68][1] * mat_B[139][1] +
                mat_A[68][2] * mat_B[147][1] +
                mat_A[68][3] * mat_B[155][1] +
                mat_A[69][0] * mat_B[163][1] +
                mat_A[69][1] * mat_B[171][1] +
                mat_A[69][2] * mat_B[179][1] +
                mat_A[69][3] * mat_B[187][1] +
                mat_A[70][0] * mat_B[195][1] +
                mat_A[70][1] * mat_B[203][1] +
                mat_A[70][2] * mat_B[211][1] +
                mat_A[70][3] * mat_B[219][1] +
                mat_A[71][0] * mat_B[227][1] +
                mat_A[71][1] * mat_B[235][1] +
                mat_A[71][2] * mat_B[243][1] +
                mat_A[71][3] * mat_B[251][1];
    mat_C[67][2] <=
                mat_A[64][0] * mat_B[3][2] +
                mat_A[64][1] * mat_B[11][2] +
                mat_A[64][2] * mat_B[19][2] +
                mat_A[64][3] * mat_B[27][2] +
                mat_A[65][0] * mat_B[35][2] +
                mat_A[65][1] * mat_B[43][2] +
                mat_A[65][2] * mat_B[51][2] +
                mat_A[65][3] * mat_B[59][2] +
                mat_A[66][0] * mat_B[67][2] +
                mat_A[66][1] * mat_B[75][2] +
                mat_A[66][2] * mat_B[83][2] +
                mat_A[66][3] * mat_B[91][2] +
                mat_A[67][0] * mat_B[99][2] +
                mat_A[67][1] * mat_B[107][2] +
                mat_A[67][2] * mat_B[115][2] +
                mat_A[67][3] * mat_B[123][2] +
                mat_A[68][0] * mat_B[131][2] +
                mat_A[68][1] * mat_B[139][2] +
                mat_A[68][2] * mat_B[147][2] +
                mat_A[68][3] * mat_B[155][2] +
                mat_A[69][0] * mat_B[163][2] +
                mat_A[69][1] * mat_B[171][2] +
                mat_A[69][2] * mat_B[179][2] +
                mat_A[69][3] * mat_B[187][2] +
                mat_A[70][0] * mat_B[195][2] +
                mat_A[70][1] * mat_B[203][2] +
                mat_A[70][2] * mat_B[211][2] +
                mat_A[70][3] * mat_B[219][2] +
                mat_A[71][0] * mat_B[227][2] +
                mat_A[71][1] * mat_B[235][2] +
                mat_A[71][2] * mat_B[243][2] +
                mat_A[71][3] * mat_B[251][2];
    mat_C[67][3] <=
                mat_A[64][0] * mat_B[3][3] +
                mat_A[64][1] * mat_B[11][3] +
                mat_A[64][2] * mat_B[19][3] +
                mat_A[64][3] * mat_B[27][3] +
                mat_A[65][0] * mat_B[35][3] +
                mat_A[65][1] * mat_B[43][3] +
                mat_A[65][2] * mat_B[51][3] +
                mat_A[65][3] * mat_B[59][3] +
                mat_A[66][0] * mat_B[67][3] +
                mat_A[66][1] * mat_B[75][3] +
                mat_A[66][2] * mat_B[83][3] +
                mat_A[66][3] * mat_B[91][3] +
                mat_A[67][0] * mat_B[99][3] +
                mat_A[67][1] * mat_B[107][3] +
                mat_A[67][2] * mat_B[115][3] +
                mat_A[67][3] * mat_B[123][3] +
                mat_A[68][0] * mat_B[131][3] +
                mat_A[68][1] * mat_B[139][3] +
                mat_A[68][2] * mat_B[147][3] +
                mat_A[68][3] * mat_B[155][3] +
                mat_A[69][0] * mat_B[163][3] +
                mat_A[69][1] * mat_B[171][3] +
                mat_A[69][2] * mat_B[179][3] +
                mat_A[69][3] * mat_B[187][3] +
                mat_A[70][0] * mat_B[195][3] +
                mat_A[70][1] * mat_B[203][3] +
                mat_A[70][2] * mat_B[211][3] +
                mat_A[70][3] * mat_B[219][3] +
                mat_A[71][0] * mat_B[227][3] +
                mat_A[71][1] * mat_B[235][3] +
                mat_A[71][2] * mat_B[243][3] +
                mat_A[71][3] * mat_B[251][3];
    mat_C[68][0] <=
                mat_A[64][0] * mat_B[4][0] +
                mat_A[64][1] * mat_B[12][0] +
                mat_A[64][2] * mat_B[20][0] +
                mat_A[64][3] * mat_B[28][0] +
                mat_A[65][0] * mat_B[36][0] +
                mat_A[65][1] * mat_B[44][0] +
                mat_A[65][2] * mat_B[52][0] +
                mat_A[65][3] * mat_B[60][0] +
                mat_A[66][0] * mat_B[68][0] +
                mat_A[66][1] * mat_B[76][0] +
                mat_A[66][2] * mat_B[84][0] +
                mat_A[66][3] * mat_B[92][0] +
                mat_A[67][0] * mat_B[100][0] +
                mat_A[67][1] * mat_B[108][0] +
                mat_A[67][2] * mat_B[116][0] +
                mat_A[67][3] * mat_B[124][0] +
                mat_A[68][0] * mat_B[132][0] +
                mat_A[68][1] * mat_B[140][0] +
                mat_A[68][2] * mat_B[148][0] +
                mat_A[68][3] * mat_B[156][0] +
                mat_A[69][0] * mat_B[164][0] +
                mat_A[69][1] * mat_B[172][0] +
                mat_A[69][2] * mat_B[180][0] +
                mat_A[69][3] * mat_B[188][0] +
                mat_A[70][0] * mat_B[196][0] +
                mat_A[70][1] * mat_B[204][0] +
                mat_A[70][2] * mat_B[212][0] +
                mat_A[70][3] * mat_B[220][0] +
                mat_A[71][0] * mat_B[228][0] +
                mat_A[71][1] * mat_B[236][0] +
                mat_A[71][2] * mat_B[244][0] +
                mat_A[71][3] * mat_B[252][0];
    mat_C[68][1] <=
                mat_A[64][0] * mat_B[4][1] +
                mat_A[64][1] * mat_B[12][1] +
                mat_A[64][2] * mat_B[20][1] +
                mat_A[64][3] * mat_B[28][1] +
                mat_A[65][0] * mat_B[36][1] +
                mat_A[65][1] * mat_B[44][1] +
                mat_A[65][2] * mat_B[52][1] +
                mat_A[65][3] * mat_B[60][1] +
                mat_A[66][0] * mat_B[68][1] +
                mat_A[66][1] * mat_B[76][1] +
                mat_A[66][2] * mat_B[84][1] +
                mat_A[66][3] * mat_B[92][1] +
                mat_A[67][0] * mat_B[100][1] +
                mat_A[67][1] * mat_B[108][1] +
                mat_A[67][2] * mat_B[116][1] +
                mat_A[67][3] * mat_B[124][1] +
                mat_A[68][0] * mat_B[132][1] +
                mat_A[68][1] * mat_B[140][1] +
                mat_A[68][2] * mat_B[148][1] +
                mat_A[68][3] * mat_B[156][1] +
                mat_A[69][0] * mat_B[164][1] +
                mat_A[69][1] * mat_B[172][1] +
                mat_A[69][2] * mat_B[180][1] +
                mat_A[69][3] * mat_B[188][1] +
                mat_A[70][0] * mat_B[196][1] +
                mat_A[70][1] * mat_B[204][1] +
                mat_A[70][2] * mat_B[212][1] +
                mat_A[70][3] * mat_B[220][1] +
                mat_A[71][0] * mat_B[228][1] +
                mat_A[71][1] * mat_B[236][1] +
                mat_A[71][2] * mat_B[244][1] +
                mat_A[71][3] * mat_B[252][1];
    mat_C[68][2] <=
                mat_A[64][0] * mat_B[4][2] +
                mat_A[64][1] * mat_B[12][2] +
                mat_A[64][2] * mat_B[20][2] +
                mat_A[64][3] * mat_B[28][2] +
                mat_A[65][0] * mat_B[36][2] +
                mat_A[65][1] * mat_B[44][2] +
                mat_A[65][2] * mat_B[52][2] +
                mat_A[65][3] * mat_B[60][2] +
                mat_A[66][0] * mat_B[68][2] +
                mat_A[66][1] * mat_B[76][2] +
                mat_A[66][2] * mat_B[84][2] +
                mat_A[66][3] * mat_B[92][2] +
                mat_A[67][0] * mat_B[100][2] +
                mat_A[67][1] * mat_B[108][2] +
                mat_A[67][2] * mat_B[116][2] +
                mat_A[67][3] * mat_B[124][2] +
                mat_A[68][0] * mat_B[132][2] +
                mat_A[68][1] * mat_B[140][2] +
                mat_A[68][2] * mat_B[148][2] +
                mat_A[68][3] * mat_B[156][2] +
                mat_A[69][0] * mat_B[164][2] +
                mat_A[69][1] * mat_B[172][2] +
                mat_A[69][2] * mat_B[180][2] +
                mat_A[69][3] * mat_B[188][2] +
                mat_A[70][0] * mat_B[196][2] +
                mat_A[70][1] * mat_B[204][2] +
                mat_A[70][2] * mat_B[212][2] +
                mat_A[70][3] * mat_B[220][2] +
                mat_A[71][0] * mat_B[228][2] +
                mat_A[71][1] * mat_B[236][2] +
                mat_A[71][2] * mat_B[244][2] +
                mat_A[71][3] * mat_B[252][2];
    mat_C[68][3] <=
                mat_A[64][0] * mat_B[4][3] +
                mat_A[64][1] * mat_B[12][3] +
                mat_A[64][2] * mat_B[20][3] +
                mat_A[64][3] * mat_B[28][3] +
                mat_A[65][0] * mat_B[36][3] +
                mat_A[65][1] * mat_B[44][3] +
                mat_A[65][2] * mat_B[52][3] +
                mat_A[65][3] * mat_B[60][3] +
                mat_A[66][0] * mat_B[68][3] +
                mat_A[66][1] * mat_B[76][3] +
                mat_A[66][2] * mat_B[84][3] +
                mat_A[66][3] * mat_B[92][3] +
                mat_A[67][0] * mat_B[100][3] +
                mat_A[67][1] * mat_B[108][3] +
                mat_A[67][2] * mat_B[116][3] +
                mat_A[67][3] * mat_B[124][3] +
                mat_A[68][0] * mat_B[132][3] +
                mat_A[68][1] * mat_B[140][3] +
                mat_A[68][2] * mat_B[148][3] +
                mat_A[68][3] * mat_B[156][3] +
                mat_A[69][0] * mat_B[164][3] +
                mat_A[69][1] * mat_B[172][3] +
                mat_A[69][2] * mat_B[180][3] +
                mat_A[69][3] * mat_B[188][3] +
                mat_A[70][0] * mat_B[196][3] +
                mat_A[70][1] * mat_B[204][3] +
                mat_A[70][2] * mat_B[212][3] +
                mat_A[70][3] * mat_B[220][3] +
                mat_A[71][0] * mat_B[228][3] +
                mat_A[71][1] * mat_B[236][3] +
                mat_A[71][2] * mat_B[244][3] +
                mat_A[71][3] * mat_B[252][3];
    mat_C[69][0] <=
                mat_A[64][0] * mat_B[5][0] +
                mat_A[64][1] * mat_B[13][0] +
                mat_A[64][2] * mat_B[21][0] +
                mat_A[64][3] * mat_B[29][0] +
                mat_A[65][0] * mat_B[37][0] +
                mat_A[65][1] * mat_B[45][0] +
                mat_A[65][2] * mat_B[53][0] +
                mat_A[65][3] * mat_B[61][0] +
                mat_A[66][0] * mat_B[69][0] +
                mat_A[66][1] * mat_B[77][0] +
                mat_A[66][2] * mat_B[85][0] +
                mat_A[66][3] * mat_B[93][0] +
                mat_A[67][0] * mat_B[101][0] +
                mat_A[67][1] * mat_B[109][0] +
                mat_A[67][2] * mat_B[117][0] +
                mat_A[67][3] * mat_B[125][0] +
                mat_A[68][0] * mat_B[133][0] +
                mat_A[68][1] * mat_B[141][0] +
                mat_A[68][2] * mat_B[149][0] +
                mat_A[68][3] * mat_B[157][0] +
                mat_A[69][0] * mat_B[165][0] +
                mat_A[69][1] * mat_B[173][0] +
                mat_A[69][2] * mat_B[181][0] +
                mat_A[69][3] * mat_B[189][0] +
                mat_A[70][0] * mat_B[197][0] +
                mat_A[70][1] * mat_B[205][0] +
                mat_A[70][2] * mat_B[213][0] +
                mat_A[70][3] * mat_B[221][0] +
                mat_A[71][0] * mat_B[229][0] +
                mat_A[71][1] * mat_B[237][0] +
                mat_A[71][2] * mat_B[245][0] +
                mat_A[71][3] * mat_B[253][0];
    mat_C[69][1] <=
                mat_A[64][0] * mat_B[5][1] +
                mat_A[64][1] * mat_B[13][1] +
                mat_A[64][2] * mat_B[21][1] +
                mat_A[64][3] * mat_B[29][1] +
                mat_A[65][0] * mat_B[37][1] +
                mat_A[65][1] * mat_B[45][1] +
                mat_A[65][2] * mat_B[53][1] +
                mat_A[65][3] * mat_B[61][1] +
                mat_A[66][0] * mat_B[69][1] +
                mat_A[66][1] * mat_B[77][1] +
                mat_A[66][2] * mat_B[85][1] +
                mat_A[66][3] * mat_B[93][1] +
                mat_A[67][0] * mat_B[101][1] +
                mat_A[67][1] * mat_B[109][1] +
                mat_A[67][2] * mat_B[117][1] +
                mat_A[67][3] * mat_B[125][1] +
                mat_A[68][0] * mat_B[133][1] +
                mat_A[68][1] * mat_B[141][1] +
                mat_A[68][2] * mat_B[149][1] +
                mat_A[68][3] * mat_B[157][1] +
                mat_A[69][0] * mat_B[165][1] +
                mat_A[69][1] * mat_B[173][1] +
                mat_A[69][2] * mat_B[181][1] +
                mat_A[69][3] * mat_B[189][1] +
                mat_A[70][0] * mat_B[197][1] +
                mat_A[70][1] * mat_B[205][1] +
                mat_A[70][2] * mat_B[213][1] +
                mat_A[70][3] * mat_B[221][1] +
                mat_A[71][0] * mat_B[229][1] +
                mat_A[71][1] * mat_B[237][1] +
                mat_A[71][2] * mat_B[245][1] +
                mat_A[71][3] * mat_B[253][1];
    mat_C[69][2] <=
                mat_A[64][0] * mat_B[5][2] +
                mat_A[64][1] * mat_B[13][2] +
                mat_A[64][2] * mat_B[21][2] +
                mat_A[64][3] * mat_B[29][2] +
                mat_A[65][0] * mat_B[37][2] +
                mat_A[65][1] * mat_B[45][2] +
                mat_A[65][2] * mat_B[53][2] +
                mat_A[65][3] * mat_B[61][2] +
                mat_A[66][0] * mat_B[69][2] +
                mat_A[66][1] * mat_B[77][2] +
                mat_A[66][2] * mat_B[85][2] +
                mat_A[66][3] * mat_B[93][2] +
                mat_A[67][0] * mat_B[101][2] +
                mat_A[67][1] * mat_B[109][2] +
                mat_A[67][2] * mat_B[117][2] +
                mat_A[67][3] * mat_B[125][2] +
                mat_A[68][0] * mat_B[133][2] +
                mat_A[68][1] * mat_B[141][2] +
                mat_A[68][2] * mat_B[149][2] +
                mat_A[68][3] * mat_B[157][2] +
                mat_A[69][0] * mat_B[165][2] +
                mat_A[69][1] * mat_B[173][2] +
                mat_A[69][2] * mat_B[181][2] +
                mat_A[69][3] * mat_B[189][2] +
                mat_A[70][0] * mat_B[197][2] +
                mat_A[70][1] * mat_B[205][2] +
                mat_A[70][2] * mat_B[213][2] +
                mat_A[70][3] * mat_B[221][2] +
                mat_A[71][0] * mat_B[229][2] +
                mat_A[71][1] * mat_B[237][2] +
                mat_A[71][2] * mat_B[245][2] +
                mat_A[71][3] * mat_B[253][2];
    mat_C[69][3] <=
                mat_A[64][0] * mat_B[5][3] +
                mat_A[64][1] * mat_B[13][3] +
                mat_A[64][2] * mat_B[21][3] +
                mat_A[64][3] * mat_B[29][3] +
                mat_A[65][0] * mat_B[37][3] +
                mat_A[65][1] * mat_B[45][3] +
                mat_A[65][2] * mat_B[53][3] +
                mat_A[65][3] * mat_B[61][3] +
                mat_A[66][0] * mat_B[69][3] +
                mat_A[66][1] * mat_B[77][3] +
                mat_A[66][2] * mat_B[85][3] +
                mat_A[66][3] * mat_B[93][3] +
                mat_A[67][0] * mat_B[101][3] +
                mat_A[67][1] * mat_B[109][3] +
                mat_A[67][2] * mat_B[117][3] +
                mat_A[67][3] * mat_B[125][3] +
                mat_A[68][0] * mat_B[133][3] +
                mat_A[68][1] * mat_B[141][3] +
                mat_A[68][2] * mat_B[149][3] +
                mat_A[68][3] * mat_B[157][3] +
                mat_A[69][0] * mat_B[165][3] +
                mat_A[69][1] * mat_B[173][3] +
                mat_A[69][2] * mat_B[181][3] +
                mat_A[69][3] * mat_B[189][3] +
                mat_A[70][0] * mat_B[197][3] +
                mat_A[70][1] * mat_B[205][3] +
                mat_A[70][2] * mat_B[213][3] +
                mat_A[70][3] * mat_B[221][3] +
                mat_A[71][0] * mat_B[229][3] +
                mat_A[71][1] * mat_B[237][3] +
                mat_A[71][2] * mat_B[245][3] +
                mat_A[71][3] * mat_B[253][3];
    mat_C[70][0] <=
                mat_A[64][0] * mat_B[6][0] +
                mat_A[64][1] * mat_B[14][0] +
                mat_A[64][2] * mat_B[22][0] +
                mat_A[64][3] * mat_B[30][0] +
                mat_A[65][0] * mat_B[38][0] +
                mat_A[65][1] * mat_B[46][0] +
                mat_A[65][2] * mat_B[54][0] +
                mat_A[65][3] * mat_B[62][0] +
                mat_A[66][0] * mat_B[70][0] +
                mat_A[66][1] * mat_B[78][0] +
                mat_A[66][2] * mat_B[86][0] +
                mat_A[66][3] * mat_B[94][0] +
                mat_A[67][0] * mat_B[102][0] +
                mat_A[67][1] * mat_B[110][0] +
                mat_A[67][2] * mat_B[118][0] +
                mat_A[67][3] * mat_B[126][0] +
                mat_A[68][0] * mat_B[134][0] +
                mat_A[68][1] * mat_B[142][0] +
                mat_A[68][2] * mat_B[150][0] +
                mat_A[68][3] * mat_B[158][0] +
                mat_A[69][0] * mat_B[166][0] +
                mat_A[69][1] * mat_B[174][0] +
                mat_A[69][2] * mat_B[182][0] +
                mat_A[69][3] * mat_B[190][0] +
                mat_A[70][0] * mat_B[198][0] +
                mat_A[70][1] * mat_B[206][0] +
                mat_A[70][2] * mat_B[214][0] +
                mat_A[70][3] * mat_B[222][0] +
                mat_A[71][0] * mat_B[230][0] +
                mat_A[71][1] * mat_B[238][0] +
                mat_A[71][2] * mat_B[246][0] +
                mat_A[71][3] * mat_B[254][0];
    mat_C[70][1] <=
                mat_A[64][0] * mat_B[6][1] +
                mat_A[64][1] * mat_B[14][1] +
                mat_A[64][2] * mat_B[22][1] +
                mat_A[64][3] * mat_B[30][1] +
                mat_A[65][0] * mat_B[38][1] +
                mat_A[65][1] * mat_B[46][1] +
                mat_A[65][2] * mat_B[54][1] +
                mat_A[65][3] * mat_B[62][1] +
                mat_A[66][0] * mat_B[70][1] +
                mat_A[66][1] * mat_B[78][1] +
                mat_A[66][2] * mat_B[86][1] +
                mat_A[66][3] * mat_B[94][1] +
                mat_A[67][0] * mat_B[102][1] +
                mat_A[67][1] * mat_B[110][1] +
                mat_A[67][2] * mat_B[118][1] +
                mat_A[67][3] * mat_B[126][1] +
                mat_A[68][0] * mat_B[134][1] +
                mat_A[68][1] * mat_B[142][1] +
                mat_A[68][2] * mat_B[150][1] +
                mat_A[68][3] * mat_B[158][1] +
                mat_A[69][0] * mat_B[166][1] +
                mat_A[69][1] * mat_B[174][1] +
                mat_A[69][2] * mat_B[182][1] +
                mat_A[69][3] * mat_B[190][1] +
                mat_A[70][0] * mat_B[198][1] +
                mat_A[70][1] * mat_B[206][1] +
                mat_A[70][2] * mat_B[214][1] +
                mat_A[70][3] * mat_B[222][1] +
                mat_A[71][0] * mat_B[230][1] +
                mat_A[71][1] * mat_B[238][1] +
                mat_A[71][2] * mat_B[246][1] +
                mat_A[71][3] * mat_B[254][1];
    mat_C[70][2] <=
                mat_A[64][0] * mat_B[6][2] +
                mat_A[64][1] * mat_B[14][2] +
                mat_A[64][2] * mat_B[22][2] +
                mat_A[64][3] * mat_B[30][2] +
                mat_A[65][0] * mat_B[38][2] +
                mat_A[65][1] * mat_B[46][2] +
                mat_A[65][2] * mat_B[54][2] +
                mat_A[65][3] * mat_B[62][2] +
                mat_A[66][0] * mat_B[70][2] +
                mat_A[66][1] * mat_B[78][2] +
                mat_A[66][2] * mat_B[86][2] +
                mat_A[66][3] * mat_B[94][2] +
                mat_A[67][0] * mat_B[102][2] +
                mat_A[67][1] * mat_B[110][2] +
                mat_A[67][2] * mat_B[118][2] +
                mat_A[67][3] * mat_B[126][2] +
                mat_A[68][0] * mat_B[134][2] +
                mat_A[68][1] * mat_B[142][2] +
                mat_A[68][2] * mat_B[150][2] +
                mat_A[68][3] * mat_B[158][2] +
                mat_A[69][0] * mat_B[166][2] +
                mat_A[69][1] * mat_B[174][2] +
                mat_A[69][2] * mat_B[182][2] +
                mat_A[69][3] * mat_B[190][2] +
                mat_A[70][0] * mat_B[198][2] +
                mat_A[70][1] * mat_B[206][2] +
                mat_A[70][2] * mat_B[214][2] +
                mat_A[70][3] * mat_B[222][2] +
                mat_A[71][0] * mat_B[230][2] +
                mat_A[71][1] * mat_B[238][2] +
                mat_A[71][2] * mat_B[246][2] +
                mat_A[71][3] * mat_B[254][2];
    mat_C[70][3] <=
                mat_A[64][0] * mat_B[6][3] +
                mat_A[64][1] * mat_B[14][3] +
                mat_A[64][2] * mat_B[22][3] +
                mat_A[64][3] * mat_B[30][3] +
                mat_A[65][0] * mat_B[38][3] +
                mat_A[65][1] * mat_B[46][3] +
                mat_A[65][2] * mat_B[54][3] +
                mat_A[65][3] * mat_B[62][3] +
                mat_A[66][0] * mat_B[70][3] +
                mat_A[66][1] * mat_B[78][3] +
                mat_A[66][2] * mat_B[86][3] +
                mat_A[66][3] * mat_B[94][3] +
                mat_A[67][0] * mat_B[102][3] +
                mat_A[67][1] * mat_B[110][3] +
                mat_A[67][2] * mat_B[118][3] +
                mat_A[67][3] * mat_B[126][3] +
                mat_A[68][0] * mat_B[134][3] +
                mat_A[68][1] * mat_B[142][3] +
                mat_A[68][2] * mat_B[150][3] +
                mat_A[68][3] * mat_B[158][3] +
                mat_A[69][0] * mat_B[166][3] +
                mat_A[69][1] * mat_B[174][3] +
                mat_A[69][2] * mat_B[182][3] +
                mat_A[69][3] * mat_B[190][3] +
                mat_A[70][0] * mat_B[198][3] +
                mat_A[70][1] * mat_B[206][3] +
                mat_A[70][2] * mat_B[214][3] +
                mat_A[70][3] * mat_B[222][3] +
                mat_A[71][0] * mat_B[230][3] +
                mat_A[71][1] * mat_B[238][3] +
                mat_A[71][2] * mat_B[246][3] +
                mat_A[71][3] * mat_B[254][3];
    mat_C[71][0] <=
                mat_A[64][0] * mat_B[7][0] +
                mat_A[64][1] * mat_B[15][0] +
                mat_A[64][2] * mat_B[23][0] +
                mat_A[64][3] * mat_B[31][0] +
                mat_A[65][0] * mat_B[39][0] +
                mat_A[65][1] * mat_B[47][0] +
                mat_A[65][2] * mat_B[55][0] +
                mat_A[65][3] * mat_B[63][0] +
                mat_A[66][0] * mat_B[71][0] +
                mat_A[66][1] * mat_B[79][0] +
                mat_A[66][2] * mat_B[87][0] +
                mat_A[66][3] * mat_B[95][0] +
                mat_A[67][0] * mat_B[103][0] +
                mat_A[67][1] * mat_B[111][0] +
                mat_A[67][2] * mat_B[119][0] +
                mat_A[67][3] * mat_B[127][0] +
                mat_A[68][0] * mat_B[135][0] +
                mat_A[68][1] * mat_B[143][0] +
                mat_A[68][2] * mat_B[151][0] +
                mat_A[68][3] * mat_B[159][0] +
                mat_A[69][0] * mat_B[167][0] +
                mat_A[69][1] * mat_B[175][0] +
                mat_A[69][2] * mat_B[183][0] +
                mat_A[69][3] * mat_B[191][0] +
                mat_A[70][0] * mat_B[199][0] +
                mat_A[70][1] * mat_B[207][0] +
                mat_A[70][2] * mat_B[215][0] +
                mat_A[70][3] * mat_B[223][0] +
                mat_A[71][0] * mat_B[231][0] +
                mat_A[71][1] * mat_B[239][0] +
                mat_A[71][2] * mat_B[247][0] +
                mat_A[71][3] * mat_B[255][0];
    mat_C[71][1] <=
                mat_A[64][0] * mat_B[7][1] +
                mat_A[64][1] * mat_B[15][1] +
                mat_A[64][2] * mat_B[23][1] +
                mat_A[64][3] * mat_B[31][1] +
                mat_A[65][0] * mat_B[39][1] +
                mat_A[65][1] * mat_B[47][1] +
                mat_A[65][2] * mat_B[55][1] +
                mat_A[65][3] * mat_B[63][1] +
                mat_A[66][0] * mat_B[71][1] +
                mat_A[66][1] * mat_B[79][1] +
                mat_A[66][2] * mat_B[87][1] +
                mat_A[66][3] * mat_B[95][1] +
                mat_A[67][0] * mat_B[103][1] +
                mat_A[67][1] * mat_B[111][1] +
                mat_A[67][2] * mat_B[119][1] +
                mat_A[67][3] * mat_B[127][1] +
                mat_A[68][0] * mat_B[135][1] +
                mat_A[68][1] * mat_B[143][1] +
                mat_A[68][2] * mat_B[151][1] +
                mat_A[68][3] * mat_B[159][1] +
                mat_A[69][0] * mat_B[167][1] +
                mat_A[69][1] * mat_B[175][1] +
                mat_A[69][2] * mat_B[183][1] +
                mat_A[69][3] * mat_B[191][1] +
                mat_A[70][0] * mat_B[199][1] +
                mat_A[70][1] * mat_B[207][1] +
                mat_A[70][2] * mat_B[215][1] +
                mat_A[70][3] * mat_B[223][1] +
                mat_A[71][0] * mat_B[231][1] +
                mat_A[71][1] * mat_B[239][1] +
                mat_A[71][2] * mat_B[247][1] +
                mat_A[71][3] * mat_B[255][1];
    mat_C[71][2] <=
                mat_A[64][0] * mat_B[7][2] +
                mat_A[64][1] * mat_B[15][2] +
                mat_A[64][2] * mat_B[23][2] +
                mat_A[64][3] * mat_B[31][2] +
                mat_A[65][0] * mat_B[39][2] +
                mat_A[65][1] * mat_B[47][2] +
                mat_A[65][2] * mat_B[55][2] +
                mat_A[65][3] * mat_B[63][2] +
                mat_A[66][0] * mat_B[71][2] +
                mat_A[66][1] * mat_B[79][2] +
                mat_A[66][2] * mat_B[87][2] +
                mat_A[66][3] * mat_B[95][2] +
                mat_A[67][0] * mat_B[103][2] +
                mat_A[67][1] * mat_B[111][2] +
                mat_A[67][2] * mat_B[119][2] +
                mat_A[67][3] * mat_B[127][2] +
                mat_A[68][0] * mat_B[135][2] +
                mat_A[68][1] * mat_B[143][2] +
                mat_A[68][2] * mat_B[151][2] +
                mat_A[68][3] * mat_B[159][2] +
                mat_A[69][0] * mat_B[167][2] +
                mat_A[69][1] * mat_B[175][2] +
                mat_A[69][2] * mat_B[183][2] +
                mat_A[69][3] * mat_B[191][2] +
                mat_A[70][0] * mat_B[199][2] +
                mat_A[70][1] * mat_B[207][2] +
                mat_A[70][2] * mat_B[215][2] +
                mat_A[70][3] * mat_B[223][2] +
                mat_A[71][0] * mat_B[231][2] +
                mat_A[71][1] * mat_B[239][2] +
                mat_A[71][2] * mat_B[247][2] +
                mat_A[71][3] * mat_B[255][2];
    mat_C[71][3] <=
                mat_A[64][0] * mat_B[7][3] +
                mat_A[64][1] * mat_B[15][3] +
                mat_A[64][2] * mat_B[23][3] +
                mat_A[64][3] * mat_B[31][3] +
                mat_A[65][0] * mat_B[39][3] +
                mat_A[65][1] * mat_B[47][3] +
                mat_A[65][2] * mat_B[55][3] +
                mat_A[65][3] * mat_B[63][3] +
                mat_A[66][0] * mat_B[71][3] +
                mat_A[66][1] * mat_B[79][3] +
                mat_A[66][2] * mat_B[87][3] +
                mat_A[66][3] * mat_B[95][3] +
                mat_A[67][0] * mat_B[103][3] +
                mat_A[67][1] * mat_B[111][3] +
                mat_A[67][2] * mat_B[119][3] +
                mat_A[67][3] * mat_B[127][3] +
                mat_A[68][0] * mat_B[135][3] +
                mat_A[68][1] * mat_B[143][3] +
                mat_A[68][2] * mat_B[151][3] +
                mat_A[68][3] * mat_B[159][3] +
                mat_A[69][0] * mat_B[167][3] +
                mat_A[69][1] * mat_B[175][3] +
                mat_A[69][2] * mat_B[183][3] +
                mat_A[69][3] * mat_B[191][3] +
                mat_A[70][0] * mat_B[199][3] +
                mat_A[70][1] * mat_B[207][3] +
                mat_A[70][2] * mat_B[215][3] +
                mat_A[70][3] * mat_B[223][3] +
                mat_A[71][0] * mat_B[231][3] +
                mat_A[71][1] * mat_B[239][3] +
                mat_A[71][2] * mat_B[247][3] +
                mat_A[71][3] * mat_B[255][3];
    mat_C[72][0] <=
                mat_A[72][0] * mat_B[0][0] +
                mat_A[72][1] * mat_B[8][0] +
                mat_A[72][2] * mat_B[16][0] +
                mat_A[72][3] * mat_B[24][0] +
                mat_A[73][0] * mat_B[32][0] +
                mat_A[73][1] * mat_B[40][0] +
                mat_A[73][2] * mat_B[48][0] +
                mat_A[73][3] * mat_B[56][0] +
                mat_A[74][0] * mat_B[64][0] +
                mat_A[74][1] * mat_B[72][0] +
                mat_A[74][2] * mat_B[80][0] +
                mat_A[74][3] * mat_B[88][0] +
                mat_A[75][0] * mat_B[96][0] +
                mat_A[75][1] * mat_B[104][0] +
                mat_A[75][2] * mat_B[112][0] +
                mat_A[75][3] * mat_B[120][0] +
                mat_A[76][0] * mat_B[128][0] +
                mat_A[76][1] * mat_B[136][0] +
                mat_A[76][2] * mat_B[144][0] +
                mat_A[76][3] * mat_B[152][0] +
                mat_A[77][0] * mat_B[160][0] +
                mat_A[77][1] * mat_B[168][0] +
                mat_A[77][2] * mat_B[176][0] +
                mat_A[77][3] * mat_B[184][0] +
                mat_A[78][0] * mat_B[192][0] +
                mat_A[78][1] * mat_B[200][0] +
                mat_A[78][2] * mat_B[208][0] +
                mat_A[78][3] * mat_B[216][0] +
                mat_A[79][0] * mat_B[224][0] +
                mat_A[79][1] * mat_B[232][0] +
                mat_A[79][2] * mat_B[240][0] +
                mat_A[79][3] * mat_B[248][0];
    mat_C[72][1] <=
                mat_A[72][0] * mat_B[0][1] +
                mat_A[72][1] * mat_B[8][1] +
                mat_A[72][2] * mat_B[16][1] +
                mat_A[72][3] * mat_B[24][1] +
                mat_A[73][0] * mat_B[32][1] +
                mat_A[73][1] * mat_B[40][1] +
                mat_A[73][2] * mat_B[48][1] +
                mat_A[73][3] * mat_B[56][1] +
                mat_A[74][0] * mat_B[64][1] +
                mat_A[74][1] * mat_B[72][1] +
                mat_A[74][2] * mat_B[80][1] +
                mat_A[74][3] * mat_B[88][1] +
                mat_A[75][0] * mat_B[96][1] +
                mat_A[75][1] * mat_B[104][1] +
                mat_A[75][2] * mat_B[112][1] +
                mat_A[75][3] * mat_B[120][1] +
                mat_A[76][0] * mat_B[128][1] +
                mat_A[76][1] * mat_B[136][1] +
                mat_A[76][2] * mat_B[144][1] +
                mat_A[76][3] * mat_B[152][1] +
                mat_A[77][0] * mat_B[160][1] +
                mat_A[77][1] * mat_B[168][1] +
                mat_A[77][2] * mat_B[176][1] +
                mat_A[77][3] * mat_B[184][1] +
                mat_A[78][0] * mat_B[192][1] +
                mat_A[78][1] * mat_B[200][1] +
                mat_A[78][2] * mat_B[208][1] +
                mat_A[78][3] * mat_B[216][1] +
                mat_A[79][0] * mat_B[224][1] +
                mat_A[79][1] * mat_B[232][1] +
                mat_A[79][2] * mat_B[240][1] +
                mat_A[79][3] * mat_B[248][1];
    mat_C[72][2] <=
                mat_A[72][0] * mat_B[0][2] +
                mat_A[72][1] * mat_B[8][2] +
                mat_A[72][2] * mat_B[16][2] +
                mat_A[72][3] * mat_B[24][2] +
                mat_A[73][0] * mat_B[32][2] +
                mat_A[73][1] * mat_B[40][2] +
                mat_A[73][2] * mat_B[48][2] +
                mat_A[73][3] * mat_B[56][2] +
                mat_A[74][0] * mat_B[64][2] +
                mat_A[74][1] * mat_B[72][2] +
                mat_A[74][2] * mat_B[80][2] +
                mat_A[74][3] * mat_B[88][2] +
                mat_A[75][0] * mat_B[96][2] +
                mat_A[75][1] * mat_B[104][2] +
                mat_A[75][2] * mat_B[112][2] +
                mat_A[75][3] * mat_B[120][2] +
                mat_A[76][0] * mat_B[128][2] +
                mat_A[76][1] * mat_B[136][2] +
                mat_A[76][2] * mat_B[144][2] +
                mat_A[76][3] * mat_B[152][2] +
                mat_A[77][0] * mat_B[160][2] +
                mat_A[77][1] * mat_B[168][2] +
                mat_A[77][2] * mat_B[176][2] +
                mat_A[77][3] * mat_B[184][2] +
                mat_A[78][0] * mat_B[192][2] +
                mat_A[78][1] * mat_B[200][2] +
                mat_A[78][2] * mat_B[208][2] +
                mat_A[78][3] * mat_B[216][2] +
                mat_A[79][0] * mat_B[224][2] +
                mat_A[79][1] * mat_B[232][2] +
                mat_A[79][2] * mat_B[240][2] +
                mat_A[79][3] * mat_B[248][2];
    mat_C[72][3] <=
                mat_A[72][0] * mat_B[0][3] +
                mat_A[72][1] * mat_B[8][3] +
                mat_A[72][2] * mat_B[16][3] +
                mat_A[72][3] * mat_B[24][3] +
                mat_A[73][0] * mat_B[32][3] +
                mat_A[73][1] * mat_B[40][3] +
                mat_A[73][2] * mat_B[48][3] +
                mat_A[73][3] * mat_B[56][3] +
                mat_A[74][0] * mat_B[64][3] +
                mat_A[74][1] * mat_B[72][3] +
                mat_A[74][2] * mat_B[80][3] +
                mat_A[74][3] * mat_B[88][3] +
                mat_A[75][0] * mat_B[96][3] +
                mat_A[75][1] * mat_B[104][3] +
                mat_A[75][2] * mat_B[112][3] +
                mat_A[75][3] * mat_B[120][3] +
                mat_A[76][0] * mat_B[128][3] +
                mat_A[76][1] * mat_B[136][3] +
                mat_A[76][2] * mat_B[144][3] +
                mat_A[76][3] * mat_B[152][3] +
                mat_A[77][0] * mat_B[160][3] +
                mat_A[77][1] * mat_B[168][3] +
                mat_A[77][2] * mat_B[176][3] +
                mat_A[77][3] * mat_B[184][3] +
                mat_A[78][0] * mat_B[192][3] +
                mat_A[78][1] * mat_B[200][3] +
                mat_A[78][2] * mat_B[208][3] +
                mat_A[78][3] * mat_B[216][3] +
                mat_A[79][0] * mat_B[224][3] +
                mat_A[79][1] * mat_B[232][3] +
                mat_A[79][2] * mat_B[240][3] +
                mat_A[79][3] * mat_B[248][3];
    mat_C[73][0] <=
                mat_A[72][0] * mat_B[1][0] +
                mat_A[72][1] * mat_B[9][0] +
                mat_A[72][2] * mat_B[17][0] +
                mat_A[72][3] * mat_B[25][0] +
                mat_A[73][0] * mat_B[33][0] +
                mat_A[73][1] * mat_B[41][0] +
                mat_A[73][2] * mat_B[49][0] +
                mat_A[73][3] * mat_B[57][0] +
                mat_A[74][0] * mat_B[65][0] +
                mat_A[74][1] * mat_B[73][0] +
                mat_A[74][2] * mat_B[81][0] +
                mat_A[74][3] * mat_B[89][0] +
                mat_A[75][0] * mat_B[97][0] +
                mat_A[75][1] * mat_B[105][0] +
                mat_A[75][2] * mat_B[113][0] +
                mat_A[75][3] * mat_B[121][0] +
                mat_A[76][0] * mat_B[129][0] +
                mat_A[76][1] * mat_B[137][0] +
                mat_A[76][2] * mat_B[145][0] +
                mat_A[76][3] * mat_B[153][0] +
                mat_A[77][0] * mat_B[161][0] +
                mat_A[77][1] * mat_B[169][0] +
                mat_A[77][2] * mat_B[177][0] +
                mat_A[77][3] * mat_B[185][0] +
                mat_A[78][0] * mat_B[193][0] +
                mat_A[78][1] * mat_B[201][0] +
                mat_A[78][2] * mat_B[209][0] +
                mat_A[78][3] * mat_B[217][0] +
                mat_A[79][0] * mat_B[225][0] +
                mat_A[79][1] * mat_B[233][0] +
                mat_A[79][2] * mat_B[241][0] +
                mat_A[79][3] * mat_B[249][0];
    mat_C[73][1] <=
                mat_A[72][0] * mat_B[1][1] +
                mat_A[72][1] * mat_B[9][1] +
                mat_A[72][2] * mat_B[17][1] +
                mat_A[72][3] * mat_B[25][1] +
                mat_A[73][0] * mat_B[33][1] +
                mat_A[73][1] * mat_B[41][1] +
                mat_A[73][2] * mat_B[49][1] +
                mat_A[73][3] * mat_B[57][1] +
                mat_A[74][0] * mat_B[65][1] +
                mat_A[74][1] * mat_B[73][1] +
                mat_A[74][2] * mat_B[81][1] +
                mat_A[74][3] * mat_B[89][1] +
                mat_A[75][0] * mat_B[97][1] +
                mat_A[75][1] * mat_B[105][1] +
                mat_A[75][2] * mat_B[113][1] +
                mat_A[75][3] * mat_B[121][1] +
                mat_A[76][0] * mat_B[129][1] +
                mat_A[76][1] * mat_B[137][1] +
                mat_A[76][2] * mat_B[145][1] +
                mat_A[76][3] * mat_B[153][1] +
                mat_A[77][0] * mat_B[161][1] +
                mat_A[77][1] * mat_B[169][1] +
                mat_A[77][2] * mat_B[177][1] +
                mat_A[77][3] * mat_B[185][1] +
                mat_A[78][0] * mat_B[193][1] +
                mat_A[78][1] * mat_B[201][1] +
                mat_A[78][2] * mat_B[209][1] +
                mat_A[78][3] * mat_B[217][1] +
                mat_A[79][0] * mat_B[225][1] +
                mat_A[79][1] * mat_B[233][1] +
                mat_A[79][2] * mat_B[241][1] +
                mat_A[79][3] * mat_B[249][1];
    mat_C[73][2] <=
                mat_A[72][0] * mat_B[1][2] +
                mat_A[72][1] * mat_B[9][2] +
                mat_A[72][2] * mat_B[17][2] +
                mat_A[72][3] * mat_B[25][2] +
                mat_A[73][0] * mat_B[33][2] +
                mat_A[73][1] * mat_B[41][2] +
                mat_A[73][2] * mat_B[49][2] +
                mat_A[73][3] * mat_B[57][2] +
                mat_A[74][0] * mat_B[65][2] +
                mat_A[74][1] * mat_B[73][2] +
                mat_A[74][2] * mat_B[81][2] +
                mat_A[74][3] * mat_B[89][2] +
                mat_A[75][0] * mat_B[97][2] +
                mat_A[75][1] * mat_B[105][2] +
                mat_A[75][2] * mat_B[113][2] +
                mat_A[75][3] * mat_B[121][2] +
                mat_A[76][0] * mat_B[129][2] +
                mat_A[76][1] * mat_B[137][2] +
                mat_A[76][2] * mat_B[145][2] +
                mat_A[76][3] * mat_B[153][2] +
                mat_A[77][0] * mat_B[161][2] +
                mat_A[77][1] * mat_B[169][2] +
                mat_A[77][2] * mat_B[177][2] +
                mat_A[77][3] * mat_B[185][2] +
                mat_A[78][0] * mat_B[193][2] +
                mat_A[78][1] * mat_B[201][2] +
                mat_A[78][2] * mat_B[209][2] +
                mat_A[78][3] * mat_B[217][2] +
                mat_A[79][0] * mat_B[225][2] +
                mat_A[79][1] * mat_B[233][2] +
                mat_A[79][2] * mat_B[241][2] +
                mat_A[79][3] * mat_B[249][2];
    mat_C[73][3] <=
                mat_A[72][0] * mat_B[1][3] +
                mat_A[72][1] * mat_B[9][3] +
                mat_A[72][2] * mat_B[17][3] +
                mat_A[72][3] * mat_B[25][3] +
                mat_A[73][0] * mat_B[33][3] +
                mat_A[73][1] * mat_B[41][3] +
                mat_A[73][2] * mat_B[49][3] +
                mat_A[73][3] * mat_B[57][3] +
                mat_A[74][0] * mat_B[65][3] +
                mat_A[74][1] * mat_B[73][3] +
                mat_A[74][2] * mat_B[81][3] +
                mat_A[74][3] * mat_B[89][3] +
                mat_A[75][0] * mat_B[97][3] +
                mat_A[75][1] * mat_B[105][3] +
                mat_A[75][2] * mat_B[113][3] +
                mat_A[75][3] * mat_B[121][3] +
                mat_A[76][0] * mat_B[129][3] +
                mat_A[76][1] * mat_B[137][3] +
                mat_A[76][2] * mat_B[145][3] +
                mat_A[76][3] * mat_B[153][3] +
                mat_A[77][0] * mat_B[161][3] +
                mat_A[77][1] * mat_B[169][3] +
                mat_A[77][2] * mat_B[177][3] +
                mat_A[77][3] * mat_B[185][3] +
                mat_A[78][0] * mat_B[193][3] +
                mat_A[78][1] * mat_B[201][3] +
                mat_A[78][2] * mat_B[209][3] +
                mat_A[78][3] * mat_B[217][3] +
                mat_A[79][0] * mat_B[225][3] +
                mat_A[79][1] * mat_B[233][3] +
                mat_A[79][2] * mat_B[241][3] +
                mat_A[79][3] * mat_B[249][3];
    mat_C[74][0] <=
                mat_A[72][0] * mat_B[2][0] +
                mat_A[72][1] * mat_B[10][0] +
                mat_A[72][2] * mat_B[18][0] +
                mat_A[72][3] * mat_B[26][0] +
                mat_A[73][0] * mat_B[34][0] +
                mat_A[73][1] * mat_B[42][0] +
                mat_A[73][2] * mat_B[50][0] +
                mat_A[73][3] * mat_B[58][0] +
                mat_A[74][0] * mat_B[66][0] +
                mat_A[74][1] * mat_B[74][0] +
                mat_A[74][2] * mat_B[82][0] +
                mat_A[74][3] * mat_B[90][0] +
                mat_A[75][0] * mat_B[98][0] +
                mat_A[75][1] * mat_B[106][0] +
                mat_A[75][2] * mat_B[114][0] +
                mat_A[75][3] * mat_B[122][0] +
                mat_A[76][0] * mat_B[130][0] +
                mat_A[76][1] * mat_B[138][0] +
                mat_A[76][2] * mat_B[146][0] +
                mat_A[76][3] * mat_B[154][0] +
                mat_A[77][0] * mat_B[162][0] +
                mat_A[77][1] * mat_B[170][0] +
                mat_A[77][2] * mat_B[178][0] +
                mat_A[77][3] * mat_B[186][0] +
                mat_A[78][0] * mat_B[194][0] +
                mat_A[78][1] * mat_B[202][0] +
                mat_A[78][2] * mat_B[210][0] +
                mat_A[78][3] * mat_B[218][0] +
                mat_A[79][0] * mat_B[226][0] +
                mat_A[79][1] * mat_B[234][0] +
                mat_A[79][2] * mat_B[242][0] +
                mat_A[79][3] * mat_B[250][0];
    mat_C[74][1] <=
                mat_A[72][0] * mat_B[2][1] +
                mat_A[72][1] * mat_B[10][1] +
                mat_A[72][2] * mat_B[18][1] +
                mat_A[72][3] * mat_B[26][1] +
                mat_A[73][0] * mat_B[34][1] +
                mat_A[73][1] * mat_B[42][1] +
                mat_A[73][2] * mat_B[50][1] +
                mat_A[73][3] * mat_B[58][1] +
                mat_A[74][0] * mat_B[66][1] +
                mat_A[74][1] * mat_B[74][1] +
                mat_A[74][2] * mat_B[82][1] +
                mat_A[74][3] * mat_B[90][1] +
                mat_A[75][0] * mat_B[98][1] +
                mat_A[75][1] * mat_B[106][1] +
                mat_A[75][2] * mat_B[114][1] +
                mat_A[75][3] * mat_B[122][1] +
                mat_A[76][0] * mat_B[130][1] +
                mat_A[76][1] * mat_B[138][1] +
                mat_A[76][2] * mat_B[146][1] +
                mat_A[76][3] * mat_B[154][1] +
                mat_A[77][0] * mat_B[162][1] +
                mat_A[77][1] * mat_B[170][1] +
                mat_A[77][2] * mat_B[178][1] +
                mat_A[77][3] * mat_B[186][1] +
                mat_A[78][0] * mat_B[194][1] +
                mat_A[78][1] * mat_B[202][1] +
                mat_A[78][2] * mat_B[210][1] +
                mat_A[78][3] * mat_B[218][1] +
                mat_A[79][0] * mat_B[226][1] +
                mat_A[79][1] * mat_B[234][1] +
                mat_A[79][2] * mat_B[242][1] +
                mat_A[79][3] * mat_B[250][1];
    mat_C[74][2] <=
                mat_A[72][0] * mat_B[2][2] +
                mat_A[72][1] * mat_B[10][2] +
                mat_A[72][2] * mat_B[18][2] +
                mat_A[72][3] * mat_B[26][2] +
                mat_A[73][0] * mat_B[34][2] +
                mat_A[73][1] * mat_B[42][2] +
                mat_A[73][2] * mat_B[50][2] +
                mat_A[73][3] * mat_B[58][2] +
                mat_A[74][0] * mat_B[66][2] +
                mat_A[74][1] * mat_B[74][2] +
                mat_A[74][2] * mat_B[82][2] +
                mat_A[74][3] * mat_B[90][2] +
                mat_A[75][0] * mat_B[98][2] +
                mat_A[75][1] * mat_B[106][2] +
                mat_A[75][2] * mat_B[114][2] +
                mat_A[75][3] * mat_B[122][2] +
                mat_A[76][0] * mat_B[130][2] +
                mat_A[76][1] * mat_B[138][2] +
                mat_A[76][2] * mat_B[146][2] +
                mat_A[76][3] * mat_B[154][2] +
                mat_A[77][0] * mat_B[162][2] +
                mat_A[77][1] * mat_B[170][2] +
                mat_A[77][2] * mat_B[178][2] +
                mat_A[77][3] * mat_B[186][2] +
                mat_A[78][0] * mat_B[194][2] +
                mat_A[78][1] * mat_B[202][2] +
                mat_A[78][2] * mat_B[210][2] +
                mat_A[78][3] * mat_B[218][2] +
                mat_A[79][0] * mat_B[226][2] +
                mat_A[79][1] * mat_B[234][2] +
                mat_A[79][2] * mat_B[242][2] +
                mat_A[79][3] * mat_B[250][2];
    mat_C[74][3] <=
                mat_A[72][0] * mat_B[2][3] +
                mat_A[72][1] * mat_B[10][3] +
                mat_A[72][2] * mat_B[18][3] +
                mat_A[72][3] * mat_B[26][3] +
                mat_A[73][0] * mat_B[34][3] +
                mat_A[73][1] * mat_B[42][3] +
                mat_A[73][2] * mat_B[50][3] +
                mat_A[73][3] * mat_B[58][3] +
                mat_A[74][0] * mat_B[66][3] +
                mat_A[74][1] * mat_B[74][3] +
                mat_A[74][2] * mat_B[82][3] +
                mat_A[74][3] * mat_B[90][3] +
                mat_A[75][0] * mat_B[98][3] +
                mat_A[75][1] * mat_B[106][3] +
                mat_A[75][2] * mat_B[114][3] +
                mat_A[75][3] * mat_B[122][3] +
                mat_A[76][0] * mat_B[130][3] +
                mat_A[76][1] * mat_B[138][3] +
                mat_A[76][2] * mat_B[146][3] +
                mat_A[76][3] * mat_B[154][3] +
                mat_A[77][0] * mat_B[162][3] +
                mat_A[77][1] * mat_B[170][3] +
                mat_A[77][2] * mat_B[178][3] +
                mat_A[77][3] * mat_B[186][3] +
                mat_A[78][0] * mat_B[194][3] +
                mat_A[78][1] * mat_B[202][3] +
                mat_A[78][2] * mat_B[210][3] +
                mat_A[78][3] * mat_B[218][3] +
                mat_A[79][0] * mat_B[226][3] +
                mat_A[79][1] * mat_B[234][3] +
                mat_A[79][2] * mat_B[242][3] +
                mat_A[79][3] * mat_B[250][3];
    mat_C[75][0] <=
                mat_A[72][0] * mat_B[3][0] +
                mat_A[72][1] * mat_B[11][0] +
                mat_A[72][2] * mat_B[19][0] +
                mat_A[72][3] * mat_B[27][0] +
                mat_A[73][0] * mat_B[35][0] +
                mat_A[73][1] * mat_B[43][0] +
                mat_A[73][2] * mat_B[51][0] +
                mat_A[73][3] * mat_B[59][0] +
                mat_A[74][0] * mat_B[67][0] +
                mat_A[74][1] * mat_B[75][0] +
                mat_A[74][2] * mat_B[83][0] +
                mat_A[74][3] * mat_B[91][0] +
                mat_A[75][0] * mat_B[99][0] +
                mat_A[75][1] * mat_B[107][0] +
                mat_A[75][2] * mat_B[115][0] +
                mat_A[75][3] * mat_B[123][0] +
                mat_A[76][0] * mat_B[131][0] +
                mat_A[76][1] * mat_B[139][0] +
                mat_A[76][2] * mat_B[147][0] +
                mat_A[76][3] * mat_B[155][0] +
                mat_A[77][0] * mat_B[163][0] +
                mat_A[77][1] * mat_B[171][0] +
                mat_A[77][2] * mat_B[179][0] +
                mat_A[77][3] * mat_B[187][0] +
                mat_A[78][0] * mat_B[195][0] +
                mat_A[78][1] * mat_B[203][0] +
                mat_A[78][2] * mat_B[211][0] +
                mat_A[78][3] * mat_B[219][0] +
                mat_A[79][0] * mat_B[227][0] +
                mat_A[79][1] * mat_B[235][0] +
                mat_A[79][2] * mat_B[243][0] +
                mat_A[79][3] * mat_B[251][0];
    mat_C[75][1] <=
                mat_A[72][0] * mat_B[3][1] +
                mat_A[72][1] * mat_B[11][1] +
                mat_A[72][2] * mat_B[19][1] +
                mat_A[72][3] * mat_B[27][1] +
                mat_A[73][0] * mat_B[35][1] +
                mat_A[73][1] * mat_B[43][1] +
                mat_A[73][2] * mat_B[51][1] +
                mat_A[73][3] * mat_B[59][1] +
                mat_A[74][0] * mat_B[67][1] +
                mat_A[74][1] * mat_B[75][1] +
                mat_A[74][2] * mat_B[83][1] +
                mat_A[74][3] * mat_B[91][1] +
                mat_A[75][0] * mat_B[99][1] +
                mat_A[75][1] * mat_B[107][1] +
                mat_A[75][2] * mat_B[115][1] +
                mat_A[75][3] * mat_B[123][1] +
                mat_A[76][0] * mat_B[131][1] +
                mat_A[76][1] * mat_B[139][1] +
                mat_A[76][2] * mat_B[147][1] +
                mat_A[76][3] * mat_B[155][1] +
                mat_A[77][0] * mat_B[163][1] +
                mat_A[77][1] * mat_B[171][1] +
                mat_A[77][2] * mat_B[179][1] +
                mat_A[77][3] * mat_B[187][1] +
                mat_A[78][0] * mat_B[195][1] +
                mat_A[78][1] * mat_B[203][1] +
                mat_A[78][2] * mat_B[211][1] +
                mat_A[78][3] * mat_B[219][1] +
                mat_A[79][0] * mat_B[227][1] +
                mat_A[79][1] * mat_B[235][1] +
                mat_A[79][2] * mat_B[243][1] +
                mat_A[79][3] * mat_B[251][1];
    mat_C[75][2] <=
                mat_A[72][0] * mat_B[3][2] +
                mat_A[72][1] * mat_B[11][2] +
                mat_A[72][2] * mat_B[19][2] +
                mat_A[72][3] * mat_B[27][2] +
                mat_A[73][0] * mat_B[35][2] +
                mat_A[73][1] * mat_B[43][2] +
                mat_A[73][2] * mat_B[51][2] +
                mat_A[73][3] * mat_B[59][2] +
                mat_A[74][0] * mat_B[67][2] +
                mat_A[74][1] * mat_B[75][2] +
                mat_A[74][2] * mat_B[83][2] +
                mat_A[74][3] * mat_B[91][2] +
                mat_A[75][0] * mat_B[99][2] +
                mat_A[75][1] * mat_B[107][2] +
                mat_A[75][2] * mat_B[115][2] +
                mat_A[75][3] * mat_B[123][2] +
                mat_A[76][0] * mat_B[131][2] +
                mat_A[76][1] * mat_B[139][2] +
                mat_A[76][2] * mat_B[147][2] +
                mat_A[76][3] * mat_B[155][2] +
                mat_A[77][0] * mat_B[163][2] +
                mat_A[77][1] * mat_B[171][2] +
                mat_A[77][2] * mat_B[179][2] +
                mat_A[77][3] * mat_B[187][2] +
                mat_A[78][0] * mat_B[195][2] +
                mat_A[78][1] * mat_B[203][2] +
                mat_A[78][2] * mat_B[211][2] +
                mat_A[78][3] * mat_B[219][2] +
                mat_A[79][0] * mat_B[227][2] +
                mat_A[79][1] * mat_B[235][2] +
                mat_A[79][2] * mat_B[243][2] +
                mat_A[79][3] * mat_B[251][2];
    mat_C[75][3] <=
                mat_A[72][0] * mat_B[3][3] +
                mat_A[72][1] * mat_B[11][3] +
                mat_A[72][2] * mat_B[19][3] +
                mat_A[72][3] * mat_B[27][3] +
                mat_A[73][0] * mat_B[35][3] +
                mat_A[73][1] * mat_B[43][3] +
                mat_A[73][2] * mat_B[51][3] +
                mat_A[73][3] * mat_B[59][3] +
                mat_A[74][0] * mat_B[67][3] +
                mat_A[74][1] * mat_B[75][3] +
                mat_A[74][2] * mat_B[83][3] +
                mat_A[74][3] * mat_B[91][3] +
                mat_A[75][0] * mat_B[99][3] +
                mat_A[75][1] * mat_B[107][3] +
                mat_A[75][2] * mat_B[115][3] +
                mat_A[75][3] * mat_B[123][3] +
                mat_A[76][0] * mat_B[131][3] +
                mat_A[76][1] * mat_B[139][3] +
                mat_A[76][2] * mat_B[147][3] +
                mat_A[76][3] * mat_B[155][3] +
                mat_A[77][0] * mat_B[163][3] +
                mat_A[77][1] * mat_B[171][3] +
                mat_A[77][2] * mat_B[179][3] +
                mat_A[77][3] * mat_B[187][3] +
                mat_A[78][0] * mat_B[195][3] +
                mat_A[78][1] * mat_B[203][3] +
                mat_A[78][2] * mat_B[211][3] +
                mat_A[78][3] * mat_B[219][3] +
                mat_A[79][0] * mat_B[227][3] +
                mat_A[79][1] * mat_B[235][3] +
                mat_A[79][2] * mat_B[243][3] +
                mat_A[79][3] * mat_B[251][3];
    mat_C[76][0] <=
                mat_A[72][0] * mat_B[4][0] +
                mat_A[72][1] * mat_B[12][0] +
                mat_A[72][2] * mat_B[20][0] +
                mat_A[72][3] * mat_B[28][0] +
                mat_A[73][0] * mat_B[36][0] +
                mat_A[73][1] * mat_B[44][0] +
                mat_A[73][2] * mat_B[52][0] +
                mat_A[73][3] * mat_B[60][0] +
                mat_A[74][0] * mat_B[68][0] +
                mat_A[74][1] * mat_B[76][0] +
                mat_A[74][2] * mat_B[84][0] +
                mat_A[74][3] * mat_B[92][0] +
                mat_A[75][0] * mat_B[100][0] +
                mat_A[75][1] * mat_B[108][0] +
                mat_A[75][2] * mat_B[116][0] +
                mat_A[75][3] * mat_B[124][0] +
                mat_A[76][0] * mat_B[132][0] +
                mat_A[76][1] * mat_B[140][0] +
                mat_A[76][2] * mat_B[148][0] +
                mat_A[76][3] * mat_B[156][0] +
                mat_A[77][0] * mat_B[164][0] +
                mat_A[77][1] * mat_B[172][0] +
                mat_A[77][2] * mat_B[180][0] +
                mat_A[77][3] * mat_B[188][0] +
                mat_A[78][0] * mat_B[196][0] +
                mat_A[78][1] * mat_B[204][0] +
                mat_A[78][2] * mat_B[212][0] +
                mat_A[78][3] * mat_B[220][0] +
                mat_A[79][0] * mat_B[228][0] +
                mat_A[79][1] * mat_B[236][0] +
                mat_A[79][2] * mat_B[244][0] +
                mat_A[79][3] * mat_B[252][0];
    mat_C[76][1] <=
                mat_A[72][0] * mat_B[4][1] +
                mat_A[72][1] * mat_B[12][1] +
                mat_A[72][2] * mat_B[20][1] +
                mat_A[72][3] * mat_B[28][1] +
                mat_A[73][0] * mat_B[36][1] +
                mat_A[73][1] * mat_B[44][1] +
                mat_A[73][2] * mat_B[52][1] +
                mat_A[73][3] * mat_B[60][1] +
                mat_A[74][0] * mat_B[68][1] +
                mat_A[74][1] * mat_B[76][1] +
                mat_A[74][2] * mat_B[84][1] +
                mat_A[74][3] * mat_B[92][1] +
                mat_A[75][0] * mat_B[100][1] +
                mat_A[75][1] * mat_B[108][1] +
                mat_A[75][2] * mat_B[116][1] +
                mat_A[75][3] * mat_B[124][1] +
                mat_A[76][0] * mat_B[132][1] +
                mat_A[76][1] * mat_B[140][1] +
                mat_A[76][2] * mat_B[148][1] +
                mat_A[76][3] * mat_B[156][1] +
                mat_A[77][0] * mat_B[164][1] +
                mat_A[77][1] * mat_B[172][1] +
                mat_A[77][2] * mat_B[180][1] +
                mat_A[77][3] * mat_B[188][1] +
                mat_A[78][0] * mat_B[196][1] +
                mat_A[78][1] * mat_B[204][1] +
                mat_A[78][2] * mat_B[212][1] +
                mat_A[78][3] * mat_B[220][1] +
                mat_A[79][0] * mat_B[228][1] +
                mat_A[79][1] * mat_B[236][1] +
                mat_A[79][2] * mat_B[244][1] +
                mat_A[79][3] * mat_B[252][1];
    mat_C[76][2] <=
                mat_A[72][0] * mat_B[4][2] +
                mat_A[72][1] * mat_B[12][2] +
                mat_A[72][2] * mat_B[20][2] +
                mat_A[72][3] * mat_B[28][2] +
                mat_A[73][0] * mat_B[36][2] +
                mat_A[73][1] * mat_B[44][2] +
                mat_A[73][2] * mat_B[52][2] +
                mat_A[73][3] * mat_B[60][2] +
                mat_A[74][0] * mat_B[68][2] +
                mat_A[74][1] * mat_B[76][2] +
                mat_A[74][2] * mat_B[84][2] +
                mat_A[74][3] * mat_B[92][2] +
                mat_A[75][0] * mat_B[100][2] +
                mat_A[75][1] * mat_B[108][2] +
                mat_A[75][2] * mat_B[116][2] +
                mat_A[75][3] * mat_B[124][2] +
                mat_A[76][0] * mat_B[132][2] +
                mat_A[76][1] * mat_B[140][2] +
                mat_A[76][2] * mat_B[148][2] +
                mat_A[76][3] * mat_B[156][2] +
                mat_A[77][0] * mat_B[164][2] +
                mat_A[77][1] * mat_B[172][2] +
                mat_A[77][2] * mat_B[180][2] +
                mat_A[77][3] * mat_B[188][2] +
                mat_A[78][0] * mat_B[196][2] +
                mat_A[78][1] * mat_B[204][2] +
                mat_A[78][2] * mat_B[212][2] +
                mat_A[78][3] * mat_B[220][2] +
                mat_A[79][0] * mat_B[228][2] +
                mat_A[79][1] * mat_B[236][2] +
                mat_A[79][2] * mat_B[244][2] +
                mat_A[79][3] * mat_B[252][2];
    mat_C[76][3] <=
                mat_A[72][0] * mat_B[4][3] +
                mat_A[72][1] * mat_B[12][3] +
                mat_A[72][2] * mat_B[20][3] +
                mat_A[72][3] * mat_B[28][3] +
                mat_A[73][0] * mat_B[36][3] +
                mat_A[73][1] * mat_B[44][3] +
                mat_A[73][2] * mat_B[52][3] +
                mat_A[73][3] * mat_B[60][3] +
                mat_A[74][0] * mat_B[68][3] +
                mat_A[74][1] * mat_B[76][3] +
                mat_A[74][2] * mat_B[84][3] +
                mat_A[74][3] * mat_B[92][3] +
                mat_A[75][0] * mat_B[100][3] +
                mat_A[75][1] * mat_B[108][3] +
                mat_A[75][2] * mat_B[116][3] +
                mat_A[75][3] * mat_B[124][3] +
                mat_A[76][0] * mat_B[132][3] +
                mat_A[76][1] * mat_B[140][3] +
                mat_A[76][2] * mat_B[148][3] +
                mat_A[76][3] * mat_B[156][3] +
                mat_A[77][0] * mat_B[164][3] +
                mat_A[77][1] * mat_B[172][3] +
                mat_A[77][2] * mat_B[180][3] +
                mat_A[77][3] * mat_B[188][3] +
                mat_A[78][0] * mat_B[196][3] +
                mat_A[78][1] * mat_B[204][3] +
                mat_A[78][2] * mat_B[212][3] +
                mat_A[78][3] * mat_B[220][3] +
                mat_A[79][0] * mat_B[228][3] +
                mat_A[79][1] * mat_B[236][3] +
                mat_A[79][2] * mat_B[244][3] +
                mat_A[79][3] * mat_B[252][3];
    mat_C[77][0] <=
                mat_A[72][0] * mat_B[5][0] +
                mat_A[72][1] * mat_B[13][0] +
                mat_A[72][2] * mat_B[21][0] +
                mat_A[72][3] * mat_B[29][0] +
                mat_A[73][0] * mat_B[37][0] +
                mat_A[73][1] * mat_B[45][0] +
                mat_A[73][2] * mat_B[53][0] +
                mat_A[73][3] * mat_B[61][0] +
                mat_A[74][0] * mat_B[69][0] +
                mat_A[74][1] * mat_B[77][0] +
                mat_A[74][2] * mat_B[85][0] +
                mat_A[74][3] * mat_B[93][0] +
                mat_A[75][0] * mat_B[101][0] +
                mat_A[75][1] * mat_B[109][0] +
                mat_A[75][2] * mat_B[117][0] +
                mat_A[75][3] * mat_B[125][0] +
                mat_A[76][0] * mat_B[133][0] +
                mat_A[76][1] * mat_B[141][0] +
                mat_A[76][2] * mat_B[149][0] +
                mat_A[76][3] * mat_B[157][0] +
                mat_A[77][0] * mat_B[165][0] +
                mat_A[77][1] * mat_B[173][0] +
                mat_A[77][2] * mat_B[181][0] +
                mat_A[77][3] * mat_B[189][0] +
                mat_A[78][0] * mat_B[197][0] +
                mat_A[78][1] * mat_B[205][0] +
                mat_A[78][2] * mat_B[213][0] +
                mat_A[78][3] * mat_B[221][0] +
                mat_A[79][0] * mat_B[229][0] +
                mat_A[79][1] * mat_B[237][0] +
                mat_A[79][2] * mat_B[245][0] +
                mat_A[79][3] * mat_B[253][0];
    mat_C[77][1] <=
                mat_A[72][0] * mat_B[5][1] +
                mat_A[72][1] * mat_B[13][1] +
                mat_A[72][2] * mat_B[21][1] +
                mat_A[72][3] * mat_B[29][1] +
                mat_A[73][0] * mat_B[37][1] +
                mat_A[73][1] * mat_B[45][1] +
                mat_A[73][2] * mat_B[53][1] +
                mat_A[73][3] * mat_B[61][1] +
                mat_A[74][0] * mat_B[69][1] +
                mat_A[74][1] * mat_B[77][1] +
                mat_A[74][2] * mat_B[85][1] +
                mat_A[74][3] * mat_B[93][1] +
                mat_A[75][0] * mat_B[101][1] +
                mat_A[75][1] * mat_B[109][1] +
                mat_A[75][2] * mat_B[117][1] +
                mat_A[75][3] * mat_B[125][1] +
                mat_A[76][0] * mat_B[133][1] +
                mat_A[76][1] * mat_B[141][1] +
                mat_A[76][2] * mat_B[149][1] +
                mat_A[76][3] * mat_B[157][1] +
                mat_A[77][0] * mat_B[165][1] +
                mat_A[77][1] * mat_B[173][1] +
                mat_A[77][2] * mat_B[181][1] +
                mat_A[77][3] * mat_B[189][1] +
                mat_A[78][0] * mat_B[197][1] +
                mat_A[78][1] * mat_B[205][1] +
                mat_A[78][2] * mat_B[213][1] +
                mat_A[78][3] * mat_B[221][1] +
                mat_A[79][0] * mat_B[229][1] +
                mat_A[79][1] * mat_B[237][1] +
                mat_A[79][2] * mat_B[245][1] +
                mat_A[79][3] * mat_B[253][1];
    mat_C[77][2] <=
                mat_A[72][0] * mat_B[5][2] +
                mat_A[72][1] * mat_B[13][2] +
                mat_A[72][2] * mat_B[21][2] +
                mat_A[72][3] * mat_B[29][2] +
                mat_A[73][0] * mat_B[37][2] +
                mat_A[73][1] * mat_B[45][2] +
                mat_A[73][2] * mat_B[53][2] +
                mat_A[73][3] * mat_B[61][2] +
                mat_A[74][0] * mat_B[69][2] +
                mat_A[74][1] * mat_B[77][2] +
                mat_A[74][2] * mat_B[85][2] +
                mat_A[74][3] * mat_B[93][2] +
                mat_A[75][0] * mat_B[101][2] +
                mat_A[75][1] * mat_B[109][2] +
                mat_A[75][2] * mat_B[117][2] +
                mat_A[75][3] * mat_B[125][2] +
                mat_A[76][0] * mat_B[133][2] +
                mat_A[76][1] * mat_B[141][2] +
                mat_A[76][2] * mat_B[149][2] +
                mat_A[76][3] * mat_B[157][2] +
                mat_A[77][0] * mat_B[165][2] +
                mat_A[77][1] * mat_B[173][2] +
                mat_A[77][2] * mat_B[181][2] +
                mat_A[77][3] * mat_B[189][2] +
                mat_A[78][0] * mat_B[197][2] +
                mat_A[78][1] * mat_B[205][2] +
                mat_A[78][2] * mat_B[213][2] +
                mat_A[78][3] * mat_B[221][2] +
                mat_A[79][0] * mat_B[229][2] +
                mat_A[79][1] * mat_B[237][2] +
                mat_A[79][2] * mat_B[245][2] +
                mat_A[79][3] * mat_B[253][2];
    mat_C[77][3] <=
                mat_A[72][0] * mat_B[5][3] +
                mat_A[72][1] * mat_B[13][3] +
                mat_A[72][2] * mat_B[21][3] +
                mat_A[72][3] * mat_B[29][3] +
                mat_A[73][0] * mat_B[37][3] +
                mat_A[73][1] * mat_B[45][3] +
                mat_A[73][2] * mat_B[53][3] +
                mat_A[73][3] * mat_B[61][3] +
                mat_A[74][0] * mat_B[69][3] +
                mat_A[74][1] * mat_B[77][3] +
                mat_A[74][2] * mat_B[85][3] +
                mat_A[74][3] * mat_B[93][3] +
                mat_A[75][0] * mat_B[101][3] +
                mat_A[75][1] * mat_B[109][3] +
                mat_A[75][2] * mat_B[117][3] +
                mat_A[75][3] * mat_B[125][3] +
                mat_A[76][0] * mat_B[133][3] +
                mat_A[76][1] * mat_B[141][3] +
                mat_A[76][2] * mat_B[149][3] +
                mat_A[76][3] * mat_B[157][3] +
                mat_A[77][0] * mat_B[165][3] +
                mat_A[77][1] * mat_B[173][3] +
                mat_A[77][2] * mat_B[181][3] +
                mat_A[77][3] * mat_B[189][3] +
                mat_A[78][0] * mat_B[197][3] +
                mat_A[78][1] * mat_B[205][3] +
                mat_A[78][2] * mat_B[213][3] +
                mat_A[78][3] * mat_B[221][3] +
                mat_A[79][0] * mat_B[229][3] +
                mat_A[79][1] * mat_B[237][3] +
                mat_A[79][2] * mat_B[245][3] +
                mat_A[79][3] * mat_B[253][3];
    mat_C[78][0] <=
                mat_A[72][0] * mat_B[6][0] +
                mat_A[72][1] * mat_B[14][0] +
                mat_A[72][2] * mat_B[22][0] +
                mat_A[72][3] * mat_B[30][0] +
                mat_A[73][0] * mat_B[38][0] +
                mat_A[73][1] * mat_B[46][0] +
                mat_A[73][2] * mat_B[54][0] +
                mat_A[73][3] * mat_B[62][0] +
                mat_A[74][0] * mat_B[70][0] +
                mat_A[74][1] * mat_B[78][0] +
                mat_A[74][2] * mat_B[86][0] +
                mat_A[74][3] * mat_B[94][0] +
                mat_A[75][0] * mat_B[102][0] +
                mat_A[75][1] * mat_B[110][0] +
                mat_A[75][2] * mat_B[118][0] +
                mat_A[75][3] * mat_B[126][0] +
                mat_A[76][0] * mat_B[134][0] +
                mat_A[76][1] * mat_B[142][0] +
                mat_A[76][2] * mat_B[150][0] +
                mat_A[76][3] * mat_B[158][0] +
                mat_A[77][0] * mat_B[166][0] +
                mat_A[77][1] * mat_B[174][0] +
                mat_A[77][2] * mat_B[182][0] +
                mat_A[77][3] * mat_B[190][0] +
                mat_A[78][0] * mat_B[198][0] +
                mat_A[78][1] * mat_B[206][0] +
                mat_A[78][2] * mat_B[214][0] +
                mat_A[78][3] * mat_B[222][0] +
                mat_A[79][0] * mat_B[230][0] +
                mat_A[79][1] * mat_B[238][0] +
                mat_A[79][2] * mat_B[246][0] +
                mat_A[79][3] * mat_B[254][0];
    mat_C[78][1] <=
                mat_A[72][0] * mat_B[6][1] +
                mat_A[72][1] * mat_B[14][1] +
                mat_A[72][2] * mat_B[22][1] +
                mat_A[72][3] * mat_B[30][1] +
                mat_A[73][0] * mat_B[38][1] +
                mat_A[73][1] * mat_B[46][1] +
                mat_A[73][2] * mat_B[54][1] +
                mat_A[73][3] * mat_B[62][1] +
                mat_A[74][0] * mat_B[70][1] +
                mat_A[74][1] * mat_B[78][1] +
                mat_A[74][2] * mat_B[86][1] +
                mat_A[74][3] * mat_B[94][1] +
                mat_A[75][0] * mat_B[102][1] +
                mat_A[75][1] * mat_B[110][1] +
                mat_A[75][2] * mat_B[118][1] +
                mat_A[75][3] * mat_B[126][1] +
                mat_A[76][0] * mat_B[134][1] +
                mat_A[76][1] * mat_B[142][1] +
                mat_A[76][2] * mat_B[150][1] +
                mat_A[76][3] * mat_B[158][1] +
                mat_A[77][0] * mat_B[166][1] +
                mat_A[77][1] * mat_B[174][1] +
                mat_A[77][2] * mat_B[182][1] +
                mat_A[77][3] * mat_B[190][1] +
                mat_A[78][0] * mat_B[198][1] +
                mat_A[78][1] * mat_B[206][1] +
                mat_A[78][2] * mat_B[214][1] +
                mat_A[78][3] * mat_B[222][1] +
                mat_A[79][0] * mat_B[230][1] +
                mat_A[79][1] * mat_B[238][1] +
                mat_A[79][2] * mat_B[246][1] +
                mat_A[79][3] * mat_B[254][1];
    mat_C[78][2] <=
                mat_A[72][0] * mat_B[6][2] +
                mat_A[72][1] * mat_B[14][2] +
                mat_A[72][2] * mat_B[22][2] +
                mat_A[72][3] * mat_B[30][2] +
                mat_A[73][0] * mat_B[38][2] +
                mat_A[73][1] * mat_B[46][2] +
                mat_A[73][2] * mat_B[54][2] +
                mat_A[73][3] * mat_B[62][2] +
                mat_A[74][0] * mat_B[70][2] +
                mat_A[74][1] * mat_B[78][2] +
                mat_A[74][2] * mat_B[86][2] +
                mat_A[74][3] * mat_B[94][2] +
                mat_A[75][0] * mat_B[102][2] +
                mat_A[75][1] * mat_B[110][2] +
                mat_A[75][2] * mat_B[118][2] +
                mat_A[75][3] * mat_B[126][2] +
                mat_A[76][0] * mat_B[134][2] +
                mat_A[76][1] * mat_B[142][2] +
                mat_A[76][2] * mat_B[150][2] +
                mat_A[76][3] * mat_B[158][2] +
                mat_A[77][0] * mat_B[166][2] +
                mat_A[77][1] * mat_B[174][2] +
                mat_A[77][2] * mat_B[182][2] +
                mat_A[77][3] * mat_B[190][2] +
                mat_A[78][0] * mat_B[198][2] +
                mat_A[78][1] * mat_B[206][2] +
                mat_A[78][2] * mat_B[214][2] +
                mat_A[78][3] * mat_B[222][2] +
                mat_A[79][0] * mat_B[230][2] +
                mat_A[79][1] * mat_B[238][2] +
                mat_A[79][2] * mat_B[246][2] +
                mat_A[79][3] * mat_B[254][2];
    mat_C[78][3] <=
                mat_A[72][0] * mat_B[6][3] +
                mat_A[72][1] * mat_B[14][3] +
                mat_A[72][2] * mat_B[22][3] +
                mat_A[72][3] * mat_B[30][3] +
                mat_A[73][0] * mat_B[38][3] +
                mat_A[73][1] * mat_B[46][3] +
                mat_A[73][2] * mat_B[54][3] +
                mat_A[73][3] * mat_B[62][3] +
                mat_A[74][0] * mat_B[70][3] +
                mat_A[74][1] * mat_B[78][3] +
                mat_A[74][2] * mat_B[86][3] +
                mat_A[74][3] * mat_B[94][3] +
                mat_A[75][0] * mat_B[102][3] +
                mat_A[75][1] * mat_B[110][3] +
                mat_A[75][2] * mat_B[118][3] +
                mat_A[75][3] * mat_B[126][3] +
                mat_A[76][0] * mat_B[134][3] +
                mat_A[76][1] * mat_B[142][3] +
                mat_A[76][2] * mat_B[150][3] +
                mat_A[76][3] * mat_B[158][3] +
                mat_A[77][0] * mat_B[166][3] +
                mat_A[77][1] * mat_B[174][3] +
                mat_A[77][2] * mat_B[182][3] +
                mat_A[77][3] * mat_B[190][3] +
                mat_A[78][0] * mat_B[198][3] +
                mat_A[78][1] * mat_B[206][3] +
                mat_A[78][2] * mat_B[214][3] +
                mat_A[78][3] * mat_B[222][3] +
                mat_A[79][0] * mat_B[230][3] +
                mat_A[79][1] * mat_B[238][3] +
                mat_A[79][2] * mat_B[246][3] +
                mat_A[79][3] * mat_B[254][3];
    mat_C[79][0] <=
                mat_A[72][0] * mat_B[7][0] +
                mat_A[72][1] * mat_B[15][0] +
                mat_A[72][2] * mat_B[23][0] +
                mat_A[72][3] * mat_B[31][0] +
                mat_A[73][0] * mat_B[39][0] +
                mat_A[73][1] * mat_B[47][0] +
                mat_A[73][2] * mat_B[55][0] +
                mat_A[73][3] * mat_B[63][0] +
                mat_A[74][0] * mat_B[71][0] +
                mat_A[74][1] * mat_B[79][0] +
                mat_A[74][2] * mat_B[87][0] +
                mat_A[74][3] * mat_B[95][0] +
                mat_A[75][0] * mat_B[103][0] +
                mat_A[75][1] * mat_B[111][0] +
                mat_A[75][2] * mat_B[119][0] +
                mat_A[75][3] * mat_B[127][0] +
                mat_A[76][0] * mat_B[135][0] +
                mat_A[76][1] * mat_B[143][0] +
                mat_A[76][2] * mat_B[151][0] +
                mat_A[76][3] * mat_B[159][0] +
                mat_A[77][0] * mat_B[167][0] +
                mat_A[77][1] * mat_B[175][0] +
                mat_A[77][2] * mat_B[183][0] +
                mat_A[77][3] * mat_B[191][0] +
                mat_A[78][0] * mat_B[199][0] +
                mat_A[78][1] * mat_B[207][0] +
                mat_A[78][2] * mat_B[215][0] +
                mat_A[78][3] * mat_B[223][0] +
                mat_A[79][0] * mat_B[231][0] +
                mat_A[79][1] * mat_B[239][0] +
                mat_A[79][2] * mat_B[247][0] +
                mat_A[79][3] * mat_B[255][0];
    mat_C[79][1] <=
                mat_A[72][0] * mat_B[7][1] +
                mat_A[72][1] * mat_B[15][1] +
                mat_A[72][2] * mat_B[23][1] +
                mat_A[72][3] * mat_B[31][1] +
                mat_A[73][0] * mat_B[39][1] +
                mat_A[73][1] * mat_B[47][1] +
                mat_A[73][2] * mat_B[55][1] +
                mat_A[73][3] * mat_B[63][1] +
                mat_A[74][0] * mat_B[71][1] +
                mat_A[74][1] * mat_B[79][1] +
                mat_A[74][2] * mat_B[87][1] +
                mat_A[74][3] * mat_B[95][1] +
                mat_A[75][0] * mat_B[103][1] +
                mat_A[75][1] * mat_B[111][1] +
                mat_A[75][2] * mat_B[119][1] +
                mat_A[75][3] * mat_B[127][1] +
                mat_A[76][0] * mat_B[135][1] +
                mat_A[76][1] * mat_B[143][1] +
                mat_A[76][2] * mat_B[151][1] +
                mat_A[76][3] * mat_B[159][1] +
                mat_A[77][0] * mat_B[167][1] +
                mat_A[77][1] * mat_B[175][1] +
                mat_A[77][2] * mat_B[183][1] +
                mat_A[77][3] * mat_B[191][1] +
                mat_A[78][0] * mat_B[199][1] +
                mat_A[78][1] * mat_B[207][1] +
                mat_A[78][2] * mat_B[215][1] +
                mat_A[78][3] * mat_B[223][1] +
                mat_A[79][0] * mat_B[231][1] +
                mat_A[79][1] * mat_B[239][1] +
                mat_A[79][2] * mat_B[247][1] +
                mat_A[79][3] * mat_B[255][1];
    mat_C[79][2] <=
                mat_A[72][0] * mat_B[7][2] +
                mat_A[72][1] * mat_B[15][2] +
                mat_A[72][2] * mat_B[23][2] +
                mat_A[72][3] * mat_B[31][2] +
                mat_A[73][0] * mat_B[39][2] +
                mat_A[73][1] * mat_B[47][2] +
                mat_A[73][2] * mat_B[55][2] +
                mat_A[73][3] * mat_B[63][2] +
                mat_A[74][0] * mat_B[71][2] +
                mat_A[74][1] * mat_B[79][2] +
                mat_A[74][2] * mat_B[87][2] +
                mat_A[74][3] * mat_B[95][2] +
                mat_A[75][0] * mat_B[103][2] +
                mat_A[75][1] * mat_B[111][2] +
                mat_A[75][2] * mat_B[119][2] +
                mat_A[75][3] * mat_B[127][2] +
                mat_A[76][0] * mat_B[135][2] +
                mat_A[76][1] * mat_B[143][2] +
                mat_A[76][2] * mat_B[151][2] +
                mat_A[76][3] * mat_B[159][2] +
                mat_A[77][0] * mat_B[167][2] +
                mat_A[77][1] * mat_B[175][2] +
                mat_A[77][2] * mat_B[183][2] +
                mat_A[77][3] * mat_B[191][2] +
                mat_A[78][0] * mat_B[199][2] +
                mat_A[78][1] * mat_B[207][2] +
                mat_A[78][2] * mat_B[215][2] +
                mat_A[78][3] * mat_B[223][2] +
                mat_A[79][0] * mat_B[231][2] +
                mat_A[79][1] * mat_B[239][2] +
                mat_A[79][2] * mat_B[247][2] +
                mat_A[79][3] * mat_B[255][2];
    mat_C[79][3] <=
                mat_A[72][0] * mat_B[7][3] +
                mat_A[72][1] * mat_B[15][3] +
                mat_A[72][2] * mat_B[23][3] +
                mat_A[72][3] * mat_B[31][3] +
                mat_A[73][0] * mat_B[39][3] +
                mat_A[73][1] * mat_B[47][3] +
                mat_A[73][2] * mat_B[55][3] +
                mat_A[73][3] * mat_B[63][3] +
                mat_A[74][0] * mat_B[71][3] +
                mat_A[74][1] * mat_B[79][3] +
                mat_A[74][2] * mat_B[87][3] +
                mat_A[74][3] * mat_B[95][3] +
                mat_A[75][0] * mat_B[103][3] +
                mat_A[75][1] * mat_B[111][3] +
                mat_A[75][2] * mat_B[119][3] +
                mat_A[75][3] * mat_B[127][3] +
                mat_A[76][0] * mat_B[135][3] +
                mat_A[76][1] * mat_B[143][3] +
                mat_A[76][2] * mat_B[151][3] +
                mat_A[76][3] * mat_B[159][3] +
                mat_A[77][0] * mat_B[167][3] +
                mat_A[77][1] * mat_B[175][3] +
                mat_A[77][2] * mat_B[183][3] +
                mat_A[77][3] * mat_B[191][3] +
                mat_A[78][0] * mat_B[199][3] +
                mat_A[78][1] * mat_B[207][3] +
                mat_A[78][2] * mat_B[215][3] +
                mat_A[78][3] * mat_B[223][3] +
                mat_A[79][0] * mat_B[231][3] +
                mat_A[79][1] * mat_B[239][3] +
                mat_A[79][2] * mat_B[247][3] +
                mat_A[79][3] * mat_B[255][3];
    mat_C[80][0] <=
                mat_A[80][0] * mat_B[0][0] +
                mat_A[80][1] * mat_B[8][0] +
                mat_A[80][2] * mat_B[16][0] +
                mat_A[80][3] * mat_B[24][0] +
                mat_A[81][0] * mat_B[32][0] +
                mat_A[81][1] * mat_B[40][0] +
                mat_A[81][2] * mat_B[48][0] +
                mat_A[81][3] * mat_B[56][0] +
                mat_A[82][0] * mat_B[64][0] +
                mat_A[82][1] * mat_B[72][0] +
                mat_A[82][2] * mat_B[80][0] +
                mat_A[82][3] * mat_B[88][0] +
                mat_A[83][0] * mat_B[96][0] +
                mat_A[83][1] * mat_B[104][0] +
                mat_A[83][2] * mat_B[112][0] +
                mat_A[83][3] * mat_B[120][0] +
                mat_A[84][0] * mat_B[128][0] +
                mat_A[84][1] * mat_B[136][0] +
                mat_A[84][2] * mat_B[144][0] +
                mat_A[84][3] * mat_B[152][0] +
                mat_A[85][0] * mat_B[160][0] +
                mat_A[85][1] * mat_B[168][0] +
                mat_A[85][2] * mat_B[176][0] +
                mat_A[85][3] * mat_B[184][0] +
                mat_A[86][0] * mat_B[192][0] +
                mat_A[86][1] * mat_B[200][0] +
                mat_A[86][2] * mat_B[208][0] +
                mat_A[86][3] * mat_B[216][0] +
                mat_A[87][0] * mat_B[224][0] +
                mat_A[87][1] * mat_B[232][0] +
                mat_A[87][2] * mat_B[240][0] +
                mat_A[87][3] * mat_B[248][0];
    mat_C[80][1] <=
                mat_A[80][0] * mat_B[0][1] +
                mat_A[80][1] * mat_B[8][1] +
                mat_A[80][2] * mat_B[16][1] +
                mat_A[80][3] * mat_B[24][1] +
                mat_A[81][0] * mat_B[32][1] +
                mat_A[81][1] * mat_B[40][1] +
                mat_A[81][2] * mat_B[48][1] +
                mat_A[81][3] * mat_B[56][1] +
                mat_A[82][0] * mat_B[64][1] +
                mat_A[82][1] * mat_B[72][1] +
                mat_A[82][2] * mat_B[80][1] +
                mat_A[82][3] * mat_B[88][1] +
                mat_A[83][0] * mat_B[96][1] +
                mat_A[83][1] * mat_B[104][1] +
                mat_A[83][2] * mat_B[112][1] +
                mat_A[83][3] * mat_B[120][1] +
                mat_A[84][0] * mat_B[128][1] +
                mat_A[84][1] * mat_B[136][1] +
                mat_A[84][2] * mat_B[144][1] +
                mat_A[84][3] * mat_B[152][1] +
                mat_A[85][0] * mat_B[160][1] +
                mat_A[85][1] * mat_B[168][1] +
                mat_A[85][2] * mat_B[176][1] +
                mat_A[85][3] * mat_B[184][1] +
                mat_A[86][0] * mat_B[192][1] +
                mat_A[86][1] * mat_B[200][1] +
                mat_A[86][2] * mat_B[208][1] +
                mat_A[86][3] * mat_B[216][1] +
                mat_A[87][0] * mat_B[224][1] +
                mat_A[87][1] * mat_B[232][1] +
                mat_A[87][2] * mat_B[240][1] +
                mat_A[87][3] * mat_B[248][1];
    mat_C[80][2] <=
                mat_A[80][0] * mat_B[0][2] +
                mat_A[80][1] * mat_B[8][2] +
                mat_A[80][2] * mat_B[16][2] +
                mat_A[80][3] * mat_B[24][2] +
                mat_A[81][0] * mat_B[32][2] +
                mat_A[81][1] * mat_B[40][2] +
                mat_A[81][2] * mat_B[48][2] +
                mat_A[81][3] * mat_B[56][2] +
                mat_A[82][0] * mat_B[64][2] +
                mat_A[82][1] * mat_B[72][2] +
                mat_A[82][2] * mat_B[80][2] +
                mat_A[82][3] * mat_B[88][2] +
                mat_A[83][0] * mat_B[96][2] +
                mat_A[83][1] * mat_B[104][2] +
                mat_A[83][2] * mat_B[112][2] +
                mat_A[83][3] * mat_B[120][2] +
                mat_A[84][0] * mat_B[128][2] +
                mat_A[84][1] * mat_B[136][2] +
                mat_A[84][2] * mat_B[144][2] +
                mat_A[84][3] * mat_B[152][2] +
                mat_A[85][0] * mat_B[160][2] +
                mat_A[85][1] * mat_B[168][2] +
                mat_A[85][2] * mat_B[176][2] +
                mat_A[85][3] * mat_B[184][2] +
                mat_A[86][0] * mat_B[192][2] +
                mat_A[86][1] * mat_B[200][2] +
                mat_A[86][2] * mat_B[208][2] +
                mat_A[86][3] * mat_B[216][2] +
                mat_A[87][0] * mat_B[224][2] +
                mat_A[87][1] * mat_B[232][2] +
                mat_A[87][2] * mat_B[240][2] +
                mat_A[87][3] * mat_B[248][2];
    mat_C[80][3] <=
                mat_A[80][0] * mat_B[0][3] +
                mat_A[80][1] * mat_B[8][3] +
                mat_A[80][2] * mat_B[16][3] +
                mat_A[80][3] * mat_B[24][3] +
                mat_A[81][0] * mat_B[32][3] +
                mat_A[81][1] * mat_B[40][3] +
                mat_A[81][2] * mat_B[48][3] +
                mat_A[81][3] * mat_B[56][3] +
                mat_A[82][0] * mat_B[64][3] +
                mat_A[82][1] * mat_B[72][3] +
                mat_A[82][2] * mat_B[80][3] +
                mat_A[82][3] * mat_B[88][3] +
                mat_A[83][0] * mat_B[96][3] +
                mat_A[83][1] * mat_B[104][3] +
                mat_A[83][2] * mat_B[112][3] +
                mat_A[83][3] * mat_B[120][3] +
                mat_A[84][0] * mat_B[128][3] +
                mat_A[84][1] * mat_B[136][3] +
                mat_A[84][2] * mat_B[144][3] +
                mat_A[84][3] * mat_B[152][3] +
                mat_A[85][0] * mat_B[160][3] +
                mat_A[85][1] * mat_B[168][3] +
                mat_A[85][2] * mat_B[176][3] +
                mat_A[85][3] * mat_B[184][3] +
                mat_A[86][0] * mat_B[192][3] +
                mat_A[86][1] * mat_B[200][3] +
                mat_A[86][2] * mat_B[208][3] +
                mat_A[86][3] * mat_B[216][3] +
                mat_A[87][0] * mat_B[224][3] +
                mat_A[87][1] * mat_B[232][3] +
                mat_A[87][2] * mat_B[240][3] +
                mat_A[87][3] * mat_B[248][3];
    mat_C[81][0] <=
                mat_A[80][0] * mat_B[1][0] +
                mat_A[80][1] * mat_B[9][0] +
                mat_A[80][2] * mat_B[17][0] +
                mat_A[80][3] * mat_B[25][0] +
                mat_A[81][0] * mat_B[33][0] +
                mat_A[81][1] * mat_B[41][0] +
                mat_A[81][2] * mat_B[49][0] +
                mat_A[81][3] * mat_B[57][0] +
                mat_A[82][0] * mat_B[65][0] +
                mat_A[82][1] * mat_B[73][0] +
                mat_A[82][2] * mat_B[81][0] +
                mat_A[82][3] * mat_B[89][0] +
                mat_A[83][0] * mat_B[97][0] +
                mat_A[83][1] * mat_B[105][0] +
                mat_A[83][2] * mat_B[113][0] +
                mat_A[83][3] * mat_B[121][0] +
                mat_A[84][0] * mat_B[129][0] +
                mat_A[84][1] * mat_B[137][0] +
                mat_A[84][2] * mat_B[145][0] +
                mat_A[84][3] * mat_B[153][0] +
                mat_A[85][0] * mat_B[161][0] +
                mat_A[85][1] * mat_B[169][0] +
                mat_A[85][2] * mat_B[177][0] +
                mat_A[85][3] * mat_B[185][0] +
                mat_A[86][0] * mat_B[193][0] +
                mat_A[86][1] * mat_B[201][0] +
                mat_A[86][2] * mat_B[209][0] +
                mat_A[86][3] * mat_B[217][0] +
                mat_A[87][0] * mat_B[225][0] +
                mat_A[87][1] * mat_B[233][0] +
                mat_A[87][2] * mat_B[241][0] +
                mat_A[87][3] * mat_B[249][0];
    mat_C[81][1] <=
                mat_A[80][0] * mat_B[1][1] +
                mat_A[80][1] * mat_B[9][1] +
                mat_A[80][2] * mat_B[17][1] +
                mat_A[80][3] * mat_B[25][1] +
                mat_A[81][0] * mat_B[33][1] +
                mat_A[81][1] * mat_B[41][1] +
                mat_A[81][2] * mat_B[49][1] +
                mat_A[81][3] * mat_B[57][1] +
                mat_A[82][0] * mat_B[65][1] +
                mat_A[82][1] * mat_B[73][1] +
                mat_A[82][2] * mat_B[81][1] +
                mat_A[82][3] * mat_B[89][1] +
                mat_A[83][0] * mat_B[97][1] +
                mat_A[83][1] * mat_B[105][1] +
                mat_A[83][2] * mat_B[113][1] +
                mat_A[83][3] * mat_B[121][1] +
                mat_A[84][0] * mat_B[129][1] +
                mat_A[84][1] * mat_B[137][1] +
                mat_A[84][2] * mat_B[145][1] +
                mat_A[84][3] * mat_B[153][1] +
                mat_A[85][0] * mat_B[161][1] +
                mat_A[85][1] * mat_B[169][1] +
                mat_A[85][2] * mat_B[177][1] +
                mat_A[85][3] * mat_B[185][1] +
                mat_A[86][0] * mat_B[193][1] +
                mat_A[86][1] * mat_B[201][1] +
                mat_A[86][2] * mat_B[209][1] +
                mat_A[86][3] * mat_B[217][1] +
                mat_A[87][0] * mat_B[225][1] +
                mat_A[87][1] * mat_B[233][1] +
                mat_A[87][2] * mat_B[241][1] +
                mat_A[87][3] * mat_B[249][1];
    mat_C[81][2] <=
                mat_A[80][0] * mat_B[1][2] +
                mat_A[80][1] * mat_B[9][2] +
                mat_A[80][2] * mat_B[17][2] +
                mat_A[80][3] * mat_B[25][2] +
                mat_A[81][0] * mat_B[33][2] +
                mat_A[81][1] * mat_B[41][2] +
                mat_A[81][2] * mat_B[49][2] +
                mat_A[81][3] * mat_B[57][2] +
                mat_A[82][0] * mat_B[65][2] +
                mat_A[82][1] * mat_B[73][2] +
                mat_A[82][2] * mat_B[81][2] +
                mat_A[82][3] * mat_B[89][2] +
                mat_A[83][0] * mat_B[97][2] +
                mat_A[83][1] * mat_B[105][2] +
                mat_A[83][2] * mat_B[113][2] +
                mat_A[83][3] * mat_B[121][2] +
                mat_A[84][0] * mat_B[129][2] +
                mat_A[84][1] * mat_B[137][2] +
                mat_A[84][2] * mat_B[145][2] +
                mat_A[84][3] * mat_B[153][2] +
                mat_A[85][0] * mat_B[161][2] +
                mat_A[85][1] * mat_B[169][2] +
                mat_A[85][2] * mat_B[177][2] +
                mat_A[85][3] * mat_B[185][2] +
                mat_A[86][0] * mat_B[193][2] +
                mat_A[86][1] * mat_B[201][2] +
                mat_A[86][2] * mat_B[209][2] +
                mat_A[86][3] * mat_B[217][2] +
                mat_A[87][0] * mat_B[225][2] +
                mat_A[87][1] * mat_B[233][2] +
                mat_A[87][2] * mat_B[241][2] +
                mat_A[87][3] * mat_B[249][2];
    mat_C[81][3] <=
                mat_A[80][0] * mat_B[1][3] +
                mat_A[80][1] * mat_B[9][3] +
                mat_A[80][2] * mat_B[17][3] +
                mat_A[80][3] * mat_B[25][3] +
                mat_A[81][0] * mat_B[33][3] +
                mat_A[81][1] * mat_B[41][3] +
                mat_A[81][2] * mat_B[49][3] +
                mat_A[81][3] * mat_B[57][3] +
                mat_A[82][0] * mat_B[65][3] +
                mat_A[82][1] * mat_B[73][3] +
                mat_A[82][2] * mat_B[81][3] +
                mat_A[82][3] * mat_B[89][3] +
                mat_A[83][0] * mat_B[97][3] +
                mat_A[83][1] * mat_B[105][3] +
                mat_A[83][2] * mat_B[113][3] +
                mat_A[83][3] * mat_B[121][3] +
                mat_A[84][0] * mat_B[129][3] +
                mat_A[84][1] * mat_B[137][3] +
                mat_A[84][2] * mat_B[145][3] +
                mat_A[84][3] * mat_B[153][3] +
                mat_A[85][0] * mat_B[161][3] +
                mat_A[85][1] * mat_B[169][3] +
                mat_A[85][2] * mat_B[177][3] +
                mat_A[85][3] * mat_B[185][3] +
                mat_A[86][0] * mat_B[193][3] +
                mat_A[86][1] * mat_B[201][3] +
                mat_A[86][2] * mat_B[209][3] +
                mat_A[86][3] * mat_B[217][3] +
                mat_A[87][0] * mat_B[225][3] +
                mat_A[87][1] * mat_B[233][3] +
                mat_A[87][2] * mat_B[241][3] +
                mat_A[87][3] * mat_B[249][3];
    mat_C[82][0] <=
                mat_A[80][0] * mat_B[2][0] +
                mat_A[80][1] * mat_B[10][0] +
                mat_A[80][2] * mat_B[18][0] +
                mat_A[80][3] * mat_B[26][0] +
                mat_A[81][0] * mat_B[34][0] +
                mat_A[81][1] * mat_B[42][0] +
                mat_A[81][2] * mat_B[50][0] +
                mat_A[81][3] * mat_B[58][0] +
                mat_A[82][0] * mat_B[66][0] +
                mat_A[82][1] * mat_B[74][0] +
                mat_A[82][2] * mat_B[82][0] +
                mat_A[82][3] * mat_B[90][0] +
                mat_A[83][0] * mat_B[98][0] +
                mat_A[83][1] * mat_B[106][0] +
                mat_A[83][2] * mat_B[114][0] +
                mat_A[83][3] * mat_B[122][0] +
                mat_A[84][0] * mat_B[130][0] +
                mat_A[84][1] * mat_B[138][0] +
                mat_A[84][2] * mat_B[146][0] +
                mat_A[84][3] * mat_B[154][0] +
                mat_A[85][0] * mat_B[162][0] +
                mat_A[85][1] * mat_B[170][0] +
                mat_A[85][2] * mat_B[178][0] +
                mat_A[85][3] * mat_B[186][0] +
                mat_A[86][0] * mat_B[194][0] +
                mat_A[86][1] * mat_B[202][0] +
                mat_A[86][2] * mat_B[210][0] +
                mat_A[86][3] * mat_B[218][0] +
                mat_A[87][0] * mat_B[226][0] +
                mat_A[87][1] * mat_B[234][0] +
                mat_A[87][2] * mat_B[242][0] +
                mat_A[87][3] * mat_B[250][0];
    mat_C[82][1] <=
                mat_A[80][0] * mat_B[2][1] +
                mat_A[80][1] * mat_B[10][1] +
                mat_A[80][2] * mat_B[18][1] +
                mat_A[80][3] * mat_B[26][1] +
                mat_A[81][0] * mat_B[34][1] +
                mat_A[81][1] * mat_B[42][1] +
                mat_A[81][2] * mat_B[50][1] +
                mat_A[81][3] * mat_B[58][1] +
                mat_A[82][0] * mat_B[66][1] +
                mat_A[82][1] * mat_B[74][1] +
                mat_A[82][2] * mat_B[82][1] +
                mat_A[82][3] * mat_B[90][1] +
                mat_A[83][0] * mat_B[98][1] +
                mat_A[83][1] * mat_B[106][1] +
                mat_A[83][2] * mat_B[114][1] +
                mat_A[83][3] * mat_B[122][1] +
                mat_A[84][0] * mat_B[130][1] +
                mat_A[84][1] * mat_B[138][1] +
                mat_A[84][2] * mat_B[146][1] +
                mat_A[84][3] * mat_B[154][1] +
                mat_A[85][0] * mat_B[162][1] +
                mat_A[85][1] * mat_B[170][1] +
                mat_A[85][2] * mat_B[178][1] +
                mat_A[85][3] * mat_B[186][1] +
                mat_A[86][0] * mat_B[194][1] +
                mat_A[86][1] * mat_B[202][1] +
                mat_A[86][2] * mat_B[210][1] +
                mat_A[86][3] * mat_B[218][1] +
                mat_A[87][0] * mat_B[226][1] +
                mat_A[87][1] * mat_B[234][1] +
                mat_A[87][2] * mat_B[242][1] +
                mat_A[87][3] * mat_B[250][1];
    mat_C[82][2] <=
                mat_A[80][0] * mat_B[2][2] +
                mat_A[80][1] * mat_B[10][2] +
                mat_A[80][2] * mat_B[18][2] +
                mat_A[80][3] * mat_B[26][2] +
                mat_A[81][0] * mat_B[34][2] +
                mat_A[81][1] * mat_B[42][2] +
                mat_A[81][2] * mat_B[50][2] +
                mat_A[81][3] * mat_B[58][2] +
                mat_A[82][0] * mat_B[66][2] +
                mat_A[82][1] * mat_B[74][2] +
                mat_A[82][2] * mat_B[82][2] +
                mat_A[82][3] * mat_B[90][2] +
                mat_A[83][0] * mat_B[98][2] +
                mat_A[83][1] * mat_B[106][2] +
                mat_A[83][2] * mat_B[114][2] +
                mat_A[83][3] * mat_B[122][2] +
                mat_A[84][0] * mat_B[130][2] +
                mat_A[84][1] * mat_B[138][2] +
                mat_A[84][2] * mat_B[146][2] +
                mat_A[84][3] * mat_B[154][2] +
                mat_A[85][0] * mat_B[162][2] +
                mat_A[85][1] * mat_B[170][2] +
                mat_A[85][2] * mat_B[178][2] +
                mat_A[85][3] * mat_B[186][2] +
                mat_A[86][0] * mat_B[194][2] +
                mat_A[86][1] * mat_B[202][2] +
                mat_A[86][2] * mat_B[210][2] +
                mat_A[86][3] * mat_B[218][2] +
                mat_A[87][0] * mat_B[226][2] +
                mat_A[87][1] * mat_B[234][2] +
                mat_A[87][2] * mat_B[242][2] +
                mat_A[87][3] * mat_B[250][2];
    mat_C[82][3] <=
                mat_A[80][0] * mat_B[2][3] +
                mat_A[80][1] * mat_B[10][3] +
                mat_A[80][2] * mat_B[18][3] +
                mat_A[80][3] * mat_B[26][3] +
                mat_A[81][0] * mat_B[34][3] +
                mat_A[81][1] * mat_B[42][3] +
                mat_A[81][2] * mat_B[50][3] +
                mat_A[81][3] * mat_B[58][3] +
                mat_A[82][0] * mat_B[66][3] +
                mat_A[82][1] * mat_B[74][3] +
                mat_A[82][2] * mat_B[82][3] +
                mat_A[82][3] * mat_B[90][3] +
                mat_A[83][0] * mat_B[98][3] +
                mat_A[83][1] * mat_B[106][3] +
                mat_A[83][2] * mat_B[114][3] +
                mat_A[83][3] * mat_B[122][3] +
                mat_A[84][0] * mat_B[130][3] +
                mat_A[84][1] * mat_B[138][3] +
                mat_A[84][2] * mat_B[146][3] +
                mat_A[84][3] * mat_B[154][3] +
                mat_A[85][0] * mat_B[162][3] +
                mat_A[85][1] * mat_B[170][3] +
                mat_A[85][2] * mat_B[178][3] +
                mat_A[85][3] * mat_B[186][3] +
                mat_A[86][0] * mat_B[194][3] +
                mat_A[86][1] * mat_B[202][3] +
                mat_A[86][2] * mat_B[210][3] +
                mat_A[86][3] * mat_B[218][3] +
                mat_A[87][0] * mat_B[226][3] +
                mat_A[87][1] * mat_B[234][3] +
                mat_A[87][2] * mat_B[242][3] +
                mat_A[87][3] * mat_B[250][3];
    mat_C[83][0] <=
                mat_A[80][0] * mat_B[3][0] +
                mat_A[80][1] * mat_B[11][0] +
                mat_A[80][2] * mat_B[19][0] +
                mat_A[80][3] * mat_B[27][0] +
                mat_A[81][0] * mat_B[35][0] +
                mat_A[81][1] * mat_B[43][0] +
                mat_A[81][2] * mat_B[51][0] +
                mat_A[81][3] * mat_B[59][0] +
                mat_A[82][0] * mat_B[67][0] +
                mat_A[82][1] * mat_B[75][0] +
                mat_A[82][2] * mat_B[83][0] +
                mat_A[82][3] * mat_B[91][0] +
                mat_A[83][0] * mat_B[99][0] +
                mat_A[83][1] * mat_B[107][0] +
                mat_A[83][2] * mat_B[115][0] +
                mat_A[83][3] * mat_B[123][0] +
                mat_A[84][0] * mat_B[131][0] +
                mat_A[84][1] * mat_B[139][0] +
                mat_A[84][2] * mat_B[147][0] +
                mat_A[84][3] * mat_B[155][0] +
                mat_A[85][0] * mat_B[163][0] +
                mat_A[85][1] * mat_B[171][0] +
                mat_A[85][2] * mat_B[179][0] +
                mat_A[85][3] * mat_B[187][0] +
                mat_A[86][0] * mat_B[195][0] +
                mat_A[86][1] * mat_B[203][0] +
                mat_A[86][2] * mat_B[211][0] +
                mat_A[86][3] * mat_B[219][0] +
                mat_A[87][0] * mat_B[227][0] +
                mat_A[87][1] * mat_B[235][0] +
                mat_A[87][2] * mat_B[243][0] +
                mat_A[87][3] * mat_B[251][0];
    mat_C[83][1] <=
                mat_A[80][0] * mat_B[3][1] +
                mat_A[80][1] * mat_B[11][1] +
                mat_A[80][2] * mat_B[19][1] +
                mat_A[80][3] * mat_B[27][1] +
                mat_A[81][0] * mat_B[35][1] +
                mat_A[81][1] * mat_B[43][1] +
                mat_A[81][2] * mat_B[51][1] +
                mat_A[81][3] * mat_B[59][1] +
                mat_A[82][0] * mat_B[67][1] +
                mat_A[82][1] * mat_B[75][1] +
                mat_A[82][2] * mat_B[83][1] +
                mat_A[82][3] * mat_B[91][1] +
                mat_A[83][0] * mat_B[99][1] +
                mat_A[83][1] * mat_B[107][1] +
                mat_A[83][2] * mat_B[115][1] +
                mat_A[83][3] * mat_B[123][1] +
                mat_A[84][0] * mat_B[131][1] +
                mat_A[84][1] * mat_B[139][1] +
                mat_A[84][2] * mat_B[147][1] +
                mat_A[84][3] * mat_B[155][1] +
                mat_A[85][0] * mat_B[163][1] +
                mat_A[85][1] * mat_B[171][1] +
                mat_A[85][2] * mat_B[179][1] +
                mat_A[85][3] * mat_B[187][1] +
                mat_A[86][0] * mat_B[195][1] +
                mat_A[86][1] * mat_B[203][1] +
                mat_A[86][2] * mat_B[211][1] +
                mat_A[86][3] * mat_B[219][1] +
                mat_A[87][0] * mat_B[227][1] +
                mat_A[87][1] * mat_B[235][1] +
                mat_A[87][2] * mat_B[243][1] +
                mat_A[87][3] * mat_B[251][1];
    mat_C[83][2] <=
                mat_A[80][0] * mat_B[3][2] +
                mat_A[80][1] * mat_B[11][2] +
                mat_A[80][2] * mat_B[19][2] +
                mat_A[80][3] * mat_B[27][2] +
                mat_A[81][0] * mat_B[35][2] +
                mat_A[81][1] * mat_B[43][2] +
                mat_A[81][2] * mat_B[51][2] +
                mat_A[81][3] * mat_B[59][2] +
                mat_A[82][0] * mat_B[67][2] +
                mat_A[82][1] * mat_B[75][2] +
                mat_A[82][2] * mat_B[83][2] +
                mat_A[82][3] * mat_B[91][2] +
                mat_A[83][0] * mat_B[99][2] +
                mat_A[83][1] * mat_B[107][2] +
                mat_A[83][2] * mat_B[115][2] +
                mat_A[83][3] * mat_B[123][2] +
                mat_A[84][0] * mat_B[131][2] +
                mat_A[84][1] * mat_B[139][2] +
                mat_A[84][2] * mat_B[147][2] +
                mat_A[84][3] * mat_B[155][2] +
                mat_A[85][0] * mat_B[163][2] +
                mat_A[85][1] * mat_B[171][2] +
                mat_A[85][2] * mat_B[179][2] +
                mat_A[85][3] * mat_B[187][2] +
                mat_A[86][0] * mat_B[195][2] +
                mat_A[86][1] * mat_B[203][2] +
                mat_A[86][2] * mat_B[211][2] +
                mat_A[86][3] * mat_B[219][2] +
                mat_A[87][0] * mat_B[227][2] +
                mat_A[87][1] * mat_B[235][2] +
                mat_A[87][2] * mat_B[243][2] +
                mat_A[87][3] * mat_B[251][2];
    mat_C[83][3] <=
                mat_A[80][0] * mat_B[3][3] +
                mat_A[80][1] * mat_B[11][3] +
                mat_A[80][2] * mat_B[19][3] +
                mat_A[80][3] * mat_B[27][3] +
                mat_A[81][0] * mat_B[35][3] +
                mat_A[81][1] * mat_B[43][3] +
                mat_A[81][2] * mat_B[51][3] +
                mat_A[81][3] * mat_B[59][3] +
                mat_A[82][0] * mat_B[67][3] +
                mat_A[82][1] * mat_B[75][3] +
                mat_A[82][2] * mat_B[83][3] +
                mat_A[82][3] * mat_B[91][3] +
                mat_A[83][0] * mat_B[99][3] +
                mat_A[83][1] * mat_B[107][3] +
                mat_A[83][2] * mat_B[115][3] +
                mat_A[83][3] * mat_B[123][3] +
                mat_A[84][0] * mat_B[131][3] +
                mat_A[84][1] * mat_B[139][3] +
                mat_A[84][2] * mat_B[147][3] +
                mat_A[84][3] * mat_B[155][3] +
                mat_A[85][0] * mat_B[163][3] +
                mat_A[85][1] * mat_B[171][3] +
                mat_A[85][2] * mat_B[179][3] +
                mat_A[85][3] * mat_B[187][3] +
                mat_A[86][0] * mat_B[195][3] +
                mat_A[86][1] * mat_B[203][3] +
                mat_A[86][2] * mat_B[211][3] +
                mat_A[86][3] * mat_B[219][3] +
                mat_A[87][0] * mat_B[227][3] +
                mat_A[87][1] * mat_B[235][3] +
                mat_A[87][2] * mat_B[243][3] +
                mat_A[87][3] * mat_B[251][3];
    mat_C[84][0] <=
                mat_A[80][0] * mat_B[4][0] +
                mat_A[80][1] * mat_B[12][0] +
                mat_A[80][2] * mat_B[20][0] +
                mat_A[80][3] * mat_B[28][0] +
                mat_A[81][0] * mat_B[36][0] +
                mat_A[81][1] * mat_B[44][0] +
                mat_A[81][2] * mat_B[52][0] +
                mat_A[81][3] * mat_B[60][0] +
                mat_A[82][0] * mat_B[68][0] +
                mat_A[82][1] * mat_B[76][0] +
                mat_A[82][2] * mat_B[84][0] +
                mat_A[82][3] * mat_B[92][0] +
                mat_A[83][0] * mat_B[100][0] +
                mat_A[83][1] * mat_B[108][0] +
                mat_A[83][2] * mat_B[116][0] +
                mat_A[83][3] * mat_B[124][0] +
                mat_A[84][0] * mat_B[132][0] +
                mat_A[84][1] * mat_B[140][0] +
                mat_A[84][2] * mat_B[148][0] +
                mat_A[84][3] * mat_B[156][0] +
                mat_A[85][0] * mat_B[164][0] +
                mat_A[85][1] * mat_B[172][0] +
                mat_A[85][2] * mat_B[180][0] +
                mat_A[85][3] * mat_B[188][0] +
                mat_A[86][0] * mat_B[196][0] +
                mat_A[86][1] * mat_B[204][0] +
                mat_A[86][2] * mat_B[212][0] +
                mat_A[86][3] * mat_B[220][0] +
                mat_A[87][0] * mat_B[228][0] +
                mat_A[87][1] * mat_B[236][0] +
                mat_A[87][2] * mat_B[244][0] +
                mat_A[87][3] * mat_B[252][0];
    mat_C[84][1] <=
                mat_A[80][0] * mat_B[4][1] +
                mat_A[80][1] * mat_B[12][1] +
                mat_A[80][2] * mat_B[20][1] +
                mat_A[80][3] * mat_B[28][1] +
                mat_A[81][0] * mat_B[36][1] +
                mat_A[81][1] * mat_B[44][1] +
                mat_A[81][2] * mat_B[52][1] +
                mat_A[81][3] * mat_B[60][1] +
                mat_A[82][0] * mat_B[68][1] +
                mat_A[82][1] * mat_B[76][1] +
                mat_A[82][2] * mat_B[84][1] +
                mat_A[82][3] * mat_B[92][1] +
                mat_A[83][0] * mat_B[100][1] +
                mat_A[83][1] * mat_B[108][1] +
                mat_A[83][2] * mat_B[116][1] +
                mat_A[83][3] * mat_B[124][1] +
                mat_A[84][0] * mat_B[132][1] +
                mat_A[84][1] * mat_B[140][1] +
                mat_A[84][2] * mat_B[148][1] +
                mat_A[84][3] * mat_B[156][1] +
                mat_A[85][0] * mat_B[164][1] +
                mat_A[85][1] * mat_B[172][1] +
                mat_A[85][2] * mat_B[180][1] +
                mat_A[85][3] * mat_B[188][1] +
                mat_A[86][0] * mat_B[196][1] +
                mat_A[86][1] * mat_B[204][1] +
                mat_A[86][2] * mat_B[212][1] +
                mat_A[86][3] * mat_B[220][1] +
                mat_A[87][0] * mat_B[228][1] +
                mat_A[87][1] * mat_B[236][1] +
                mat_A[87][2] * mat_B[244][1] +
                mat_A[87][3] * mat_B[252][1];
    mat_C[84][2] <=
                mat_A[80][0] * mat_B[4][2] +
                mat_A[80][1] * mat_B[12][2] +
                mat_A[80][2] * mat_B[20][2] +
                mat_A[80][3] * mat_B[28][2] +
                mat_A[81][0] * mat_B[36][2] +
                mat_A[81][1] * mat_B[44][2] +
                mat_A[81][2] * mat_B[52][2] +
                mat_A[81][3] * mat_B[60][2] +
                mat_A[82][0] * mat_B[68][2] +
                mat_A[82][1] * mat_B[76][2] +
                mat_A[82][2] * mat_B[84][2] +
                mat_A[82][3] * mat_B[92][2] +
                mat_A[83][0] * mat_B[100][2] +
                mat_A[83][1] * mat_B[108][2] +
                mat_A[83][2] * mat_B[116][2] +
                mat_A[83][3] * mat_B[124][2] +
                mat_A[84][0] * mat_B[132][2] +
                mat_A[84][1] * mat_B[140][2] +
                mat_A[84][2] * mat_B[148][2] +
                mat_A[84][3] * mat_B[156][2] +
                mat_A[85][0] * mat_B[164][2] +
                mat_A[85][1] * mat_B[172][2] +
                mat_A[85][2] * mat_B[180][2] +
                mat_A[85][3] * mat_B[188][2] +
                mat_A[86][0] * mat_B[196][2] +
                mat_A[86][1] * mat_B[204][2] +
                mat_A[86][2] * mat_B[212][2] +
                mat_A[86][3] * mat_B[220][2] +
                mat_A[87][0] * mat_B[228][2] +
                mat_A[87][1] * mat_B[236][2] +
                mat_A[87][2] * mat_B[244][2] +
                mat_A[87][3] * mat_B[252][2];
    mat_C[84][3] <=
                mat_A[80][0] * mat_B[4][3] +
                mat_A[80][1] * mat_B[12][3] +
                mat_A[80][2] * mat_B[20][3] +
                mat_A[80][3] * mat_B[28][3] +
                mat_A[81][0] * mat_B[36][3] +
                mat_A[81][1] * mat_B[44][3] +
                mat_A[81][2] * mat_B[52][3] +
                mat_A[81][3] * mat_B[60][3] +
                mat_A[82][0] * mat_B[68][3] +
                mat_A[82][1] * mat_B[76][3] +
                mat_A[82][2] * mat_B[84][3] +
                mat_A[82][3] * mat_B[92][3] +
                mat_A[83][0] * mat_B[100][3] +
                mat_A[83][1] * mat_B[108][3] +
                mat_A[83][2] * mat_B[116][3] +
                mat_A[83][3] * mat_B[124][3] +
                mat_A[84][0] * mat_B[132][3] +
                mat_A[84][1] * mat_B[140][3] +
                mat_A[84][2] * mat_B[148][3] +
                mat_A[84][3] * mat_B[156][3] +
                mat_A[85][0] * mat_B[164][3] +
                mat_A[85][1] * mat_B[172][3] +
                mat_A[85][2] * mat_B[180][3] +
                mat_A[85][3] * mat_B[188][3] +
                mat_A[86][0] * mat_B[196][3] +
                mat_A[86][1] * mat_B[204][3] +
                mat_A[86][2] * mat_B[212][3] +
                mat_A[86][3] * mat_B[220][3] +
                mat_A[87][0] * mat_B[228][3] +
                mat_A[87][1] * mat_B[236][3] +
                mat_A[87][2] * mat_B[244][3] +
                mat_A[87][3] * mat_B[252][3];
    mat_C[85][0] <=
                mat_A[80][0] * mat_B[5][0] +
                mat_A[80][1] * mat_B[13][0] +
                mat_A[80][2] * mat_B[21][0] +
                mat_A[80][3] * mat_B[29][0] +
                mat_A[81][0] * mat_B[37][0] +
                mat_A[81][1] * mat_B[45][0] +
                mat_A[81][2] * mat_B[53][0] +
                mat_A[81][3] * mat_B[61][0] +
                mat_A[82][0] * mat_B[69][0] +
                mat_A[82][1] * mat_B[77][0] +
                mat_A[82][2] * mat_B[85][0] +
                mat_A[82][3] * mat_B[93][0] +
                mat_A[83][0] * mat_B[101][0] +
                mat_A[83][1] * mat_B[109][0] +
                mat_A[83][2] * mat_B[117][0] +
                mat_A[83][3] * mat_B[125][0] +
                mat_A[84][0] * mat_B[133][0] +
                mat_A[84][1] * mat_B[141][0] +
                mat_A[84][2] * mat_B[149][0] +
                mat_A[84][3] * mat_B[157][0] +
                mat_A[85][0] * mat_B[165][0] +
                mat_A[85][1] * mat_B[173][0] +
                mat_A[85][2] * mat_B[181][0] +
                mat_A[85][3] * mat_B[189][0] +
                mat_A[86][0] * mat_B[197][0] +
                mat_A[86][1] * mat_B[205][0] +
                mat_A[86][2] * mat_B[213][0] +
                mat_A[86][3] * mat_B[221][0] +
                mat_A[87][0] * mat_B[229][0] +
                mat_A[87][1] * mat_B[237][0] +
                mat_A[87][2] * mat_B[245][0] +
                mat_A[87][3] * mat_B[253][0];
    mat_C[85][1] <=
                mat_A[80][0] * mat_B[5][1] +
                mat_A[80][1] * mat_B[13][1] +
                mat_A[80][2] * mat_B[21][1] +
                mat_A[80][3] * mat_B[29][1] +
                mat_A[81][0] * mat_B[37][1] +
                mat_A[81][1] * mat_B[45][1] +
                mat_A[81][2] * mat_B[53][1] +
                mat_A[81][3] * mat_B[61][1] +
                mat_A[82][0] * mat_B[69][1] +
                mat_A[82][1] * mat_B[77][1] +
                mat_A[82][2] * mat_B[85][1] +
                mat_A[82][3] * mat_B[93][1] +
                mat_A[83][0] * mat_B[101][1] +
                mat_A[83][1] * mat_B[109][1] +
                mat_A[83][2] * mat_B[117][1] +
                mat_A[83][3] * mat_B[125][1] +
                mat_A[84][0] * mat_B[133][1] +
                mat_A[84][1] * mat_B[141][1] +
                mat_A[84][2] * mat_B[149][1] +
                mat_A[84][3] * mat_B[157][1] +
                mat_A[85][0] * mat_B[165][1] +
                mat_A[85][1] * mat_B[173][1] +
                mat_A[85][2] * mat_B[181][1] +
                mat_A[85][3] * mat_B[189][1] +
                mat_A[86][0] * mat_B[197][1] +
                mat_A[86][1] * mat_B[205][1] +
                mat_A[86][2] * mat_B[213][1] +
                mat_A[86][3] * mat_B[221][1] +
                mat_A[87][0] * mat_B[229][1] +
                mat_A[87][1] * mat_B[237][1] +
                mat_A[87][2] * mat_B[245][1] +
                mat_A[87][3] * mat_B[253][1];
    mat_C[85][2] <=
                mat_A[80][0] * mat_B[5][2] +
                mat_A[80][1] * mat_B[13][2] +
                mat_A[80][2] * mat_B[21][2] +
                mat_A[80][3] * mat_B[29][2] +
                mat_A[81][0] * mat_B[37][2] +
                mat_A[81][1] * mat_B[45][2] +
                mat_A[81][2] * mat_B[53][2] +
                mat_A[81][3] * mat_B[61][2] +
                mat_A[82][0] * mat_B[69][2] +
                mat_A[82][1] * mat_B[77][2] +
                mat_A[82][2] * mat_B[85][2] +
                mat_A[82][3] * mat_B[93][2] +
                mat_A[83][0] * mat_B[101][2] +
                mat_A[83][1] * mat_B[109][2] +
                mat_A[83][2] * mat_B[117][2] +
                mat_A[83][3] * mat_B[125][2] +
                mat_A[84][0] * mat_B[133][2] +
                mat_A[84][1] * mat_B[141][2] +
                mat_A[84][2] * mat_B[149][2] +
                mat_A[84][3] * mat_B[157][2] +
                mat_A[85][0] * mat_B[165][2] +
                mat_A[85][1] * mat_B[173][2] +
                mat_A[85][2] * mat_B[181][2] +
                mat_A[85][3] * mat_B[189][2] +
                mat_A[86][0] * mat_B[197][2] +
                mat_A[86][1] * mat_B[205][2] +
                mat_A[86][2] * mat_B[213][2] +
                mat_A[86][3] * mat_B[221][2] +
                mat_A[87][0] * mat_B[229][2] +
                mat_A[87][1] * mat_B[237][2] +
                mat_A[87][2] * mat_B[245][2] +
                mat_A[87][3] * mat_B[253][2];
    mat_C[85][3] <=
                mat_A[80][0] * mat_B[5][3] +
                mat_A[80][1] * mat_B[13][3] +
                mat_A[80][2] * mat_B[21][3] +
                mat_A[80][3] * mat_B[29][3] +
                mat_A[81][0] * mat_B[37][3] +
                mat_A[81][1] * mat_B[45][3] +
                mat_A[81][2] * mat_B[53][3] +
                mat_A[81][3] * mat_B[61][3] +
                mat_A[82][0] * mat_B[69][3] +
                mat_A[82][1] * mat_B[77][3] +
                mat_A[82][2] * mat_B[85][3] +
                mat_A[82][3] * mat_B[93][3] +
                mat_A[83][0] * mat_B[101][3] +
                mat_A[83][1] * mat_B[109][3] +
                mat_A[83][2] * mat_B[117][3] +
                mat_A[83][3] * mat_B[125][3] +
                mat_A[84][0] * mat_B[133][3] +
                mat_A[84][1] * mat_B[141][3] +
                mat_A[84][2] * mat_B[149][3] +
                mat_A[84][3] * mat_B[157][3] +
                mat_A[85][0] * mat_B[165][3] +
                mat_A[85][1] * mat_B[173][3] +
                mat_A[85][2] * mat_B[181][3] +
                mat_A[85][3] * mat_B[189][3] +
                mat_A[86][0] * mat_B[197][3] +
                mat_A[86][1] * mat_B[205][3] +
                mat_A[86][2] * mat_B[213][3] +
                mat_A[86][3] * mat_B[221][3] +
                mat_A[87][0] * mat_B[229][3] +
                mat_A[87][1] * mat_B[237][3] +
                mat_A[87][2] * mat_B[245][3] +
                mat_A[87][3] * mat_B[253][3];
    mat_C[86][0] <=
                mat_A[80][0] * mat_B[6][0] +
                mat_A[80][1] * mat_B[14][0] +
                mat_A[80][2] * mat_B[22][0] +
                mat_A[80][3] * mat_B[30][0] +
                mat_A[81][0] * mat_B[38][0] +
                mat_A[81][1] * mat_B[46][0] +
                mat_A[81][2] * mat_B[54][0] +
                mat_A[81][3] * mat_B[62][0] +
                mat_A[82][0] * mat_B[70][0] +
                mat_A[82][1] * mat_B[78][0] +
                mat_A[82][2] * mat_B[86][0] +
                mat_A[82][3] * mat_B[94][0] +
                mat_A[83][0] * mat_B[102][0] +
                mat_A[83][1] * mat_B[110][0] +
                mat_A[83][2] * mat_B[118][0] +
                mat_A[83][3] * mat_B[126][0] +
                mat_A[84][0] * mat_B[134][0] +
                mat_A[84][1] * mat_B[142][0] +
                mat_A[84][2] * mat_B[150][0] +
                mat_A[84][3] * mat_B[158][0] +
                mat_A[85][0] * mat_B[166][0] +
                mat_A[85][1] * mat_B[174][0] +
                mat_A[85][2] * mat_B[182][0] +
                mat_A[85][3] * mat_B[190][0] +
                mat_A[86][0] * mat_B[198][0] +
                mat_A[86][1] * mat_B[206][0] +
                mat_A[86][2] * mat_B[214][0] +
                mat_A[86][3] * mat_B[222][0] +
                mat_A[87][0] * mat_B[230][0] +
                mat_A[87][1] * mat_B[238][0] +
                mat_A[87][2] * mat_B[246][0] +
                mat_A[87][3] * mat_B[254][0];
    mat_C[86][1] <=
                mat_A[80][0] * mat_B[6][1] +
                mat_A[80][1] * mat_B[14][1] +
                mat_A[80][2] * mat_B[22][1] +
                mat_A[80][3] * mat_B[30][1] +
                mat_A[81][0] * mat_B[38][1] +
                mat_A[81][1] * mat_B[46][1] +
                mat_A[81][2] * mat_B[54][1] +
                mat_A[81][3] * mat_B[62][1] +
                mat_A[82][0] * mat_B[70][1] +
                mat_A[82][1] * mat_B[78][1] +
                mat_A[82][2] * mat_B[86][1] +
                mat_A[82][3] * mat_B[94][1] +
                mat_A[83][0] * mat_B[102][1] +
                mat_A[83][1] * mat_B[110][1] +
                mat_A[83][2] * mat_B[118][1] +
                mat_A[83][3] * mat_B[126][1] +
                mat_A[84][0] * mat_B[134][1] +
                mat_A[84][1] * mat_B[142][1] +
                mat_A[84][2] * mat_B[150][1] +
                mat_A[84][3] * mat_B[158][1] +
                mat_A[85][0] * mat_B[166][1] +
                mat_A[85][1] * mat_B[174][1] +
                mat_A[85][2] * mat_B[182][1] +
                mat_A[85][3] * mat_B[190][1] +
                mat_A[86][0] * mat_B[198][1] +
                mat_A[86][1] * mat_B[206][1] +
                mat_A[86][2] * mat_B[214][1] +
                mat_A[86][3] * mat_B[222][1] +
                mat_A[87][0] * mat_B[230][1] +
                mat_A[87][1] * mat_B[238][1] +
                mat_A[87][2] * mat_B[246][1] +
                mat_A[87][3] * mat_B[254][1];
    mat_C[86][2] <=
                mat_A[80][0] * mat_B[6][2] +
                mat_A[80][1] * mat_B[14][2] +
                mat_A[80][2] * mat_B[22][2] +
                mat_A[80][3] * mat_B[30][2] +
                mat_A[81][0] * mat_B[38][2] +
                mat_A[81][1] * mat_B[46][2] +
                mat_A[81][2] * mat_B[54][2] +
                mat_A[81][3] * mat_B[62][2] +
                mat_A[82][0] * mat_B[70][2] +
                mat_A[82][1] * mat_B[78][2] +
                mat_A[82][2] * mat_B[86][2] +
                mat_A[82][3] * mat_B[94][2] +
                mat_A[83][0] * mat_B[102][2] +
                mat_A[83][1] * mat_B[110][2] +
                mat_A[83][2] * mat_B[118][2] +
                mat_A[83][3] * mat_B[126][2] +
                mat_A[84][0] * mat_B[134][2] +
                mat_A[84][1] * mat_B[142][2] +
                mat_A[84][2] * mat_B[150][2] +
                mat_A[84][3] * mat_B[158][2] +
                mat_A[85][0] * mat_B[166][2] +
                mat_A[85][1] * mat_B[174][2] +
                mat_A[85][2] * mat_B[182][2] +
                mat_A[85][3] * mat_B[190][2] +
                mat_A[86][0] * mat_B[198][2] +
                mat_A[86][1] * mat_B[206][2] +
                mat_A[86][2] * mat_B[214][2] +
                mat_A[86][3] * mat_B[222][2] +
                mat_A[87][0] * mat_B[230][2] +
                mat_A[87][1] * mat_B[238][2] +
                mat_A[87][2] * mat_B[246][2] +
                mat_A[87][3] * mat_B[254][2];
    mat_C[86][3] <=
                mat_A[80][0] * mat_B[6][3] +
                mat_A[80][1] * mat_B[14][3] +
                mat_A[80][2] * mat_B[22][3] +
                mat_A[80][3] * mat_B[30][3] +
                mat_A[81][0] * mat_B[38][3] +
                mat_A[81][1] * mat_B[46][3] +
                mat_A[81][2] * mat_B[54][3] +
                mat_A[81][3] * mat_B[62][3] +
                mat_A[82][0] * mat_B[70][3] +
                mat_A[82][1] * mat_B[78][3] +
                mat_A[82][2] * mat_B[86][3] +
                mat_A[82][3] * mat_B[94][3] +
                mat_A[83][0] * mat_B[102][3] +
                mat_A[83][1] * mat_B[110][3] +
                mat_A[83][2] * mat_B[118][3] +
                mat_A[83][3] * mat_B[126][3] +
                mat_A[84][0] * mat_B[134][3] +
                mat_A[84][1] * mat_B[142][3] +
                mat_A[84][2] * mat_B[150][3] +
                mat_A[84][3] * mat_B[158][3] +
                mat_A[85][0] * mat_B[166][3] +
                mat_A[85][1] * mat_B[174][3] +
                mat_A[85][2] * mat_B[182][3] +
                mat_A[85][3] * mat_B[190][3] +
                mat_A[86][0] * mat_B[198][3] +
                mat_A[86][1] * mat_B[206][3] +
                mat_A[86][2] * mat_B[214][3] +
                mat_A[86][3] * mat_B[222][3] +
                mat_A[87][0] * mat_B[230][3] +
                mat_A[87][1] * mat_B[238][3] +
                mat_A[87][2] * mat_B[246][3] +
                mat_A[87][3] * mat_B[254][3];
    mat_C[87][0] <=
                mat_A[80][0] * mat_B[7][0] +
                mat_A[80][1] * mat_B[15][0] +
                mat_A[80][2] * mat_B[23][0] +
                mat_A[80][3] * mat_B[31][0] +
                mat_A[81][0] * mat_B[39][0] +
                mat_A[81][1] * mat_B[47][0] +
                mat_A[81][2] * mat_B[55][0] +
                mat_A[81][3] * mat_B[63][0] +
                mat_A[82][0] * mat_B[71][0] +
                mat_A[82][1] * mat_B[79][0] +
                mat_A[82][2] * mat_B[87][0] +
                mat_A[82][3] * mat_B[95][0] +
                mat_A[83][0] * mat_B[103][0] +
                mat_A[83][1] * mat_B[111][0] +
                mat_A[83][2] * mat_B[119][0] +
                mat_A[83][3] * mat_B[127][0] +
                mat_A[84][0] * mat_B[135][0] +
                mat_A[84][1] * mat_B[143][0] +
                mat_A[84][2] * mat_B[151][0] +
                mat_A[84][3] * mat_B[159][0] +
                mat_A[85][0] * mat_B[167][0] +
                mat_A[85][1] * mat_B[175][0] +
                mat_A[85][2] * mat_B[183][0] +
                mat_A[85][3] * mat_B[191][0] +
                mat_A[86][0] * mat_B[199][0] +
                mat_A[86][1] * mat_B[207][0] +
                mat_A[86][2] * mat_B[215][0] +
                mat_A[86][3] * mat_B[223][0] +
                mat_A[87][0] * mat_B[231][0] +
                mat_A[87][1] * mat_B[239][0] +
                mat_A[87][2] * mat_B[247][0] +
                mat_A[87][3] * mat_B[255][0];
    mat_C[87][1] <=
                mat_A[80][0] * mat_B[7][1] +
                mat_A[80][1] * mat_B[15][1] +
                mat_A[80][2] * mat_B[23][1] +
                mat_A[80][3] * mat_B[31][1] +
                mat_A[81][0] * mat_B[39][1] +
                mat_A[81][1] * mat_B[47][1] +
                mat_A[81][2] * mat_B[55][1] +
                mat_A[81][3] * mat_B[63][1] +
                mat_A[82][0] * mat_B[71][1] +
                mat_A[82][1] * mat_B[79][1] +
                mat_A[82][2] * mat_B[87][1] +
                mat_A[82][3] * mat_B[95][1] +
                mat_A[83][0] * mat_B[103][1] +
                mat_A[83][1] * mat_B[111][1] +
                mat_A[83][2] * mat_B[119][1] +
                mat_A[83][3] * mat_B[127][1] +
                mat_A[84][0] * mat_B[135][1] +
                mat_A[84][1] * mat_B[143][1] +
                mat_A[84][2] * mat_B[151][1] +
                mat_A[84][3] * mat_B[159][1] +
                mat_A[85][0] * mat_B[167][1] +
                mat_A[85][1] * mat_B[175][1] +
                mat_A[85][2] * mat_B[183][1] +
                mat_A[85][3] * mat_B[191][1] +
                mat_A[86][0] * mat_B[199][1] +
                mat_A[86][1] * mat_B[207][1] +
                mat_A[86][2] * mat_B[215][1] +
                mat_A[86][3] * mat_B[223][1] +
                mat_A[87][0] * mat_B[231][1] +
                mat_A[87][1] * mat_B[239][1] +
                mat_A[87][2] * mat_B[247][1] +
                mat_A[87][3] * mat_B[255][1];
    mat_C[87][2] <=
                mat_A[80][0] * mat_B[7][2] +
                mat_A[80][1] * mat_B[15][2] +
                mat_A[80][2] * mat_B[23][2] +
                mat_A[80][3] * mat_B[31][2] +
                mat_A[81][0] * mat_B[39][2] +
                mat_A[81][1] * mat_B[47][2] +
                mat_A[81][2] * mat_B[55][2] +
                mat_A[81][3] * mat_B[63][2] +
                mat_A[82][0] * mat_B[71][2] +
                mat_A[82][1] * mat_B[79][2] +
                mat_A[82][2] * mat_B[87][2] +
                mat_A[82][3] * mat_B[95][2] +
                mat_A[83][0] * mat_B[103][2] +
                mat_A[83][1] * mat_B[111][2] +
                mat_A[83][2] * mat_B[119][2] +
                mat_A[83][3] * mat_B[127][2] +
                mat_A[84][0] * mat_B[135][2] +
                mat_A[84][1] * mat_B[143][2] +
                mat_A[84][2] * mat_B[151][2] +
                mat_A[84][3] * mat_B[159][2] +
                mat_A[85][0] * mat_B[167][2] +
                mat_A[85][1] * mat_B[175][2] +
                mat_A[85][2] * mat_B[183][2] +
                mat_A[85][3] * mat_B[191][2] +
                mat_A[86][0] * mat_B[199][2] +
                mat_A[86][1] * mat_B[207][2] +
                mat_A[86][2] * mat_B[215][2] +
                mat_A[86][3] * mat_B[223][2] +
                mat_A[87][0] * mat_B[231][2] +
                mat_A[87][1] * mat_B[239][2] +
                mat_A[87][2] * mat_B[247][2] +
                mat_A[87][3] * mat_B[255][2];
    mat_C[87][3] <=
                mat_A[80][0] * mat_B[7][3] +
                mat_A[80][1] * mat_B[15][3] +
                mat_A[80][2] * mat_B[23][3] +
                mat_A[80][3] * mat_B[31][3] +
                mat_A[81][0] * mat_B[39][3] +
                mat_A[81][1] * mat_B[47][3] +
                mat_A[81][2] * mat_B[55][3] +
                mat_A[81][3] * mat_B[63][3] +
                mat_A[82][0] * mat_B[71][3] +
                mat_A[82][1] * mat_B[79][3] +
                mat_A[82][2] * mat_B[87][3] +
                mat_A[82][3] * mat_B[95][3] +
                mat_A[83][0] * mat_B[103][3] +
                mat_A[83][1] * mat_B[111][3] +
                mat_A[83][2] * mat_B[119][3] +
                mat_A[83][3] * mat_B[127][3] +
                mat_A[84][0] * mat_B[135][3] +
                mat_A[84][1] * mat_B[143][3] +
                mat_A[84][2] * mat_B[151][3] +
                mat_A[84][3] * mat_B[159][3] +
                mat_A[85][0] * mat_B[167][3] +
                mat_A[85][1] * mat_B[175][3] +
                mat_A[85][2] * mat_B[183][3] +
                mat_A[85][3] * mat_B[191][3] +
                mat_A[86][0] * mat_B[199][3] +
                mat_A[86][1] * mat_B[207][3] +
                mat_A[86][2] * mat_B[215][3] +
                mat_A[86][3] * mat_B[223][3] +
                mat_A[87][0] * mat_B[231][3] +
                mat_A[87][1] * mat_B[239][3] +
                mat_A[87][2] * mat_B[247][3] +
                mat_A[87][3] * mat_B[255][3];
    mat_C[88][0] <=
                mat_A[88][0] * mat_B[0][0] +
                mat_A[88][1] * mat_B[8][0] +
                mat_A[88][2] * mat_B[16][0] +
                mat_A[88][3] * mat_B[24][0] +
                mat_A[89][0] * mat_B[32][0] +
                mat_A[89][1] * mat_B[40][0] +
                mat_A[89][2] * mat_B[48][0] +
                mat_A[89][3] * mat_B[56][0] +
                mat_A[90][0] * mat_B[64][0] +
                mat_A[90][1] * mat_B[72][0] +
                mat_A[90][2] * mat_B[80][0] +
                mat_A[90][3] * mat_B[88][0] +
                mat_A[91][0] * mat_B[96][0] +
                mat_A[91][1] * mat_B[104][0] +
                mat_A[91][2] * mat_B[112][0] +
                mat_A[91][3] * mat_B[120][0] +
                mat_A[92][0] * mat_B[128][0] +
                mat_A[92][1] * mat_B[136][0] +
                mat_A[92][2] * mat_B[144][0] +
                mat_A[92][3] * mat_B[152][0] +
                mat_A[93][0] * mat_B[160][0] +
                mat_A[93][1] * mat_B[168][0] +
                mat_A[93][2] * mat_B[176][0] +
                mat_A[93][3] * mat_B[184][0] +
                mat_A[94][0] * mat_B[192][0] +
                mat_A[94][1] * mat_B[200][0] +
                mat_A[94][2] * mat_B[208][0] +
                mat_A[94][3] * mat_B[216][0] +
                mat_A[95][0] * mat_B[224][0] +
                mat_A[95][1] * mat_B[232][0] +
                mat_A[95][2] * mat_B[240][0] +
                mat_A[95][3] * mat_B[248][0];
    mat_C[88][1] <=
                mat_A[88][0] * mat_B[0][1] +
                mat_A[88][1] * mat_B[8][1] +
                mat_A[88][2] * mat_B[16][1] +
                mat_A[88][3] * mat_B[24][1] +
                mat_A[89][0] * mat_B[32][1] +
                mat_A[89][1] * mat_B[40][1] +
                mat_A[89][2] * mat_B[48][1] +
                mat_A[89][3] * mat_B[56][1] +
                mat_A[90][0] * mat_B[64][1] +
                mat_A[90][1] * mat_B[72][1] +
                mat_A[90][2] * mat_B[80][1] +
                mat_A[90][3] * mat_B[88][1] +
                mat_A[91][0] * mat_B[96][1] +
                mat_A[91][1] * mat_B[104][1] +
                mat_A[91][2] * mat_B[112][1] +
                mat_A[91][3] * mat_B[120][1] +
                mat_A[92][0] * mat_B[128][1] +
                mat_A[92][1] * mat_B[136][1] +
                mat_A[92][2] * mat_B[144][1] +
                mat_A[92][3] * mat_B[152][1] +
                mat_A[93][0] * mat_B[160][1] +
                mat_A[93][1] * mat_B[168][1] +
                mat_A[93][2] * mat_B[176][1] +
                mat_A[93][3] * mat_B[184][1] +
                mat_A[94][0] * mat_B[192][1] +
                mat_A[94][1] * mat_B[200][1] +
                mat_A[94][2] * mat_B[208][1] +
                mat_A[94][3] * mat_B[216][1] +
                mat_A[95][0] * mat_B[224][1] +
                mat_A[95][1] * mat_B[232][1] +
                mat_A[95][2] * mat_B[240][1] +
                mat_A[95][3] * mat_B[248][1];
    mat_C[88][2] <=
                mat_A[88][0] * mat_B[0][2] +
                mat_A[88][1] * mat_B[8][2] +
                mat_A[88][2] * mat_B[16][2] +
                mat_A[88][3] * mat_B[24][2] +
                mat_A[89][0] * mat_B[32][2] +
                mat_A[89][1] * mat_B[40][2] +
                mat_A[89][2] * mat_B[48][2] +
                mat_A[89][3] * mat_B[56][2] +
                mat_A[90][0] * mat_B[64][2] +
                mat_A[90][1] * mat_B[72][2] +
                mat_A[90][2] * mat_B[80][2] +
                mat_A[90][3] * mat_B[88][2] +
                mat_A[91][0] * mat_B[96][2] +
                mat_A[91][1] * mat_B[104][2] +
                mat_A[91][2] * mat_B[112][2] +
                mat_A[91][3] * mat_B[120][2] +
                mat_A[92][0] * mat_B[128][2] +
                mat_A[92][1] * mat_B[136][2] +
                mat_A[92][2] * mat_B[144][2] +
                mat_A[92][3] * mat_B[152][2] +
                mat_A[93][0] * mat_B[160][2] +
                mat_A[93][1] * mat_B[168][2] +
                mat_A[93][2] * mat_B[176][2] +
                mat_A[93][3] * mat_B[184][2] +
                mat_A[94][0] * mat_B[192][2] +
                mat_A[94][1] * mat_B[200][2] +
                mat_A[94][2] * mat_B[208][2] +
                mat_A[94][3] * mat_B[216][2] +
                mat_A[95][0] * mat_B[224][2] +
                mat_A[95][1] * mat_B[232][2] +
                mat_A[95][2] * mat_B[240][2] +
                mat_A[95][3] * mat_B[248][2];
    mat_C[88][3] <=
                mat_A[88][0] * mat_B[0][3] +
                mat_A[88][1] * mat_B[8][3] +
                mat_A[88][2] * mat_B[16][3] +
                mat_A[88][3] * mat_B[24][3] +
                mat_A[89][0] * mat_B[32][3] +
                mat_A[89][1] * mat_B[40][3] +
                mat_A[89][2] * mat_B[48][3] +
                mat_A[89][3] * mat_B[56][3] +
                mat_A[90][0] * mat_B[64][3] +
                mat_A[90][1] * mat_B[72][3] +
                mat_A[90][2] * mat_B[80][3] +
                mat_A[90][3] * mat_B[88][3] +
                mat_A[91][0] * mat_B[96][3] +
                mat_A[91][1] * mat_B[104][3] +
                mat_A[91][2] * mat_B[112][3] +
                mat_A[91][3] * mat_B[120][3] +
                mat_A[92][0] * mat_B[128][3] +
                mat_A[92][1] * mat_B[136][3] +
                mat_A[92][2] * mat_B[144][3] +
                mat_A[92][3] * mat_B[152][3] +
                mat_A[93][0] * mat_B[160][3] +
                mat_A[93][1] * mat_B[168][3] +
                mat_A[93][2] * mat_B[176][3] +
                mat_A[93][3] * mat_B[184][3] +
                mat_A[94][0] * mat_B[192][3] +
                mat_A[94][1] * mat_B[200][3] +
                mat_A[94][2] * mat_B[208][3] +
                mat_A[94][3] * mat_B[216][3] +
                mat_A[95][0] * mat_B[224][3] +
                mat_A[95][1] * mat_B[232][3] +
                mat_A[95][2] * mat_B[240][3] +
                mat_A[95][3] * mat_B[248][3];
    mat_C[89][0] <=
                mat_A[88][0] * mat_B[1][0] +
                mat_A[88][1] * mat_B[9][0] +
                mat_A[88][2] * mat_B[17][0] +
                mat_A[88][3] * mat_B[25][0] +
                mat_A[89][0] * mat_B[33][0] +
                mat_A[89][1] * mat_B[41][0] +
                mat_A[89][2] * mat_B[49][0] +
                mat_A[89][3] * mat_B[57][0] +
                mat_A[90][0] * mat_B[65][0] +
                mat_A[90][1] * mat_B[73][0] +
                mat_A[90][2] * mat_B[81][0] +
                mat_A[90][3] * mat_B[89][0] +
                mat_A[91][0] * mat_B[97][0] +
                mat_A[91][1] * mat_B[105][0] +
                mat_A[91][2] * mat_B[113][0] +
                mat_A[91][3] * mat_B[121][0] +
                mat_A[92][0] * mat_B[129][0] +
                mat_A[92][1] * mat_B[137][0] +
                mat_A[92][2] * mat_B[145][0] +
                mat_A[92][3] * mat_B[153][0] +
                mat_A[93][0] * mat_B[161][0] +
                mat_A[93][1] * mat_B[169][0] +
                mat_A[93][2] * mat_B[177][0] +
                mat_A[93][3] * mat_B[185][0] +
                mat_A[94][0] * mat_B[193][0] +
                mat_A[94][1] * mat_B[201][0] +
                mat_A[94][2] * mat_B[209][0] +
                mat_A[94][3] * mat_B[217][0] +
                mat_A[95][0] * mat_B[225][0] +
                mat_A[95][1] * mat_B[233][0] +
                mat_A[95][2] * mat_B[241][0] +
                mat_A[95][3] * mat_B[249][0];
    mat_C[89][1] <=
                mat_A[88][0] * mat_B[1][1] +
                mat_A[88][1] * mat_B[9][1] +
                mat_A[88][2] * mat_B[17][1] +
                mat_A[88][3] * mat_B[25][1] +
                mat_A[89][0] * mat_B[33][1] +
                mat_A[89][1] * mat_B[41][1] +
                mat_A[89][2] * mat_B[49][1] +
                mat_A[89][3] * mat_B[57][1] +
                mat_A[90][0] * mat_B[65][1] +
                mat_A[90][1] * mat_B[73][1] +
                mat_A[90][2] * mat_B[81][1] +
                mat_A[90][3] * mat_B[89][1] +
                mat_A[91][0] * mat_B[97][1] +
                mat_A[91][1] * mat_B[105][1] +
                mat_A[91][2] * mat_B[113][1] +
                mat_A[91][3] * mat_B[121][1] +
                mat_A[92][0] * mat_B[129][1] +
                mat_A[92][1] * mat_B[137][1] +
                mat_A[92][2] * mat_B[145][1] +
                mat_A[92][3] * mat_B[153][1] +
                mat_A[93][0] * mat_B[161][1] +
                mat_A[93][1] * mat_B[169][1] +
                mat_A[93][2] * mat_B[177][1] +
                mat_A[93][3] * mat_B[185][1] +
                mat_A[94][0] * mat_B[193][1] +
                mat_A[94][1] * mat_B[201][1] +
                mat_A[94][2] * mat_B[209][1] +
                mat_A[94][3] * mat_B[217][1] +
                mat_A[95][0] * mat_B[225][1] +
                mat_A[95][1] * mat_B[233][1] +
                mat_A[95][2] * mat_B[241][1] +
                mat_A[95][3] * mat_B[249][1];
    mat_C[89][2] <=
                mat_A[88][0] * mat_B[1][2] +
                mat_A[88][1] * mat_B[9][2] +
                mat_A[88][2] * mat_B[17][2] +
                mat_A[88][3] * mat_B[25][2] +
                mat_A[89][0] * mat_B[33][2] +
                mat_A[89][1] * mat_B[41][2] +
                mat_A[89][2] * mat_B[49][2] +
                mat_A[89][3] * mat_B[57][2] +
                mat_A[90][0] * mat_B[65][2] +
                mat_A[90][1] * mat_B[73][2] +
                mat_A[90][2] * mat_B[81][2] +
                mat_A[90][3] * mat_B[89][2] +
                mat_A[91][0] * mat_B[97][2] +
                mat_A[91][1] * mat_B[105][2] +
                mat_A[91][2] * mat_B[113][2] +
                mat_A[91][3] * mat_B[121][2] +
                mat_A[92][0] * mat_B[129][2] +
                mat_A[92][1] * mat_B[137][2] +
                mat_A[92][2] * mat_B[145][2] +
                mat_A[92][3] * mat_B[153][2] +
                mat_A[93][0] * mat_B[161][2] +
                mat_A[93][1] * mat_B[169][2] +
                mat_A[93][2] * mat_B[177][2] +
                mat_A[93][3] * mat_B[185][2] +
                mat_A[94][0] * mat_B[193][2] +
                mat_A[94][1] * mat_B[201][2] +
                mat_A[94][2] * mat_B[209][2] +
                mat_A[94][3] * mat_B[217][2] +
                mat_A[95][0] * mat_B[225][2] +
                mat_A[95][1] * mat_B[233][2] +
                mat_A[95][2] * mat_B[241][2] +
                mat_A[95][3] * mat_B[249][2];
    mat_C[89][3] <=
                mat_A[88][0] * mat_B[1][3] +
                mat_A[88][1] * mat_B[9][3] +
                mat_A[88][2] * mat_B[17][3] +
                mat_A[88][3] * mat_B[25][3] +
                mat_A[89][0] * mat_B[33][3] +
                mat_A[89][1] * mat_B[41][3] +
                mat_A[89][2] * mat_B[49][3] +
                mat_A[89][3] * mat_B[57][3] +
                mat_A[90][0] * mat_B[65][3] +
                mat_A[90][1] * mat_B[73][3] +
                mat_A[90][2] * mat_B[81][3] +
                mat_A[90][3] * mat_B[89][3] +
                mat_A[91][0] * mat_B[97][3] +
                mat_A[91][1] * mat_B[105][3] +
                mat_A[91][2] * mat_B[113][3] +
                mat_A[91][3] * mat_B[121][3] +
                mat_A[92][0] * mat_B[129][3] +
                mat_A[92][1] * mat_B[137][3] +
                mat_A[92][2] * mat_B[145][3] +
                mat_A[92][3] * mat_B[153][3] +
                mat_A[93][0] * mat_B[161][3] +
                mat_A[93][1] * mat_B[169][3] +
                mat_A[93][2] * mat_B[177][3] +
                mat_A[93][3] * mat_B[185][3] +
                mat_A[94][0] * mat_B[193][3] +
                mat_A[94][1] * mat_B[201][3] +
                mat_A[94][2] * mat_B[209][3] +
                mat_A[94][3] * mat_B[217][3] +
                mat_A[95][0] * mat_B[225][3] +
                mat_A[95][1] * mat_B[233][3] +
                mat_A[95][2] * mat_B[241][3] +
                mat_A[95][3] * mat_B[249][3];
    mat_C[90][0] <=
                mat_A[88][0] * mat_B[2][0] +
                mat_A[88][1] * mat_B[10][0] +
                mat_A[88][2] * mat_B[18][0] +
                mat_A[88][3] * mat_B[26][0] +
                mat_A[89][0] * mat_B[34][0] +
                mat_A[89][1] * mat_B[42][0] +
                mat_A[89][2] * mat_B[50][0] +
                mat_A[89][3] * mat_B[58][0] +
                mat_A[90][0] * mat_B[66][0] +
                mat_A[90][1] * mat_B[74][0] +
                mat_A[90][2] * mat_B[82][0] +
                mat_A[90][3] * mat_B[90][0] +
                mat_A[91][0] * mat_B[98][0] +
                mat_A[91][1] * mat_B[106][0] +
                mat_A[91][2] * mat_B[114][0] +
                mat_A[91][3] * mat_B[122][0] +
                mat_A[92][0] * mat_B[130][0] +
                mat_A[92][1] * mat_B[138][0] +
                mat_A[92][2] * mat_B[146][0] +
                mat_A[92][3] * mat_B[154][0] +
                mat_A[93][0] * mat_B[162][0] +
                mat_A[93][1] * mat_B[170][0] +
                mat_A[93][2] * mat_B[178][0] +
                mat_A[93][3] * mat_B[186][0] +
                mat_A[94][0] * mat_B[194][0] +
                mat_A[94][1] * mat_B[202][0] +
                mat_A[94][2] * mat_B[210][0] +
                mat_A[94][3] * mat_B[218][0] +
                mat_A[95][0] * mat_B[226][0] +
                mat_A[95][1] * mat_B[234][0] +
                mat_A[95][2] * mat_B[242][0] +
                mat_A[95][3] * mat_B[250][0];
    mat_C[90][1] <=
                mat_A[88][0] * mat_B[2][1] +
                mat_A[88][1] * mat_B[10][1] +
                mat_A[88][2] * mat_B[18][1] +
                mat_A[88][3] * mat_B[26][1] +
                mat_A[89][0] * mat_B[34][1] +
                mat_A[89][1] * mat_B[42][1] +
                mat_A[89][2] * mat_B[50][1] +
                mat_A[89][3] * mat_B[58][1] +
                mat_A[90][0] * mat_B[66][1] +
                mat_A[90][1] * mat_B[74][1] +
                mat_A[90][2] * mat_B[82][1] +
                mat_A[90][3] * mat_B[90][1] +
                mat_A[91][0] * mat_B[98][1] +
                mat_A[91][1] * mat_B[106][1] +
                mat_A[91][2] * mat_B[114][1] +
                mat_A[91][3] * mat_B[122][1] +
                mat_A[92][0] * mat_B[130][1] +
                mat_A[92][1] * mat_B[138][1] +
                mat_A[92][2] * mat_B[146][1] +
                mat_A[92][3] * mat_B[154][1] +
                mat_A[93][0] * mat_B[162][1] +
                mat_A[93][1] * mat_B[170][1] +
                mat_A[93][2] * mat_B[178][1] +
                mat_A[93][3] * mat_B[186][1] +
                mat_A[94][0] * mat_B[194][1] +
                mat_A[94][1] * mat_B[202][1] +
                mat_A[94][2] * mat_B[210][1] +
                mat_A[94][3] * mat_B[218][1] +
                mat_A[95][0] * mat_B[226][1] +
                mat_A[95][1] * mat_B[234][1] +
                mat_A[95][2] * mat_B[242][1] +
                mat_A[95][3] * mat_B[250][1];
    mat_C[90][2] <=
                mat_A[88][0] * mat_B[2][2] +
                mat_A[88][1] * mat_B[10][2] +
                mat_A[88][2] * mat_B[18][2] +
                mat_A[88][3] * mat_B[26][2] +
                mat_A[89][0] * mat_B[34][2] +
                mat_A[89][1] * mat_B[42][2] +
                mat_A[89][2] * mat_B[50][2] +
                mat_A[89][3] * mat_B[58][2] +
                mat_A[90][0] * mat_B[66][2] +
                mat_A[90][1] * mat_B[74][2] +
                mat_A[90][2] * mat_B[82][2] +
                mat_A[90][3] * mat_B[90][2] +
                mat_A[91][0] * mat_B[98][2] +
                mat_A[91][1] * mat_B[106][2] +
                mat_A[91][2] * mat_B[114][2] +
                mat_A[91][3] * mat_B[122][2] +
                mat_A[92][0] * mat_B[130][2] +
                mat_A[92][1] * mat_B[138][2] +
                mat_A[92][2] * mat_B[146][2] +
                mat_A[92][3] * mat_B[154][2] +
                mat_A[93][0] * mat_B[162][2] +
                mat_A[93][1] * mat_B[170][2] +
                mat_A[93][2] * mat_B[178][2] +
                mat_A[93][3] * mat_B[186][2] +
                mat_A[94][0] * mat_B[194][2] +
                mat_A[94][1] * mat_B[202][2] +
                mat_A[94][2] * mat_B[210][2] +
                mat_A[94][3] * mat_B[218][2] +
                mat_A[95][0] * mat_B[226][2] +
                mat_A[95][1] * mat_B[234][2] +
                mat_A[95][2] * mat_B[242][2] +
                mat_A[95][3] * mat_B[250][2];
    mat_C[90][3] <=
                mat_A[88][0] * mat_B[2][3] +
                mat_A[88][1] * mat_B[10][3] +
                mat_A[88][2] * mat_B[18][3] +
                mat_A[88][3] * mat_B[26][3] +
                mat_A[89][0] * mat_B[34][3] +
                mat_A[89][1] * mat_B[42][3] +
                mat_A[89][2] * mat_B[50][3] +
                mat_A[89][3] * mat_B[58][3] +
                mat_A[90][0] * mat_B[66][3] +
                mat_A[90][1] * mat_B[74][3] +
                mat_A[90][2] * mat_B[82][3] +
                mat_A[90][3] * mat_B[90][3] +
                mat_A[91][0] * mat_B[98][3] +
                mat_A[91][1] * mat_B[106][3] +
                mat_A[91][2] * mat_B[114][3] +
                mat_A[91][3] * mat_B[122][3] +
                mat_A[92][0] * mat_B[130][3] +
                mat_A[92][1] * mat_B[138][3] +
                mat_A[92][2] * mat_B[146][3] +
                mat_A[92][3] * mat_B[154][3] +
                mat_A[93][0] * mat_B[162][3] +
                mat_A[93][1] * mat_B[170][3] +
                mat_A[93][2] * mat_B[178][3] +
                mat_A[93][3] * mat_B[186][3] +
                mat_A[94][0] * mat_B[194][3] +
                mat_A[94][1] * mat_B[202][3] +
                mat_A[94][2] * mat_B[210][3] +
                mat_A[94][3] * mat_B[218][3] +
                mat_A[95][0] * mat_B[226][3] +
                mat_A[95][1] * mat_B[234][3] +
                mat_A[95][2] * mat_B[242][3] +
                mat_A[95][3] * mat_B[250][3];
    mat_C[91][0] <=
                mat_A[88][0] * mat_B[3][0] +
                mat_A[88][1] * mat_B[11][0] +
                mat_A[88][2] * mat_B[19][0] +
                mat_A[88][3] * mat_B[27][0] +
                mat_A[89][0] * mat_B[35][0] +
                mat_A[89][1] * mat_B[43][0] +
                mat_A[89][2] * mat_B[51][0] +
                mat_A[89][3] * mat_B[59][0] +
                mat_A[90][0] * mat_B[67][0] +
                mat_A[90][1] * mat_B[75][0] +
                mat_A[90][2] * mat_B[83][0] +
                mat_A[90][3] * mat_B[91][0] +
                mat_A[91][0] * mat_B[99][0] +
                mat_A[91][1] * mat_B[107][0] +
                mat_A[91][2] * mat_B[115][0] +
                mat_A[91][3] * mat_B[123][0] +
                mat_A[92][0] * mat_B[131][0] +
                mat_A[92][1] * mat_B[139][0] +
                mat_A[92][2] * mat_B[147][0] +
                mat_A[92][3] * mat_B[155][0] +
                mat_A[93][0] * mat_B[163][0] +
                mat_A[93][1] * mat_B[171][0] +
                mat_A[93][2] * mat_B[179][0] +
                mat_A[93][3] * mat_B[187][0] +
                mat_A[94][0] * mat_B[195][0] +
                mat_A[94][1] * mat_B[203][0] +
                mat_A[94][2] * mat_B[211][0] +
                mat_A[94][3] * mat_B[219][0] +
                mat_A[95][0] * mat_B[227][0] +
                mat_A[95][1] * mat_B[235][0] +
                mat_A[95][2] * mat_B[243][0] +
                mat_A[95][3] * mat_B[251][0];
    mat_C[91][1] <=
                mat_A[88][0] * mat_B[3][1] +
                mat_A[88][1] * mat_B[11][1] +
                mat_A[88][2] * mat_B[19][1] +
                mat_A[88][3] * mat_B[27][1] +
                mat_A[89][0] * mat_B[35][1] +
                mat_A[89][1] * mat_B[43][1] +
                mat_A[89][2] * mat_B[51][1] +
                mat_A[89][3] * mat_B[59][1] +
                mat_A[90][0] * mat_B[67][1] +
                mat_A[90][1] * mat_B[75][1] +
                mat_A[90][2] * mat_B[83][1] +
                mat_A[90][3] * mat_B[91][1] +
                mat_A[91][0] * mat_B[99][1] +
                mat_A[91][1] * mat_B[107][1] +
                mat_A[91][2] * mat_B[115][1] +
                mat_A[91][3] * mat_B[123][1] +
                mat_A[92][0] * mat_B[131][1] +
                mat_A[92][1] * mat_B[139][1] +
                mat_A[92][2] * mat_B[147][1] +
                mat_A[92][3] * mat_B[155][1] +
                mat_A[93][0] * mat_B[163][1] +
                mat_A[93][1] * mat_B[171][1] +
                mat_A[93][2] * mat_B[179][1] +
                mat_A[93][3] * mat_B[187][1] +
                mat_A[94][0] * mat_B[195][1] +
                mat_A[94][1] * mat_B[203][1] +
                mat_A[94][2] * mat_B[211][1] +
                mat_A[94][3] * mat_B[219][1] +
                mat_A[95][0] * mat_B[227][1] +
                mat_A[95][1] * mat_B[235][1] +
                mat_A[95][2] * mat_B[243][1] +
                mat_A[95][3] * mat_B[251][1];
    mat_C[91][2] <=
                mat_A[88][0] * mat_B[3][2] +
                mat_A[88][1] * mat_B[11][2] +
                mat_A[88][2] * mat_B[19][2] +
                mat_A[88][3] * mat_B[27][2] +
                mat_A[89][0] * mat_B[35][2] +
                mat_A[89][1] * mat_B[43][2] +
                mat_A[89][2] * mat_B[51][2] +
                mat_A[89][3] * mat_B[59][2] +
                mat_A[90][0] * mat_B[67][2] +
                mat_A[90][1] * mat_B[75][2] +
                mat_A[90][2] * mat_B[83][2] +
                mat_A[90][3] * mat_B[91][2] +
                mat_A[91][0] * mat_B[99][2] +
                mat_A[91][1] * mat_B[107][2] +
                mat_A[91][2] * mat_B[115][2] +
                mat_A[91][3] * mat_B[123][2] +
                mat_A[92][0] * mat_B[131][2] +
                mat_A[92][1] * mat_B[139][2] +
                mat_A[92][2] * mat_B[147][2] +
                mat_A[92][3] * mat_B[155][2] +
                mat_A[93][0] * mat_B[163][2] +
                mat_A[93][1] * mat_B[171][2] +
                mat_A[93][2] * mat_B[179][2] +
                mat_A[93][3] * mat_B[187][2] +
                mat_A[94][0] * mat_B[195][2] +
                mat_A[94][1] * mat_B[203][2] +
                mat_A[94][2] * mat_B[211][2] +
                mat_A[94][3] * mat_B[219][2] +
                mat_A[95][0] * mat_B[227][2] +
                mat_A[95][1] * mat_B[235][2] +
                mat_A[95][2] * mat_B[243][2] +
                mat_A[95][3] * mat_B[251][2];
    mat_C[91][3] <=
                mat_A[88][0] * mat_B[3][3] +
                mat_A[88][1] * mat_B[11][3] +
                mat_A[88][2] * mat_B[19][3] +
                mat_A[88][3] * mat_B[27][3] +
                mat_A[89][0] * mat_B[35][3] +
                mat_A[89][1] * mat_B[43][3] +
                mat_A[89][2] * mat_B[51][3] +
                mat_A[89][3] * mat_B[59][3] +
                mat_A[90][0] * mat_B[67][3] +
                mat_A[90][1] * mat_B[75][3] +
                mat_A[90][2] * mat_B[83][3] +
                mat_A[90][3] * mat_B[91][3] +
                mat_A[91][0] * mat_B[99][3] +
                mat_A[91][1] * mat_B[107][3] +
                mat_A[91][2] * mat_B[115][3] +
                mat_A[91][3] * mat_B[123][3] +
                mat_A[92][0] * mat_B[131][3] +
                mat_A[92][1] * mat_B[139][3] +
                mat_A[92][2] * mat_B[147][3] +
                mat_A[92][3] * mat_B[155][3] +
                mat_A[93][0] * mat_B[163][3] +
                mat_A[93][1] * mat_B[171][3] +
                mat_A[93][2] * mat_B[179][3] +
                mat_A[93][3] * mat_B[187][3] +
                mat_A[94][0] * mat_B[195][3] +
                mat_A[94][1] * mat_B[203][3] +
                mat_A[94][2] * mat_B[211][3] +
                mat_A[94][3] * mat_B[219][3] +
                mat_A[95][0] * mat_B[227][3] +
                mat_A[95][1] * mat_B[235][3] +
                mat_A[95][2] * mat_B[243][3] +
                mat_A[95][3] * mat_B[251][3];
    mat_C[92][0] <=
                mat_A[88][0] * mat_B[4][0] +
                mat_A[88][1] * mat_B[12][0] +
                mat_A[88][2] * mat_B[20][0] +
                mat_A[88][3] * mat_B[28][0] +
                mat_A[89][0] * mat_B[36][0] +
                mat_A[89][1] * mat_B[44][0] +
                mat_A[89][2] * mat_B[52][0] +
                mat_A[89][3] * mat_B[60][0] +
                mat_A[90][0] * mat_B[68][0] +
                mat_A[90][1] * mat_B[76][0] +
                mat_A[90][2] * mat_B[84][0] +
                mat_A[90][3] * mat_B[92][0] +
                mat_A[91][0] * mat_B[100][0] +
                mat_A[91][1] * mat_B[108][0] +
                mat_A[91][2] * mat_B[116][0] +
                mat_A[91][3] * mat_B[124][0] +
                mat_A[92][0] * mat_B[132][0] +
                mat_A[92][1] * mat_B[140][0] +
                mat_A[92][2] * mat_B[148][0] +
                mat_A[92][3] * mat_B[156][0] +
                mat_A[93][0] * mat_B[164][0] +
                mat_A[93][1] * mat_B[172][0] +
                mat_A[93][2] * mat_B[180][0] +
                mat_A[93][3] * mat_B[188][0] +
                mat_A[94][0] * mat_B[196][0] +
                mat_A[94][1] * mat_B[204][0] +
                mat_A[94][2] * mat_B[212][0] +
                mat_A[94][3] * mat_B[220][0] +
                mat_A[95][0] * mat_B[228][0] +
                mat_A[95][1] * mat_B[236][0] +
                mat_A[95][2] * mat_B[244][0] +
                mat_A[95][3] * mat_B[252][0];
    mat_C[92][1] <=
                mat_A[88][0] * mat_B[4][1] +
                mat_A[88][1] * mat_B[12][1] +
                mat_A[88][2] * mat_B[20][1] +
                mat_A[88][3] * mat_B[28][1] +
                mat_A[89][0] * mat_B[36][1] +
                mat_A[89][1] * mat_B[44][1] +
                mat_A[89][2] * mat_B[52][1] +
                mat_A[89][3] * mat_B[60][1] +
                mat_A[90][0] * mat_B[68][1] +
                mat_A[90][1] * mat_B[76][1] +
                mat_A[90][2] * mat_B[84][1] +
                mat_A[90][3] * mat_B[92][1] +
                mat_A[91][0] * mat_B[100][1] +
                mat_A[91][1] * mat_B[108][1] +
                mat_A[91][2] * mat_B[116][1] +
                mat_A[91][3] * mat_B[124][1] +
                mat_A[92][0] * mat_B[132][1] +
                mat_A[92][1] * mat_B[140][1] +
                mat_A[92][2] * mat_B[148][1] +
                mat_A[92][3] * mat_B[156][1] +
                mat_A[93][0] * mat_B[164][1] +
                mat_A[93][1] * mat_B[172][1] +
                mat_A[93][2] * mat_B[180][1] +
                mat_A[93][3] * mat_B[188][1] +
                mat_A[94][0] * mat_B[196][1] +
                mat_A[94][1] * mat_B[204][1] +
                mat_A[94][2] * mat_B[212][1] +
                mat_A[94][3] * mat_B[220][1] +
                mat_A[95][0] * mat_B[228][1] +
                mat_A[95][1] * mat_B[236][1] +
                mat_A[95][2] * mat_B[244][1] +
                mat_A[95][3] * mat_B[252][1];
    mat_C[92][2] <=
                mat_A[88][0] * mat_B[4][2] +
                mat_A[88][1] * mat_B[12][2] +
                mat_A[88][2] * mat_B[20][2] +
                mat_A[88][3] * mat_B[28][2] +
                mat_A[89][0] * mat_B[36][2] +
                mat_A[89][1] * mat_B[44][2] +
                mat_A[89][2] * mat_B[52][2] +
                mat_A[89][3] * mat_B[60][2] +
                mat_A[90][0] * mat_B[68][2] +
                mat_A[90][1] * mat_B[76][2] +
                mat_A[90][2] * mat_B[84][2] +
                mat_A[90][3] * mat_B[92][2] +
                mat_A[91][0] * mat_B[100][2] +
                mat_A[91][1] * mat_B[108][2] +
                mat_A[91][2] * mat_B[116][2] +
                mat_A[91][3] * mat_B[124][2] +
                mat_A[92][0] * mat_B[132][2] +
                mat_A[92][1] * mat_B[140][2] +
                mat_A[92][2] * mat_B[148][2] +
                mat_A[92][3] * mat_B[156][2] +
                mat_A[93][0] * mat_B[164][2] +
                mat_A[93][1] * mat_B[172][2] +
                mat_A[93][2] * mat_B[180][2] +
                mat_A[93][3] * mat_B[188][2] +
                mat_A[94][0] * mat_B[196][2] +
                mat_A[94][1] * mat_B[204][2] +
                mat_A[94][2] * mat_B[212][2] +
                mat_A[94][3] * mat_B[220][2] +
                mat_A[95][0] * mat_B[228][2] +
                mat_A[95][1] * mat_B[236][2] +
                mat_A[95][2] * mat_B[244][2] +
                mat_A[95][3] * mat_B[252][2];
    mat_C[92][3] <=
                mat_A[88][0] * mat_B[4][3] +
                mat_A[88][1] * mat_B[12][3] +
                mat_A[88][2] * mat_B[20][3] +
                mat_A[88][3] * mat_B[28][3] +
                mat_A[89][0] * mat_B[36][3] +
                mat_A[89][1] * mat_B[44][3] +
                mat_A[89][2] * mat_B[52][3] +
                mat_A[89][3] * mat_B[60][3] +
                mat_A[90][0] * mat_B[68][3] +
                mat_A[90][1] * mat_B[76][3] +
                mat_A[90][2] * mat_B[84][3] +
                mat_A[90][3] * mat_B[92][3] +
                mat_A[91][0] * mat_B[100][3] +
                mat_A[91][1] * mat_B[108][3] +
                mat_A[91][2] * mat_B[116][3] +
                mat_A[91][3] * mat_B[124][3] +
                mat_A[92][0] * mat_B[132][3] +
                mat_A[92][1] * mat_B[140][3] +
                mat_A[92][2] * mat_B[148][3] +
                mat_A[92][3] * mat_B[156][3] +
                mat_A[93][0] * mat_B[164][3] +
                mat_A[93][1] * mat_B[172][3] +
                mat_A[93][2] * mat_B[180][3] +
                mat_A[93][3] * mat_B[188][3] +
                mat_A[94][0] * mat_B[196][3] +
                mat_A[94][1] * mat_B[204][3] +
                mat_A[94][2] * mat_B[212][3] +
                mat_A[94][3] * mat_B[220][3] +
                mat_A[95][0] * mat_B[228][3] +
                mat_A[95][1] * mat_B[236][3] +
                mat_A[95][2] * mat_B[244][3] +
                mat_A[95][3] * mat_B[252][3];
    mat_C[93][0] <=
                mat_A[88][0] * mat_B[5][0] +
                mat_A[88][1] * mat_B[13][0] +
                mat_A[88][2] * mat_B[21][0] +
                mat_A[88][3] * mat_B[29][0] +
                mat_A[89][0] * mat_B[37][0] +
                mat_A[89][1] * mat_B[45][0] +
                mat_A[89][2] * mat_B[53][0] +
                mat_A[89][3] * mat_B[61][0] +
                mat_A[90][0] * mat_B[69][0] +
                mat_A[90][1] * mat_B[77][0] +
                mat_A[90][2] * mat_B[85][0] +
                mat_A[90][3] * mat_B[93][0] +
                mat_A[91][0] * mat_B[101][0] +
                mat_A[91][1] * mat_B[109][0] +
                mat_A[91][2] * mat_B[117][0] +
                mat_A[91][3] * mat_B[125][0] +
                mat_A[92][0] * mat_B[133][0] +
                mat_A[92][1] * mat_B[141][0] +
                mat_A[92][2] * mat_B[149][0] +
                mat_A[92][3] * mat_B[157][0] +
                mat_A[93][0] * mat_B[165][0] +
                mat_A[93][1] * mat_B[173][0] +
                mat_A[93][2] * mat_B[181][0] +
                mat_A[93][3] * mat_B[189][0] +
                mat_A[94][0] * mat_B[197][0] +
                mat_A[94][1] * mat_B[205][0] +
                mat_A[94][2] * mat_B[213][0] +
                mat_A[94][3] * mat_B[221][0] +
                mat_A[95][0] * mat_B[229][0] +
                mat_A[95][1] * mat_B[237][0] +
                mat_A[95][2] * mat_B[245][0] +
                mat_A[95][3] * mat_B[253][0];
    mat_C[93][1] <=
                mat_A[88][0] * mat_B[5][1] +
                mat_A[88][1] * mat_B[13][1] +
                mat_A[88][2] * mat_B[21][1] +
                mat_A[88][3] * mat_B[29][1] +
                mat_A[89][0] * mat_B[37][1] +
                mat_A[89][1] * mat_B[45][1] +
                mat_A[89][2] * mat_B[53][1] +
                mat_A[89][3] * mat_B[61][1] +
                mat_A[90][0] * mat_B[69][1] +
                mat_A[90][1] * mat_B[77][1] +
                mat_A[90][2] * mat_B[85][1] +
                mat_A[90][3] * mat_B[93][1] +
                mat_A[91][0] * mat_B[101][1] +
                mat_A[91][1] * mat_B[109][1] +
                mat_A[91][2] * mat_B[117][1] +
                mat_A[91][3] * mat_B[125][1] +
                mat_A[92][0] * mat_B[133][1] +
                mat_A[92][1] * mat_B[141][1] +
                mat_A[92][2] * mat_B[149][1] +
                mat_A[92][3] * mat_B[157][1] +
                mat_A[93][0] * mat_B[165][1] +
                mat_A[93][1] * mat_B[173][1] +
                mat_A[93][2] * mat_B[181][1] +
                mat_A[93][3] * mat_B[189][1] +
                mat_A[94][0] * mat_B[197][1] +
                mat_A[94][1] * mat_B[205][1] +
                mat_A[94][2] * mat_B[213][1] +
                mat_A[94][3] * mat_B[221][1] +
                mat_A[95][0] * mat_B[229][1] +
                mat_A[95][1] * mat_B[237][1] +
                mat_A[95][2] * mat_B[245][1] +
                mat_A[95][3] * mat_B[253][1];
    mat_C[93][2] <=
                mat_A[88][0] * mat_B[5][2] +
                mat_A[88][1] * mat_B[13][2] +
                mat_A[88][2] * mat_B[21][2] +
                mat_A[88][3] * mat_B[29][2] +
                mat_A[89][0] * mat_B[37][2] +
                mat_A[89][1] * mat_B[45][2] +
                mat_A[89][2] * mat_B[53][2] +
                mat_A[89][3] * mat_B[61][2] +
                mat_A[90][0] * mat_B[69][2] +
                mat_A[90][1] * mat_B[77][2] +
                mat_A[90][2] * mat_B[85][2] +
                mat_A[90][3] * mat_B[93][2] +
                mat_A[91][0] * mat_B[101][2] +
                mat_A[91][1] * mat_B[109][2] +
                mat_A[91][2] * mat_B[117][2] +
                mat_A[91][3] * mat_B[125][2] +
                mat_A[92][0] * mat_B[133][2] +
                mat_A[92][1] * mat_B[141][2] +
                mat_A[92][2] * mat_B[149][2] +
                mat_A[92][3] * mat_B[157][2] +
                mat_A[93][0] * mat_B[165][2] +
                mat_A[93][1] * mat_B[173][2] +
                mat_A[93][2] * mat_B[181][2] +
                mat_A[93][3] * mat_B[189][2] +
                mat_A[94][0] * mat_B[197][2] +
                mat_A[94][1] * mat_B[205][2] +
                mat_A[94][2] * mat_B[213][2] +
                mat_A[94][3] * mat_B[221][2] +
                mat_A[95][0] * mat_B[229][2] +
                mat_A[95][1] * mat_B[237][2] +
                mat_A[95][2] * mat_B[245][2] +
                mat_A[95][3] * mat_B[253][2];
    mat_C[93][3] <=
                mat_A[88][0] * mat_B[5][3] +
                mat_A[88][1] * mat_B[13][3] +
                mat_A[88][2] * mat_B[21][3] +
                mat_A[88][3] * mat_B[29][3] +
                mat_A[89][0] * mat_B[37][3] +
                mat_A[89][1] * mat_B[45][3] +
                mat_A[89][2] * mat_B[53][3] +
                mat_A[89][3] * mat_B[61][3] +
                mat_A[90][0] * mat_B[69][3] +
                mat_A[90][1] * mat_B[77][3] +
                mat_A[90][2] * mat_B[85][3] +
                mat_A[90][3] * mat_B[93][3] +
                mat_A[91][0] * mat_B[101][3] +
                mat_A[91][1] * mat_B[109][3] +
                mat_A[91][2] * mat_B[117][3] +
                mat_A[91][3] * mat_B[125][3] +
                mat_A[92][0] * mat_B[133][3] +
                mat_A[92][1] * mat_B[141][3] +
                mat_A[92][2] * mat_B[149][3] +
                mat_A[92][3] * mat_B[157][3] +
                mat_A[93][0] * mat_B[165][3] +
                mat_A[93][1] * mat_B[173][3] +
                mat_A[93][2] * mat_B[181][3] +
                mat_A[93][3] * mat_B[189][3] +
                mat_A[94][0] * mat_B[197][3] +
                mat_A[94][1] * mat_B[205][3] +
                mat_A[94][2] * mat_B[213][3] +
                mat_A[94][3] * mat_B[221][3] +
                mat_A[95][0] * mat_B[229][3] +
                mat_A[95][1] * mat_B[237][3] +
                mat_A[95][2] * mat_B[245][3] +
                mat_A[95][3] * mat_B[253][3];
    mat_C[94][0] <=
                mat_A[88][0] * mat_B[6][0] +
                mat_A[88][1] * mat_B[14][0] +
                mat_A[88][2] * mat_B[22][0] +
                mat_A[88][3] * mat_B[30][0] +
                mat_A[89][0] * mat_B[38][0] +
                mat_A[89][1] * mat_B[46][0] +
                mat_A[89][2] * mat_B[54][0] +
                mat_A[89][3] * mat_B[62][0] +
                mat_A[90][0] * mat_B[70][0] +
                mat_A[90][1] * mat_B[78][0] +
                mat_A[90][2] * mat_B[86][0] +
                mat_A[90][3] * mat_B[94][0] +
                mat_A[91][0] * mat_B[102][0] +
                mat_A[91][1] * mat_B[110][0] +
                mat_A[91][2] * mat_B[118][0] +
                mat_A[91][3] * mat_B[126][0] +
                mat_A[92][0] * mat_B[134][0] +
                mat_A[92][1] * mat_B[142][0] +
                mat_A[92][2] * mat_B[150][0] +
                mat_A[92][3] * mat_B[158][0] +
                mat_A[93][0] * mat_B[166][0] +
                mat_A[93][1] * mat_B[174][0] +
                mat_A[93][2] * mat_B[182][0] +
                mat_A[93][3] * mat_B[190][0] +
                mat_A[94][0] * mat_B[198][0] +
                mat_A[94][1] * mat_B[206][0] +
                mat_A[94][2] * mat_B[214][0] +
                mat_A[94][3] * mat_B[222][0] +
                mat_A[95][0] * mat_B[230][0] +
                mat_A[95][1] * mat_B[238][0] +
                mat_A[95][2] * mat_B[246][0] +
                mat_A[95][3] * mat_B[254][0];
    mat_C[94][1] <=
                mat_A[88][0] * mat_B[6][1] +
                mat_A[88][1] * mat_B[14][1] +
                mat_A[88][2] * mat_B[22][1] +
                mat_A[88][3] * mat_B[30][1] +
                mat_A[89][0] * mat_B[38][1] +
                mat_A[89][1] * mat_B[46][1] +
                mat_A[89][2] * mat_B[54][1] +
                mat_A[89][3] * mat_B[62][1] +
                mat_A[90][0] * mat_B[70][1] +
                mat_A[90][1] * mat_B[78][1] +
                mat_A[90][2] * mat_B[86][1] +
                mat_A[90][3] * mat_B[94][1] +
                mat_A[91][0] * mat_B[102][1] +
                mat_A[91][1] * mat_B[110][1] +
                mat_A[91][2] * mat_B[118][1] +
                mat_A[91][3] * mat_B[126][1] +
                mat_A[92][0] * mat_B[134][1] +
                mat_A[92][1] * mat_B[142][1] +
                mat_A[92][2] * mat_B[150][1] +
                mat_A[92][3] * mat_B[158][1] +
                mat_A[93][0] * mat_B[166][1] +
                mat_A[93][1] * mat_B[174][1] +
                mat_A[93][2] * mat_B[182][1] +
                mat_A[93][3] * mat_B[190][1] +
                mat_A[94][0] * mat_B[198][1] +
                mat_A[94][1] * mat_B[206][1] +
                mat_A[94][2] * mat_B[214][1] +
                mat_A[94][3] * mat_B[222][1] +
                mat_A[95][0] * mat_B[230][1] +
                mat_A[95][1] * mat_B[238][1] +
                mat_A[95][2] * mat_B[246][1] +
                mat_A[95][3] * mat_B[254][1];
    mat_C[94][2] <=
                mat_A[88][0] * mat_B[6][2] +
                mat_A[88][1] * mat_B[14][2] +
                mat_A[88][2] * mat_B[22][2] +
                mat_A[88][3] * mat_B[30][2] +
                mat_A[89][0] * mat_B[38][2] +
                mat_A[89][1] * mat_B[46][2] +
                mat_A[89][2] * mat_B[54][2] +
                mat_A[89][3] * mat_B[62][2] +
                mat_A[90][0] * mat_B[70][2] +
                mat_A[90][1] * mat_B[78][2] +
                mat_A[90][2] * mat_B[86][2] +
                mat_A[90][3] * mat_B[94][2] +
                mat_A[91][0] * mat_B[102][2] +
                mat_A[91][1] * mat_B[110][2] +
                mat_A[91][2] * mat_B[118][2] +
                mat_A[91][3] * mat_B[126][2] +
                mat_A[92][0] * mat_B[134][2] +
                mat_A[92][1] * mat_B[142][2] +
                mat_A[92][2] * mat_B[150][2] +
                mat_A[92][3] * mat_B[158][2] +
                mat_A[93][0] * mat_B[166][2] +
                mat_A[93][1] * mat_B[174][2] +
                mat_A[93][2] * mat_B[182][2] +
                mat_A[93][3] * mat_B[190][2] +
                mat_A[94][0] * mat_B[198][2] +
                mat_A[94][1] * mat_B[206][2] +
                mat_A[94][2] * mat_B[214][2] +
                mat_A[94][3] * mat_B[222][2] +
                mat_A[95][0] * mat_B[230][2] +
                mat_A[95][1] * mat_B[238][2] +
                mat_A[95][2] * mat_B[246][2] +
                mat_A[95][3] * mat_B[254][2];
    mat_C[94][3] <=
                mat_A[88][0] * mat_B[6][3] +
                mat_A[88][1] * mat_B[14][3] +
                mat_A[88][2] * mat_B[22][3] +
                mat_A[88][3] * mat_B[30][3] +
                mat_A[89][0] * mat_B[38][3] +
                mat_A[89][1] * mat_B[46][3] +
                mat_A[89][2] * mat_B[54][3] +
                mat_A[89][3] * mat_B[62][3] +
                mat_A[90][0] * mat_B[70][3] +
                mat_A[90][1] * mat_B[78][3] +
                mat_A[90][2] * mat_B[86][3] +
                mat_A[90][3] * mat_B[94][3] +
                mat_A[91][0] * mat_B[102][3] +
                mat_A[91][1] * mat_B[110][3] +
                mat_A[91][2] * mat_B[118][3] +
                mat_A[91][3] * mat_B[126][3] +
                mat_A[92][0] * mat_B[134][3] +
                mat_A[92][1] * mat_B[142][3] +
                mat_A[92][2] * mat_B[150][3] +
                mat_A[92][3] * mat_B[158][3] +
                mat_A[93][0] * mat_B[166][3] +
                mat_A[93][1] * mat_B[174][3] +
                mat_A[93][2] * mat_B[182][3] +
                mat_A[93][3] * mat_B[190][3] +
                mat_A[94][0] * mat_B[198][3] +
                mat_A[94][1] * mat_B[206][3] +
                mat_A[94][2] * mat_B[214][3] +
                mat_A[94][3] * mat_B[222][3] +
                mat_A[95][0] * mat_B[230][3] +
                mat_A[95][1] * mat_B[238][3] +
                mat_A[95][2] * mat_B[246][3] +
                mat_A[95][3] * mat_B[254][3];
    mat_C[95][0] <=
                mat_A[88][0] * mat_B[7][0] +
                mat_A[88][1] * mat_B[15][0] +
                mat_A[88][2] * mat_B[23][0] +
                mat_A[88][3] * mat_B[31][0] +
                mat_A[89][0] * mat_B[39][0] +
                mat_A[89][1] * mat_B[47][0] +
                mat_A[89][2] * mat_B[55][0] +
                mat_A[89][3] * mat_B[63][0] +
                mat_A[90][0] * mat_B[71][0] +
                mat_A[90][1] * mat_B[79][0] +
                mat_A[90][2] * mat_B[87][0] +
                mat_A[90][3] * mat_B[95][0] +
                mat_A[91][0] * mat_B[103][0] +
                mat_A[91][1] * mat_B[111][0] +
                mat_A[91][2] * mat_B[119][0] +
                mat_A[91][3] * mat_B[127][0] +
                mat_A[92][0] * mat_B[135][0] +
                mat_A[92][1] * mat_B[143][0] +
                mat_A[92][2] * mat_B[151][0] +
                mat_A[92][3] * mat_B[159][0] +
                mat_A[93][0] * mat_B[167][0] +
                mat_A[93][1] * mat_B[175][0] +
                mat_A[93][2] * mat_B[183][0] +
                mat_A[93][3] * mat_B[191][0] +
                mat_A[94][0] * mat_B[199][0] +
                mat_A[94][1] * mat_B[207][0] +
                mat_A[94][2] * mat_B[215][0] +
                mat_A[94][3] * mat_B[223][0] +
                mat_A[95][0] * mat_B[231][0] +
                mat_A[95][1] * mat_B[239][0] +
                mat_A[95][2] * mat_B[247][0] +
                mat_A[95][3] * mat_B[255][0];
    mat_C[95][1] <=
                mat_A[88][0] * mat_B[7][1] +
                mat_A[88][1] * mat_B[15][1] +
                mat_A[88][2] * mat_B[23][1] +
                mat_A[88][3] * mat_B[31][1] +
                mat_A[89][0] * mat_B[39][1] +
                mat_A[89][1] * mat_B[47][1] +
                mat_A[89][2] * mat_B[55][1] +
                mat_A[89][3] * mat_B[63][1] +
                mat_A[90][0] * mat_B[71][1] +
                mat_A[90][1] * mat_B[79][1] +
                mat_A[90][2] * mat_B[87][1] +
                mat_A[90][3] * mat_B[95][1] +
                mat_A[91][0] * mat_B[103][1] +
                mat_A[91][1] * mat_B[111][1] +
                mat_A[91][2] * mat_B[119][1] +
                mat_A[91][3] * mat_B[127][1] +
                mat_A[92][0] * mat_B[135][1] +
                mat_A[92][1] * mat_B[143][1] +
                mat_A[92][2] * mat_B[151][1] +
                mat_A[92][3] * mat_B[159][1] +
                mat_A[93][0] * mat_B[167][1] +
                mat_A[93][1] * mat_B[175][1] +
                mat_A[93][2] * mat_B[183][1] +
                mat_A[93][3] * mat_B[191][1] +
                mat_A[94][0] * mat_B[199][1] +
                mat_A[94][1] * mat_B[207][1] +
                mat_A[94][2] * mat_B[215][1] +
                mat_A[94][3] * mat_B[223][1] +
                mat_A[95][0] * mat_B[231][1] +
                mat_A[95][1] * mat_B[239][1] +
                mat_A[95][2] * mat_B[247][1] +
                mat_A[95][3] * mat_B[255][1];
    mat_C[95][2] <=
                mat_A[88][0] * mat_B[7][2] +
                mat_A[88][1] * mat_B[15][2] +
                mat_A[88][2] * mat_B[23][2] +
                mat_A[88][3] * mat_B[31][2] +
                mat_A[89][0] * mat_B[39][2] +
                mat_A[89][1] * mat_B[47][2] +
                mat_A[89][2] * mat_B[55][2] +
                mat_A[89][3] * mat_B[63][2] +
                mat_A[90][0] * mat_B[71][2] +
                mat_A[90][1] * mat_B[79][2] +
                mat_A[90][2] * mat_B[87][2] +
                mat_A[90][3] * mat_B[95][2] +
                mat_A[91][0] * mat_B[103][2] +
                mat_A[91][1] * mat_B[111][2] +
                mat_A[91][2] * mat_B[119][2] +
                mat_A[91][3] * mat_B[127][2] +
                mat_A[92][0] * mat_B[135][2] +
                mat_A[92][1] * mat_B[143][2] +
                mat_A[92][2] * mat_B[151][2] +
                mat_A[92][3] * mat_B[159][2] +
                mat_A[93][0] * mat_B[167][2] +
                mat_A[93][1] * mat_B[175][2] +
                mat_A[93][2] * mat_B[183][2] +
                mat_A[93][3] * mat_B[191][2] +
                mat_A[94][0] * mat_B[199][2] +
                mat_A[94][1] * mat_B[207][2] +
                mat_A[94][2] * mat_B[215][2] +
                mat_A[94][3] * mat_B[223][2] +
                mat_A[95][0] * mat_B[231][2] +
                mat_A[95][1] * mat_B[239][2] +
                mat_A[95][2] * mat_B[247][2] +
                mat_A[95][3] * mat_B[255][2];
    mat_C[95][3] <=
                mat_A[88][0] * mat_B[7][3] +
                mat_A[88][1] * mat_B[15][3] +
                mat_A[88][2] * mat_B[23][3] +
                mat_A[88][3] * mat_B[31][3] +
                mat_A[89][0] * mat_B[39][3] +
                mat_A[89][1] * mat_B[47][3] +
                mat_A[89][2] * mat_B[55][3] +
                mat_A[89][3] * mat_B[63][3] +
                mat_A[90][0] * mat_B[71][3] +
                mat_A[90][1] * mat_B[79][3] +
                mat_A[90][2] * mat_B[87][3] +
                mat_A[90][3] * mat_B[95][3] +
                mat_A[91][0] * mat_B[103][3] +
                mat_A[91][1] * mat_B[111][3] +
                mat_A[91][2] * mat_B[119][3] +
                mat_A[91][3] * mat_B[127][3] +
                mat_A[92][0] * mat_B[135][3] +
                mat_A[92][1] * mat_B[143][3] +
                mat_A[92][2] * mat_B[151][3] +
                mat_A[92][3] * mat_B[159][3] +
                mat_A[93][0] * mat_B[167][3] +
                mat_A[93][1] * mat_B[175][3] +
                mat_A[93][2] * mat_B[183][3] +
                mat_A[93][3] * mat_B[191][3] +
                mat_A[94][0] * mat_B[199][3] +
                mat_A[94][1] * mat_B[207][3] +
                mat_A[94][2] * mat_B[215][3] +
                mat_A[94][3] * mat_B[223][3] +
                mat_A[95][0] * mat_B[231][3] +
                mat_A[95][1] * mat_B[239][3] +
                mat_A[95][2] * mat_B[247][3] +
                mat_A[95][3] * mat_B[255][3];
    mat_C[96][0] <=
                mat_A[96][0] * mat_B[0][0] +
                mat_A[96][1] * mat_B[8][0] +
                mat_A[96][2] * mat_B[16][0] +
                mat_A[96][3] * mat_B[24][0] +
                mat_A[97][0] * mat_B[32][0] +
                mat_A[97][1] * mat_B[40][0] +
                mat_A[97][2] * mat_B[48][0] +
                mat_A[97][3] * mat_B[56][0] +
                mat_A[98][0] * mat_B[64][0] +
                mat_A[98][1] * mat_B[72][0] +
                mat_A[98][2] * mat_B[80][0] +
                mat_A[98][3] * mat_B[88][0] +
                mat_A[99][0] * mat_B[96][0] +
                mat_A[99][1] * mat_B[104][0] +
                mat_A[99][2] * mat_B[112][0] +
                mat_A[99][3] * mat_B[120][0] +
                mat_A[100][0] * mat_B[128][0] +
                mat_A[100][1] * mat_B[136][0] +
                mat_A[100][2] * mat_B[144][0] +
                mat_A[100][3] * mat_B[152][0] +
                mat_A[101][0] * mat_B[160][0] +
                mat_A[101][1] * mat_B[168][0] +
                mat_A[101][2] * mat_B[176][0] +
                mat_A[101][3] * mat_B[184][0] +
                mat_A[102][0] * mat_B[192][0] +
                mat_A[102][1] * mat_B[200][0] +
                mat_A[102][2] * mat_B[208][0] +
                mat_A[102][3] * mat_B[216][0] +
                mat_A[103][0] * mat_B[224][0] +
                mat_A[103][1] * mat_B[232][0] +
                mat_A[103][2] * mat_B[240][0] +
                mat_A[103][3] * mat_B[248][0];
    mat_C[96][1] <=
                mat_A[96][0] * mat_B[0][1] +
                mat_A[96][1] * mat_B[8][1] +
                mat_A[96][2] * mat_B[16][1] +
                mat_A[96][3] * mat_B[24][1] +
                mat_A[97][0] * mat_B[32][1] +
                mat_A[97][1] * mat_B[40][1] +
                mat_A[97][2] * mat_B[48][1] +
                mat_A[97][3] * mat_B[56][1] +
                mat_A[98][0] * mat_B[64][1] +
                mat_A[98][1] * mat_B[72][1] +
                mat_A[98][2] * mat_B[80][1] +
                mat_A[98][3] * mat_B[88][1] +
                mat_A[99][0] * mat_B[96][1] +
                mat_A[99][1] * mat_B[104][1] +
                mat_A[99][2] * mat_B[112][1] +
                mat_A[99][3] * mat_B[120][1] +
                mat_A[100][0] * mat_B[128][1] +
                mat_A[100][1] * mat_B[136][1] +
                mat_A[100][2] * mat_B[144][1] +
                mat_A[100][3] * mat_B[152][1] +
                mat_A[101][0] * mat_B[160][1] +
                mat_A[101][1] * mat_B[168][1] +
                mat_A[101][2] * mat_B[176][1] +
                mat_A[101][3] * mat_B[184][1] +
                mat_A[102][0] * mat_B[192][1] +
                mat_A[102][1] * mat_B[200][1] +
                mat_A[102][2] * mat_B[208][1] +
                mat_A[102][3] * mat_B[216][1] +
                mat_A[103][0] * mat_B[224][1] +
                mat_A[103][1] * mat_B[232][1] +
                mat_A[103][2] * mat_B[240][1] +
                mat_A[103][3] * mat_B[248][1];
    mat_C[96][2] <=
                mat_A[96][0] * mat_B[0][2] +
                mat_A[96][1] * mat_B[8][2] +
                mat_A[96][2] * mat_B[16][2] +
                mat_A[96][3] * mat_B[24][2] +
                mat_A[97][0] * mat_B[32][2] +
                mat_A[97][1] * mat_B[40][2] +
                mat_A[97][2] * mat_B[48][2] +
                mat_A[97][3] * mat_B[56][2] +
                mat_A[98][0] * mat_B[64][2] +
                mat_A[98][1] * mat_B[72][2] +
                mat_A[98][2] * mat_B[80][2] +
                mat_A[98][3] * mat_B[88][2] +
                mat_A[99][0] * mat_B[96][2] +
                mat_A[99][1] * mat_B[104][2] +
                mat_A[99][2] * mat_B[112][2] +
                mat_A[99][3] * mat_B[120][2] +
                mat_A[100][0] * mat_B[128][2] +
                mat_A[100][1] * mat_B[136][2] +
                mat_A[100][2] * mat_B[144][2] +
                mat_A[100][3] * mat_B[152][2] +
                mat_A[101][0] * mat_B[160][2] +
                mat_A[101][1] * mat_B[168][2] +
                mat_A[101][2] * mat_B[176][2] +
                mat_A[101][3] * mat_B[184][2] +
                mat_A[102][0] * mat_B[192][2] +
                mat_A[102][1] * mat_B[200][2] +
                mat_A[102][2] * mat_B[208][2] +
                mat_A[102][3] * mat_B[216][2] +
                mat_A[103][0] * mat_B[224][2] +
                mat_A[103][1] * mat_B[232][2] +
                mat_A[103][2] * mat_B[240][2] +
                mat_A[103][3] * mat_B[248][2];
    mat_C[96][3] <=
                mat_A[96][0] * mat_B[0][3] +
                mat_A[96][1] * mat_B[8][3] +
                mat_A[96][2] * mat_B[16][3] +
                mat_A[96][3] * mat_B[24][3] +
                mat_A[97][0] * mat_B[32][3] +
                mat_A[97][1] * mat_B[40][3] +
                mat_A[97][2] * mat_B[48][3] +
                mat_A[97][3] * mat_B[56][3] +
                mat_A[98][0] * mat_B[64][3] +
                mat_A[98][1] * mat_B[72][3] +
                mat_A[98][2] * mat_B[80][3] +
                mat_A[98][3] * mat_B[88][3] +
                mat_A[99][0] * mat_B[96][3] +
                mat_A[99][1] * mat_B[104][3] +
                mat_A[99][2] * mat_B[112][3] +
                mat_A[99][3] * mat_B[120][3] +
                mat_A[100][0] * mat_B[128][3] +
                mat_A[100][1] * mat_B[136][3] +
                mat_A[100][2] * mat_B[144][3] +
                mat_A[100][3] * mat_B[152][3] +
                mat_A[101][0] * mat_B[160][3] +
                mat_A[101][1] * mat_B[168][3] +
                mat_A[101][2] * mat_B[176][3] +
                mat_A[101][3] * mat_B[184][3] +
                mat_A[102][0] * mat_B[192][3] +
                mat_A[102][1] * mat_B[200][3] +
                mat_A[102][2] * mat_B[208][3] +
                mat_A[102][3] * mat_B[216][3] +
                mat_A[103][0] * mat_B[224][3] +
                mat_A[103][1] * mat_B[232][3] +
                mat_A[103][2] * mat_B[240][3] +
                mat_A[103][3] * mat_B[248][3];
    mat_C[97][0] <=
                mat_A[96][0] * mat_B[1][0] +
                mat_A[96][1] * mat_B[9][0] +
                mat_A[96][2] * mat_B[17][0] +
                mat_A[96][3] * mat_B[25][0] +
                mat_A[97][0] * mat_B[33][0] +
                mat_A[97][1] * mat_B[41][0] +
                mat_A[97][2] * mat_B[49][0] +
                mat_A[97][3] * mat_B[57][0] +
                mat_A[98][0] * mat_B[65][0] +
                mat_A[98][1] * mat_B[73][0] +
                mat_A[98][2] * mat_B[81][0] +
                mat_A[98][3] * mat_B[89][0] +
                mat_A[99][0] * mat_B[97][0] +
                mat_A[99][1] * mat_B[105][0] +
                mat_A[99][2] * mat_B[113][0] +
                mat_A[99][3] * mat_B[121][0] +
                mat_A[100][0] * mat_B[129][0] +
                mat_A[100][1] * mat_B[137][0] +
                mat_A[100][2] * mat_B[145][0] +
                mat_A[100][3] * mat_B[153][0] +
                mat_A[101][0] * mat_B[161][0] +
                mat_A[101][1] * mat_B[169][0] +
                mat_A[101][2] * mat_B[177][0] +
                mat_A[101][3] * mat_B[185][0] +
                mat_A[102][0] * mat_B[193][0] +
                mat_A[102][1] * mat_B[201][0] +
                mat_A[102][2] * mat_B[209][0] +
                mat_A[102][3] * mat_B[217][0] +
                mat_A[103][0] * mat_B[225][0] +
                mat_A[103][1] * mat_B[233][0] +
                mat_A[103][2] * mat_B[241][0] +
                mat_A[103][3] * mat_B[249][0];
    mat_C[97][1] <=
                mat_A[96][0] * mat_B[1][1] +
                mat_A[96][1] * mat_B[9][1] +
                mat_A[96][2] * mat_B[17][1] +
                mat_A[96][3] * mat_B[25][1] +
                mat_A[97][0] * mat_B[33][1] +
                mat_A[97][1] * mat_B[41][1] +
                mat_A[97][2] * mat_B[49][1] +
                mat_A[97][3] * mat_B[57][1] +
                mat_A[98][0] * mat_B[65][1] +
                mat_A[98][1] * mat_B[73][1] +
                mat_A[98][2] * mat_B[81][1] +
                mat_A[98][3] * mat_B[89][1] +
                mat_A[99][0] * mat_B[97][1] +
                mat_A[99][1] * mat_B[105][1] +
                mat_A[99][2] * mat_B[113][1] +
                mat_A[99][3] * mat_B[121][1] +
                mat_A[100][0] * mat_B[129][1] +
                mat_A[100][1] * mat_B[137][1] +
                mat_A[100][2] * mat_B[145][1] +
                mat_A[100][3] * mat_B[153][1] +
                mat_A[101][0] * mat_B[161][1] +
                mat_A[101][1] * mat_B[169][1] +
                mat_A[101][2] * mat_B[177][1] +
                mat_A[101][3] * mat_B[185][1] +
                mat_A[102][0] * mat_B[193][1] +
                mat_A[102][1] * mat_B[201][1] +
                mat_A[102][2] * mat_B[209][1] +
                mat_A[102][3] * mat_B[217][1] +
                mat_A[103][0] * mat_B[225][1] +
                mat_A[103][1] * mat_B[233][1] +
                mat_A[103][2] * mat_B[241][1] +
                mat_A[103][3] * mat_B[249][1];
    mat_C[97][2] <=
                mat_A[96][0] * mat_B[1][2] +
                mat_A[96][1] * mat_B[9][2] +
                mat_A[96][2] * mat_B[17][2] +
                mat_A[96][3] * mat_B[25][2] +
                mat_A[97][0] * mat_B[33][2] +
                mat_A[97][1] * mat_B[41][2] +
                mat_A[97][2] * mat_B[49][2] +
                mat_A[97][3] * mat_B[57][2] +
                mat_A[98][0] * mat_B[65][2] +
                mat_A[98][1] * mat_B[73][2] +
                mat_A[98][2] * mat_B[81][2] +
                mat_A[98][3] * mat_B[89][2] +
                mat_A[99][0] * mat_B[97][2] +
                mat_A[99][1] * mat_B[105][2] +
                mat_A[99][2] * mat_B[113][2] +
                mat_A[99][3] * mat_B[121][2] +
                mat_A[100][0] * mat_B[129][2] +
                mat_A[100][1] * mat_B[137][2] +
                mat_A[100][2] * mat_B[145][2] +
                mat_A[100][3] * mat_B[153][2] +
                mat_A[101][0] * mat_B[161][2] +
                mat_A[101][1] * mat_B[169][2] +
                mat_A[101][2] * mat_B[177][2] +
                mat_A[101][3] * mat_B[185][2] +
                mat_A[102][0] * mat_B[193][2] +
                mat_A[102][1] * mat_B[201][2] +
                mat_A[102][2] * mat_B[209][2] +
                mat_A[102][3] * mat_B[217][2] +
                mat_A[103][0] * mat_B[225][2] +
                mat_A[103][1] * mat_B[233][2] +
                mat_A[103][2] * mat_B[241][2] +
                mat_A[103][3] * mat_B[249][2];
    mat_C[97][3] <=
                mat_A[96][0] * mat_B[1][3] +
                mat_A[96][1] * mat_B[9][3] +
                mat_A[96][2] * mat_B[17][3] +
                mat_A[96][3] * mat_B[25][3] +
                mat_A[97][0] * mat_B[33][3] +
                mat_A[97][1] * mat_B[41][3] +
                mat_A[97][2] * mat_B[49][3] +
                mat_A[97][3] * mat_B[57][3] +
                mat_A[98][0] * mat_B[65][3] +
                mat_A[98][1] * mat_B[73][3] +
                mat_A[98][2] * mat_B[81][3] +
                mat_A[98][3] * mat_B[89][3] +
                mat_A[99][0] * mat_B[97][3] +
                mat_A[99][1] * mat_B[105][3] +
                mat_A[99][2] * mat_B[113][3] +
                mat_A[99][3] * mat_B[121][3] +
                mat_A[100][0] * mat_B[129][3] +
                mat_A[100][1] * mat_B[137][3] +
                mat_A[100][2] * mat_B[145][3] +
                mat_A[100][3] * mat_B[153][3] +
                mat_A[101][0] * mat_B[161][3] +
                mat_A[101][1] * mat_B[169][3] +
                mat_A[101][2] * mat_B[177][3] +
                mat_A[101][3] * mat_B[185][3] +
                mat_A[102][0] * mat_B[193][3] +
                mat_A[102][1] * mat_B[201][3] +
                mat_A[102][2] * mat_B[209][3] +
                mat_A[102][3] * mat_B[217][3] +
                mat_A[103][0] * mat_B[225][3] +
                mat_A[103][1] * mat_B[233][3] +
                mat_A[103][2] * mat_B[241][3] +
                mat_A[103][3] * mat_B[249][3];
    mat_C[98][0] <=
                mat_A[96][0] * mat_B[2][0] +
                mat_A[96][1] * mat_B[10][0] +
                mat_A[96][2] * mat_B[18][0] +
                mat_A[96][3] * mat_B[26][0] +
                mat_A[97][0] * mat_B[34][0] +
                mat_A[97][1] * mat_B[42][0] +
                mat_A[97][2] * mat_B[50][0] +
                mat_A[97][3] * mat_B[58][0] +
                mat_A[98][0] * mat_B[66][0] +
                mat_A[98][1] * mat_B[74][0] +
                mat_A[98][2] * mat_B[82][0] +
                mat_A[98][3] * mat_B[90][0] +
                mat_A[99][0] * mat_B[98][0] +
                mat_A[99][1] * mat_B[106][0] +
                mat_A[99][2] * mat_B[114][0] +
                mat_A[99][3] * mat_B[122][0] +
                mat_A[100][0] * mat_B[130][0] +
                mat_A[100][1] * mat_B[138][0] +
                mat_A[100][2] * mat_B[146][0] +
                mat_A[100][3] * mat_B[154][0] +
                mat_A[101][0] * mat_B[162][0] +
                mat_A[101][1] * mat_B[170][0] +
                mat_A[101][2] * mat_B[178][0] +
                mat_A[101][3] * mat_B[186][0] +
                mat_A[102][0] * mat_B[194][0] +
                mat_A[102][1] * mat_B[202][0] +
                mat_A[102][2] * mat_B[210][0] +
                mat_A[102][3] * mat_B[218][0] +
                mat_A[103][0] * mat_B[226][0] +
                mat_A[103][1] * mat_B[234][0] +
                mat_A[103][2] * mat_B[242][0] +
                mat_A[103][3] * mat_B[250][0];
    mat_C[98][1] <=
                mat_A[96][0] * mat_B[2][1] +
                mat_A[96][1] * mat_B[10][1] +
                mat_A[96][2] * mat_B[18][1] +
                mat_A[96][3] * mat_B[26][1] +
                mat_A[97][0] * mat_B[34][1] +
                mat_A[97][1] * mat_B[42][1] +
                mat_A[97][2] * mat_B[50][1] +
                mat_A[97][3] * mat_B[58][1] +
                mat_A[98][0] * mat_B[66][1] +
                mat_A[98][1] * mat_B[74][1] +
                mat_A[98][2] * mat_B[82][1] +
                mat_A[98][3] * mat_B[90][1] +
                mat_A[99][0] * mat_B[98][1] +
                mat_A[99][1] * mat_B[106][1] +
                mat_A[99][2] * mat_B[114][1] +
                mat_A[99][3] * mat_B[122][1] +
                mat_A[100][0] * mat_B[130][1] +
                mat_A[100][1] * mat_B[138][1] +
                mat_A[100][2] * mat_B[146][1] +
                mat_A[100][3] * mat_B[154][1] +
                mat_A[101][0] * mat_B[162][1] +
                mat_A[101][1] * mat_B[170][1] +
                mat_A[101][2] * mat_B[178][1] +
                mat_A[101][3] * mat_B[186][1] +
                mat_A[102][0] * mat_B[194][1] +
                mat_A[102][1] * mat_B[202][1] +
                mat_A[102][2] * mat_B[210][1] +
                mat_A[102][3] * mat_B[218][1] +
                mat_A[103][0] * mat_B[226][1] +
                mat_A[103][1] * mat_B[234][1] +
                mat_A[103][2] * mat_B[242][1] +
                mat_A[103][3] * mat_B[250][1];
    mat_C[98][2] <=
                mat_A[96][0] * mat_B[2][2] +
                mat_A[96][1] * mat_B[10][2] +
                mat_A[96][2] * mat_B[18][2] +
                mat_A[96][3] * mat_B[26][2] +
                mat_A[97][0] * mat_B[34][2] +
                mat_A[97][1] * mat_B[42][2] +
                mat_A[97][2] * mat_B[50][2] +
                mat_A[97][3] * mat_B[58][2] +
                mat_A[98][0] * mat_B[66][2] +
                mat_A[98][1] * mat_B[74][2] +
                mat_A[98][2] * mat_B[82][2] +
                mat_A[98][3] * mat_B[90][2] +
                mat_A[99][0] * mat_B[98][2] +
                mat_A[99][1] * mat_B[106][2] +
                mat_A[99][2] * mat_B[114][2] +
                mat_A[99][3] * mat_B[122][2] +
                mat_A[100][0] * mat_B[130][2] +
                mat_A[100][1] * mat_B[138][2] +
                mat_A[100][2] * mat_B[146][2] +
                mat_A[100][3] * mat_B[154][2] +
                mat_A[101][0] * mat_B[162][2] +
                mat_A[101][1] * mat_B[170][2] +
                mat_A[101][2] * mat_B[178][2] +
                mat_A[101][3] * mat_B[186][2] +
                mat_A[102][0] * mat_B[194][2] +
                mat_A[102][1] * mat_B[202][2] +
                mat_A[102][2] * mat_B[210][2] +
                mat_A[102][3] * mat_B[218][2] +
                mat_A[103][0] * mat_B[226][2] +
                mat_A[103][1] * mat_B[234][2] +
                mat_A[103][2] * mat_B[242][2] +
                mat_A[103][3] * mat_B[250][2];
    mat_C[98][3] <=
                mat_A[96][0] * mat_B[2][3] +
                mat_A[96][1] * mat_B[10][3] +
                mat_A[96][2] * mat_B[18][3] +
                mat_A[96][3] * mat_B[26][3] +
                mat_A[97][0] * mat_B[34][3] +
                mat_A[97][1] * mat_B[42][3] +
                mat_A[97][2] * mat_B[50][3] +
                mat_A[97][3] * mat_B[58][3] +
                mat_A[98][0] * mat_B[66][3] +
                mat_A[98][1] * mat_B[74][3] +
                mat_A[98][2] * mat_B[82][3] +
                mat_A[98][3] * mat_B[90][3] +
                mat_A[99][0] * mat_B[98][3] +
                mat_A[99][1] * mat_B[106][3] +
                mat_A[99][2] * mat_B[114][3] +
                mat_A[99][3] * mat_B[122][3] +
                mat_A[100][0] * mat_B[130][3] +
                mat_A[100][1] * mat_B[138][3] +
                mat_A[100][2] * mat_B[146][3] +
                mat_A[100][3] * mat_B[154][3] +
                mat_A[101][0] * mat_B[162][3] +
                mat_A[101][1] * mat_B[170][3] +
                mat_A[101][2] * mat_B[178][3] +
                mat_A[101][3] * mat_B[186][3] +
                mat_A[102][0] * mat_B[194][3] +
                mat_A[102][1] * mat_B[202][3] +
                mat_A[102][2] * mat_B[210][3] +
                mat_A[102][3] * mat_B[218][3] +
                mat_A[103][0] * mat_B[226][3] +
                mat_A[103][1] * mat_B[234][3] +
                mat_A[103][2] * mat_B[242][3] +
                mat_A[103][3] * mat_B[250][3];
    mat_C[99][0] <=
                mat_A[96][0] * mat_B[3][0] +
                mat_A[96][1] * mat_B[11][0] +
                mat_A[96][2] * mat_B[19][0] +
                mat_A[96][3] * mat_B[27][0] +
                mat_A[97][0] * mat_B[35][0] +
                mat_A[97][1] * mat_B[43][0] +
                mat_A[97][2] * mat_B[51][0] +
                mat_A[97][3] * mat_B[59][0] +
                mat_A[98][0] * mat_B[67][0] +
                mat_A[98][1] * mat_B[75][0] +
                mat_A[98][2] * mat_B[83][0] +
                mat_A[98][3] * mat_B[91][0] +
                mat_A[99][0] * mat_B[99][0] +
                mat_A[99][1] * mat_B[107][0] +
                mat_A[99][2] * mat_B[115][0] +
                mat_A[99][3] * mat_B[123][0] +
                mat_A[100][0] * mat_B[131][0] +
                mat_A[100][1] * mat_B[139][0] +
                mat_A[100][2] * mat_B[147][0] +
                mat_A[100][3] * mat_B[155][0] +
                mat_A[101][0] * mat_B[163][0] +
                mat_A[101][1] * mat_B[171][0] +
                mat_A[101][2] * mat_B[179][0] +
                mat_A[101][3] * mat_B[187][0] +
                mat_A[102][0] * mat_B[195][0] +
                mat_A[102][1] * mat_B[203][0] +
                mat_A[102][2] * mat_B[211][0] +
                mat_A[102][3] * mat_B[219][0] +
                mat_A[103][0] * mat_B[227][0] +
                mat_A[103][1] * mat_B[235][0] +
                mat_A[103][2] * mat_B[243][0] +
                mat_A[103][3] * mat_B[251][0];
    mat_C[99][1] <=
                mat_A[96][0] * mat_B[3][1] +
                mat_A[96][1] * mat_B[11][1] +
                mat_A[96][2] * mat_B[19][1] +
                mat_A[96][3] * mat_B[27][1] +
                mat_A[97][0] * mat_B[35][1] +
                mat_A[97][1] * mat_B[43][1] +
                mat_A[97][2] * mat_B[51][1] +
                mat_A[97][3] * mat_B[59][1] +
                mat_A[98][0] * mat_B[67][1] +
                mat_A[98][1] * mat_B[75][1] +
                mat_A[98][2] * mat_B[83][1] +
                mat_A[98][3] * mat_B[91][1] +
                mat_A[99][0] * mat_B[99][1] +
                mat_A[99][1] * mat_B[107][1] +
                mat_A[99][2] * mat_B[115][1] +
                mat_A[99][3] * mat_B[123][1] +
                mat_A[100][0] * mat_B[131][1] +
                mat_A[100][1] * mat_B[139][1] +
                mat_A[100][2] * mat_B[147][1] +
                mat_A[100][3] * mat_B[155][1] +
                mat_A[101][0] * mat_B[163][1] +
                mat_A[101][1] * mat_B[171][1] +
                mat_A[101][2] * mat_B[179][1] +
                mat_A[101][3] * mat_B[187][1] +
                mat_A[102][0] * mat_B[195][1] +
                mat_A[102][1] * mat_B[203][1] +
                mat_A[102][2] * mat_B[211][1] +
                mat_A[102][3] * mat_B[219][1] +
                mat_A[103][0] * mat_B[227][1] +
                mat_A[103][1] * mat_B[235][1] +
                mat_A[103][2] * mat_B[243][1] +
                mat_A[103][3] * mat_B[251][1];
    mat_C[99][2] <=
                mat_A[96][0] * mat_B[3][2] +
                mat_A[96][1] * mat_B[11][2] +
                mat_A[96][2] * mat_B[19][2] +
                mat_A[96][3] * mat_B[27][2] +
                mat_A[97][0] * mat_B[35][2] +
                mat_A[97][1] * mat_B[43][2] +
                mat_A[97][2] * mat_B[51][2] +
                mat_A[97][3] * mat_B[59][2] +
                mat_A[98][0] * mat_B[67][2] +
                mat_A[98][1] * mat_B[75][2] +
                mat_A[98][2] * mat_B[83][2] +
                mat_A[98][3] * mat_B[91][2] +
                mat_A[99][0] * mat_B[99][2] +
                mat_A[99][1] * mat_B[107][2] +
                mat_A[99][2] * mat_B[115][2] +
                mat_A[99][3] * mat_B[123][2] +
                mat_A[100][0] * mat_B[131][2] +
                mat_A[100][1] * mat_B[139][2] +
                mat_A[100][2] * mat_B[147][2] +
                mat_A[100][3] * mat_B[155][2] +
                mat_A[101][0] * mat_B[163][2] +
                mat_A[101][1] * mat_B[171][2] +
                mat_A[101][2] * mat_B[179][2] +
                mat_A[101][3] * mat_B[187][2] +
                mat_A[102][0] * mat_B[195][2] +
                mat_A[102][1] * mat_B[203][2] +
                mat_A[102][2] * mat_B[211][2] +
                mat_A[102][3] * mat_B[219][2] +
                mat_A[103][0] * mat_B[227][2] +
                mat_A[103][1] * mat_B[235][2] +
                mat_A[103][2] * mat_B[243][2] +
                mat_A[103][3] * mat_B[251][2];
    mat_C[99][3] <=
                mat_A[96][0] * mat_B[3][3] +
                mat_A[96][1] * mat_B[11][3] +
                mat_A[96][2] * mat_B[19][3] +
                mat_A[96][3] * mat_B[27][3] +
                mat_A[97][0] * mat_B[35][3] +
                mat_A[97][1] * mat_B[43][3] +
                mat_A[97][2] * mat_B[51][3] +
                mat_A[97][3] * mat_B[59][3] +
                mat_A[98][0] * mat_B[67][3] +
                mat_A[98][1] * mat_B[75][3] +
                mat_A[98][2] * mat_B[83][3] +
                mat_A[98][3] * mat_B[91][3] +
                mat_A[99][0] * mat_B[99][3] +
                mat_A[99][1] * mat_B[107][3] +
                mat_A[99][2] * mat_B[115][3] +
                mat_A[99][3] * mat_B[123][3] +
                mat_A[100][0] * mat_B[131][3] +
                mat_A[100][1] * mat_B[139][3] +
                mat_A[100][2] * mat_B[147][3] +
                mat_A[100][3] * mat_B[155][3] +
                mat_A[101][0] * mat_B[163][3] +
                mat_A[101][1] * mat_B[171][3] +
                mat_A[101][2] * mat_B[179][3] +
                mat_A[101][3] * mat_B[187][3] +
                mat_A[102][0] * mat_B[195][3] +
                mat_A[102][1] * mat_B[203][3] +
                mat_A[102][2] * mat_B[211][3] +
                mat_A[102][3] * mat_B[219][3] +
                mat_A[103][0] * mat_B[227][3] +
                mat_A[103][1] * mat_B[235][3] +
                mat_A[103][2] * mat_B[243][3] +
                mat_A[103][3] * mat_B[251][3];
    mat_C[100][0] <=
                mat_A[96][0] * mat_B[4][0] +
                mat_A[96][1] * mat_B[12][0] +
                mat_A[96][2] * mat_B[20][0] +
                mat_A[96][3] * mat_B[28][0] +
                mat_A[97][0] * mat_B[36][0] +
                mat_A[97][1] * mat_B[44][0] +
                mat_A[97][2] * mat_B[52][0] +
                mat_A[97][3] * mat_B[60][0] +
                mat_A[98][0] * mat_B[68][0] +
                mat_A[98][1] * mat_B[76][0] +
                mat_A[98][2] * mat_B[84][0] +
                mat_A[98][3] * mat_B[92][0] +
                mat_A[99][0] * mat_B[100][0] +
                mat_A[99][1] * mat_B[108][0] +
                mat_A[99][2] * mat_B[116][0] +
                mat_A[99][3] * mat_B[124][0] +
                mat_A[100][0] * mat_B[132][0] +
                mat_A[100][1] * mat_B[140][0] +
                mat_A[100][2] * mat_B[148][0] +
                mat_A[100][3] * mat_B[156][0] +
                mat_A[101][0] * mat_B[164][0] +
                mat_A[101][1] * mat_B[172][0] +
                mat_A[101][2] * mat_B[180][0] +
                mat_A[101][3] * mat_B[188][0] +
                mat_A[102][0] * mat_B[196][0] +
                mat_A[102][1] * mat_B[204][0] +
                mat_A[102][2] * mat_B[212][0] +
                mat_A[102][3] * mat_B[220][0] +
                mat_A[103][0] * mat_B[228][0] +
                mat_A[103][1] * mat_B[236][0] +
                mat_A[103][2] * mat_B[244][0] +
                mat_A[103][3] * mat_B[252][0];
    mat_C[100][1] <=
                mat_A[96][0] * mat_B[4][1] +
                mat_A[96][1] * mat_B[12][1] +
                mat_A[96][2] * mat_B[20][1] +
                mat_A[96][3] * mat_B[28][1] +
                mat_A[97][0] * mat_B[36][1] +
                mat_A[97][1] * mat_B[44][1] +
                mat_A[97][2] * mat_B[52][1] +
                mat_A[97][3] * mat_B[60][1] +
                mat_A[98][0] * mat_B[68][1] +
                mat_A[98][1] * mat_B[76][1] +
                mat_A[98][2] * mat_B[84][1] +
                mat_A[98][3] * mat_B[92][1] +
                mat_A[99][0] * mat_B[100][1] +
                mat_A[99][1] * mat_B[108][1] +
                mat_A[99][2] * mat_B[116][1] +
                mat_A[99][3] * mat_B[124][1] +
                mat_A[100][0] * mat_B[132][1] +
                mat_A[100][1] * mat_B[140][1] +
                mat_A[100][2] * mat_B[148][1] +
                mat_A[100][3] * mat_B[156][1] +
                mat_A[101][0] * mat_B[164][1] +
                mat_A[101][1] * mat_B[172][1] +
                mat_A[101][2] * mat_B[180][1] +
                mat_A[101][3] * mat_B[188][1] +
                mat_A[102][0] * mat_B[196][1] +
                mat_A[102][1] * mat_B[204][1] +
                mat_A[102][2] * mat_B[212][1] +
                mat_A[102][3] * mat_B[220][1] +
                mat_A[103][0] * mat_B[228][1] +
                mat_A[103][1] * mat_B[236][1] +
                mat_A[103][2] * mat_B[244][1] +
                mat_A[103][3] * mat_B[252][1];
    mat_C[100][2] <=
                mat_A[96][0] * mat_B[4][2] +
                mat_A[96][1] * mat_B[12][2] +
                mat_A[96][2] * mat_B[20][2] +
                mat_A[96][3] * mat_B[28][2] +
                mat_A[97][0] * mat_B[36][2] +
                mat_A[97][1] * mat_B[44][2] +
                mat_A[97][2] * mat_B[52][2] +
                mat_A[97][3] * mat_B[60][2] +
                mat_A[98][0] * mat_B[68][2] +
                mat_A[98][1] * mat_B[76][2] +
                mat_A[98][2] * mat_B[84][2] +
                mat_A[98][3] * mat_B[92][2] +
                mat_A[99][0] * mat_B[100][2] +
                mat_A[99][1] * mat_B[108][2] +
                mat_A[99][2] * mat_B[116][2] +
                mat_A[99][3] * mat_B[124][2] +
                mat_A[100][0] * mat_B[132][2] +
                mat_A[100][1] * mat_B[140][2] +
                mat_A[100][2] * mat_B[148][2] +
                mat_A[100][3] * mat_B[156][2] +
                mat_A[101][0] * mat_B[164][2] +
                mat_A[101][1] * mat_B[172][2] +
                mat_A[101][2] * mat_B[180][2] +
                mat_A[101][3] * mat_B[188][2] +
                mat_A[102][0] * mat_B[196][2] +
                mat_A[102][1] * mat_B[204][2] +
                mat_A[102][2] * mat_B[212][2] +
                mat_A[102][3] * mat_B[220][2] +
                mat_A[103][0] * mat_B[228][2] +
                mat_A[103][1] * mat_B[236][2] +
                mat_A[103][2] * mat_B[244][2] +
                mat_A[103][3] * mat_B[252][2];
    mat_C[100][3] <=
                mat_A[96][0] * mat_B[4][3] +
                mat_A[96][1] * mat_B[12][3] +
                mat_A[96][2] * mat_B[20][3] +
                mat_A[96][3] * mat_B[28][3] +
                mat_A[97][0] * mat_B[36][3] +
                mat_A[97][1] * mat_B[44][3] +
                mat_A[97][2] * mat_B[52][3] +
                mat_A[97][3] * mat_B[60][3] +
                mat_A[98][0] * mat_B[68][3] +
                mat_A[98][1] * mat_B[76][3] +
                mat_A[98][2] * mat_B[84][3] +
                mat_A[98][3] * mat_B[92][3] +
                mat_A[99][0] * mat_B[100][3] +
                mat_A[99][1] * mat_B[108][3] +
                mat_A[99][2] * mat_B[116][3] +
                mat_A[99][3] * mat_B[124][3] +
                mat_A[100][0] * mat_B[132][3] +
                mat_A[100][1] * mat_B[140][3] +
                mat_A[100][2] * mat_B[148][3] +
                mat_A[100][3] * mat_B[156][3] +
                mat_A[101][0] * mat_B[164][3] +
                mat_A[101][1] * mat_B[172][3] +
                mat_A[101][2] * mat_B[180][3] +
                mat_A[101][3] * mat_B[188][3] +
                mat_A[102][0] * mat_B[196][3] +
                mat_A[102][1] * mat_B[204][3] +
                mat_A[102][2] * mat_B[212][3] +
                mat_A[102][3] * mat_B[220][3] +
                mat_A[103][0] * mat_B[228][3] +
                mat_A[103][1] * mat_B[236][3] +
                mat_A[103][2] * mat_B[244][3] +
                mat_A[103][3] * mat_B[252][3];
    mat_C[101][0] <=
                mat_A[96][0] * mat_B[5][0] +
                mat_A[96][1] * mat_B[13][0] +
                mat_A[96][2] * mat_B[21][0] +
                mat_A[96][3] * mat_B[29][0] +
                mat_A[97][0] * mat_B[37][0] +
                mat_A[97][1] * mat_B[45][0] +
                mat_A[97][2] * mat_B[53][0] +
                mat_A[97][3] * mat_B[61][0] +
                mat_A[98][0] * mat_B[69][0] +
                mat_A[98][1] * mat_B[77][0] +
                mat_A[98][2] * mat_B[85][0] +
                mat_A[98][3] * mat_B[93][0] +
                mat_A[99][0] * mat_B[101][0] +
                mat_A[99][1] * mat_B[109][0] +
                mat_A[99][2] * mat_B[117][0] +
                mat_A[99][3] * mat_B[125][0] +
                mat_A[100][0] * mat_B[133][0] +
                mat_A[100][1] * mat_B[141][0] +
                mat_A[100][2] * mat_B[149][0] +
                mat_A[100][3] * mat_B[157][0] +
                mat_A[101][0] * mat_B[165][0] +
                mat_A[101][1] * mat_B[173][0] +
                mat_A[101][2] * mat_B[181][0] +
                mat_A[101][3] * mat_B[189][0] +
                mat_A[102][0] * mat_B[197][0] +
                mat_A[102][1] * mat_B[205][0] +
                mat_A[102][2] * mat_B[213][0] +
                mat_A[102][3] * mat_B[221][0] +
                mat_A[103][0] * mat_B[229][0] +
                mat_A[103][1] * mat_B[237][0] +
                mat_A[103][2] * mat_B[245][0] +
                mat_A[103][3] * mat_B[253][0];
    mat_C[101][1] <=
                mat_A[96][0] * mat_B[5][1] +
                mat_A[96][1] * mat_B[13][1] +
                mat_A[96][2] * mat_B[21][1] +
                mat_A[96][3] * mat_B[29][1] +
                mat_A[97][0] * mat_B[37][1] +
                mat_A[97][1] * mat_B[45][1] +
                mat_A[97][2] * mat_B[53][1] +
                mat_A[97][3] * mat_B[61][1] +
                mat_A[98][0] * mat_B[69][1] +
                mat_A[98][1] * mat_B[77][1] +
                mat_A[98][2] * mat_B[85][1] +
                mat_A[98][3] * mat_B[93][1] +
                mat_A[99][0] * mat_B[101][1] +
                mat_A[99][1] * mat_B[109][1] +
                mat_A[99][2] * mat_B[117][1] +
                mat_A[99][3] * mat_B[125][1] +
                mat_A[100][0] * mat_B[133][1] +
                mat_A[100][1] * mat_B[141][1] +
                mat_A[100][2] * mat_B[149][1] +
                mat_A[100][3] * mat_B[157][1] +
                mat_A[101][0] * mat_B[165][1] +
                mat_A[101][1] * mat_B[173][1] +
                mat_A[101][2] * mat_B[181][1] +
                mat_A[101][3] * mat_B[189][1] +
                mat_A[102][0] * mat_B[197][1] +
                mat_A[102][1] * mat_B[205][1] +
                mat_A[102][2] * mat_B[213][1] +
                mat_A[102][3] * mat_B[221][1] +
                mat_A[103][0] * mat_B[229][1] +
                mat_A[103][1] * mat_B[237][1] +
                mat_A[103][2] * mat_B[245][1] +
                mat_A[103][3] * mat_B[253][1];
    mat_C[101][2] <=
                mat_A[96][0] * mat_B[5][2] +
                mat_A[96][1] * mat_B[13][2] +
                mat_A[96][2] * mat_B[21][2] +
                mat_A[96][3] * mat_B[29][2] +
                mat_A[97][0] * mat_B[37][2] +
                mat_A[97][1] * mat_B[45][2] +
                mat_A[97][2] * mat_B[53][2] +
                mat_A[97][3] * mat_B[61][2] +
                mat_A[98][0] * mat_B[69][2] +
                mat_A[98][1] * mat_B[77][2] +
                mat_A[98][2] * mat_B[85][2] +
                mat_A[98][3] * mat_B[93][2] +
                mat_A[99][0] * mat_B[101][2] +
                mat_A[99][1] * mat_B[109][2] +
                mat_A[99][2] * mat_B[117][2] +
                mat_A[99][3] * mat_B[125][2] +
                mat_A[100][0] * mat_B[133][2] +
                mat_A[100][1] * mat_B[141][2] +
                mat_A[100][2] * mat_B[149][2] +
                mat_A[100][3] * mat_B[157][2] +
                mat_A[101][0] * mat_B[165][2] +
                mat_A[101][1] * mat_B[173][2] +
                mat_A[101][2] * mat_B[181][2] +
                mat_A[101][3] * mat_B[189][2] +
                mat_A[102][0] * mat_B[197][2] +
                mat_A[102][1] * mat_B[205][2] +
                mat_A[102][2] * mat_B[213][2] +
                mat_A[102][3] * mat_B[221][2] +
                mat_A[103][0] * mat_B[229][2] +
                mat_A[103][1] * mat_B[237][2] +
                mat_A[103][2] * mat_B[245][2] +
                mat_A[103][3] * mat_B[253][2];
    mat_C[101][3] <=
                mat_A[96][0] * mat_B[5][3] +
                mat_A[96][1] * mat_B[13][3] +
                mat_A[96][2] * mat_B[21][3] +
                mat_A[96][3] * mat_B[29][3] +
                mat_A[97][0] * mat_B[37][3] +
                mat_A[97][1] * mat_B[45][3] +
                mat_A[97][2] * mat_B[53][3] +
                mat_A[97][3] * mat_B[61][3] +
                mat_A[98][0] * mat_B[69][3] +
                mat_A[98][1] * mat_B[77][3] +
                mat_A[98][2] * mat_B[85][3] +
                mat_A[98][3] * mat_B[93][3] +
                mat_A[99][0] * mat_B[101][3] +
                mat_A[99][1] * mat_B[109][3] +
                mat_A[99][2] * mat_B[117][3] +
                mat_A[99][3] * mat_B[125][3] +
                mat_A[100][0] * mat_B[133][3] +
                mat_A[100][1] * mat_B[141][3] +
                mat_A[100][2] * mat_B[149][3] +
                mat_A[100][3] * mat_B[157][3] +
                mat_A[101][0] * mat_B[165][3] +
                mat_A[101][1] * mat_B[173][3] +
                mat_A[101][2] * mat_B[181][3] +
                mat_A[101][3] * mat_B[189][3] +
                mat_A[102][0] * mat_B[197][3] +
                mat_A[102][1] * mat_B[205][3] +
                mat_A[102][2] * mat_B[213][3] +
                mat_A[102][3] * mat_B[221][3] +
                mat_A[103][0] * mat_B[229][3] +
                mat_A[103][1] * mat_B[237][3] +
                mat_A[103][2] * mat_B[245][3] +
                mat_A[103][3] * mat_B[253][3];
    mat_C[102][0] <=
                mat_A[96][0] * mat_B[6][0] +
                mat_A[96][1] * mat_B[14][0] +
                mat_A[96][2] * mat_B[22][0] +
                mat_A[96][3] * mat_B[30][0] +
                mat_A[97][0] * mat_B[38][0] +
                mat_A[97][1] * mat_B[46][0] +
                mat_A[97][2] * mat_B[54][0] +
                mat_A[97][3] * mat_B[62][0] +
                mat_A[98][0] * mat_B[70][0] +
                mat_A[98][1] * mat_B[78][0] +
                mat_A[98][2] * mat_B[86][0] +
                mat_A[98][3] * mat_B[94][0] +
                mat_A[99][0] * mat_B[102][0] +
                mat_A[99][1] * mat_B[110][0] +
                mat_A[99][2] * mat_B[118][0] +
                mat_A[99][3] * mat_B[126][0] +
                mat_A[100][0] * mat_B[134][0] +
                mat_A[100][1] * mat_B[142][0] +
                mat_A[100][2] * mat_B[150][0] +
                mat_A[100][3] * mat_B[158][0] +
                mat_A[101][0] * mat_B[166][0] +
                mat_A[101][1] * mat_B[174][0] +
                mat_A[101][2] * mat_B[182][0] +
                mat_A[101][3] * mat_B[190][0] +
                mat_A[102][0] * mat_B[198][0] +
                mat_A[102][1] * mat_B[206][0] +
                mat_A[102][2] * mat_B[214][0] +
                mat_A[102][3] * mat_B[222][0] +
                mat_A[103][0] * mat_B[230][0] +
                mat_A[103][1] * mat_B[238][0] +
                mat_A[103][2] * mat_B[246][0] +
                mat_A[103][3] * mat_B[254][0];
    mat_C[102][1] <=
                mat_A[96][0] * mat_B[6][1] +
                mat_A[96][1] * mat_B[14][1] +
                mat_A[96][2] * mat_B[22][1] +
                mat_A[96][3] * mat_B[30][1] +
                mat_A[97][0] * mat_B[38][1] +
                mat_A[97][1] * mat_B[46][1] +
                mat_A[97][2] * mat_B[54][1] +
                mat_A[97][3] * mat_B[62][1] +
                mat_A[98][0] * mat_B[70][1] +
                mat_A[98][1] * mat_B[78][1] +
                mat_A[98][2] * mat_B[86][1] +
                mat_A[98][3] * mat_B[94][1] +
                mat_A[99][0] * mat_B[102][1] +
                mat_A[99][1] * mat_B[110][1] +
                mat_A[99][2] * mat_B[118][1] +
                mat_A[99][3] * mat_B[126][1] +
                mat_A[100][0] * mat_B[134][1] +
                mat_A[100][1] * mat_B[142][1] +
                mat_A[100][2] * mat_B[150][1] +
                mat_A[100][3] * mat_B[158][1] +
                mat_A[101][0] * mat_B[166][1] +
                mat_A[101][1] * mat_B[174][1] +
                mat_A[101][2] * mat_B[182][1] +
                mat_A[101][3] * mat_B[190][1] +
                mat_A[102][0] * mat_B[198][1] +
                mat_A[102][1] * mat_B[206][1] +
                mat_A[102][2] * mat_B[214][1] +
                mat_A[102][3] * mat_B[222][1] +
                mat_A[103][0] * mat_B[230][1] +
                mat_A[103][1] * mat_B[238][1] +
                mat_A[103][2] * mat_B[246][1] +
                mat_A[103][3] * mat_B[254][1];
    mat_C[102][2] <=
                mat_A[96][0] * mat_B[6][2] +
                mat_A[96][1] * mat_B[14][2] +
                mat_A[96][2] * mat_B[22][2] +
                mat_A[96][3] * mat_B[30][2] +
                mat_A[97][0] * mat_B[38][2] +
                mat_A[97][1] * mat_B[46][2] +
                mat_A[97][2] * mat_B[54][2] +
                mat_A[97][3] * mat_B[62][2] +
                mat_A[98][0] * mat_B[70][2] +
                mat_A[98][1] * mat_B[78][2] +
                mat_A[98][2] * mat_B[86][2] +
                mat_A[98][3] * mat_B[94][2] +
                mat_A[99][0] * mat_B[102][2] +
                mat_A[99][1] * mat_B[110][2] +
                mat_A[99][2] * mat_B[118][2] +
                mat_A[99][3] * mat_B[126][2] +
                mat_A[100][0] * mat_B[134][2] +
                mat_A[100][1] * mat_B[142][2] +
                mat_A[100][2] * mat_B[150][2] +
                mat_A[100][3] * mat_B[158][2] +
                mat_A[101][0] * mat_B[166][2] +
                mat_A[101][1] * mat_B[174][2] +
                mat_A[101][2] * mat_B[182][2] +
                mat_A[101][3] * mat_B[190][2] +
                mat_A[102][0] * mat_B[198][2] +
                mat_A[102][1] * mat_B[206][2] +
                mat_A[102][2] * mat_B[214][2] +
                mat_A[102][3] * mat_B[222][2] +
                mat_A[103][0] * mat_B[230][2] +
                mat_A[103][1] * mat_B[238][2] +
                mat_A[103][2] * mat_B[246][2] +
                mat_A[103][3] * mat_B[254][2];
    mat_C[102][3] <=
                mat_A[96][0] * mat_B[6][3] +
                mat_A[96][1] * mat_B[14][3] +
                mat_A[96][2] * mat_B[22][3] +
                mat_A[96][3] * mat_B[30][3] +
                mat_A[97][0] * mat_B[38][3] +
                mat_A[97][1] * mat_B[46][3] +
                mat_A[97][2] * mat_B[54][3] +
                mat_A[97][3] * mat_B[62][3] +
                mat_A[98][0] * mat_B[70][3] +
                mat_A[98][1] * mat_B[78][3] +
                mat_A[98][2] * mat_B[86][3] +
                mat_A[98][3] * mat_B[94][3] +
                mat_A[99][0] * mat_B[102][3] +
                mat_A[99][1] * mat_B[110][3] +
                mat_A[99][2] * mat_B[118][3] +
                mat_A[99][3] * mat_B[126][3] +
                mat_A[100][0] * mat_B[134][3] +
                mat_A[100][1] * mat_B[142][3] +
                mat_A[100][2] * mat_B[150][3] +
                mat_A[100][3] * mat_B[158][3] +
                mat_A[101][0] * mat_B[166][3] +
                mat_A[101][1] * mat_B[174][3] +
                mat_A[101][2] * mat_B[182][3] +
                mat_A[101][3] * mat_B[190][3] +
                mat_A[102][0] * mat_B[198][3] +
                mat_A[102][1] * mat_B[206][3] +
                mat_A[102][2] * mat_B[214][3] +
                mat_A[102][3] * mat_B[222][3] +
                mat_A[103][0] * mat_B[230][3] +
                mat_A[103][1] * mat_B[238][3] +
                mat_A[103][2] * mat_B[246][3] +
                mat_A[103][3] * mat_B[254][3];
    mat_C[103][0] <=
                mat_A[96][0] * mat_B[7][0] +
                mat_A[96][1] * mat_B[15][0] +
                mat_A[96][2] * mat_B[23][0] +
                mat_A[96][3] * mat_B[31][0] +
                mat_A[97][0] * mat_B[39][0] +
                mat_A[97][1] * mat_B[47][0] +
                mat_A[97][2] * mat_B[55][0] +
                mat_A[97][3] * mat_B[63][0] +
                mat_A[98][0] * mat_B[71][0] +
                mat_A[98][1] * mat_B[79][0] +
                mat_A[98][2] * mat_B[87][0] +
                mat_A[98][3] * mat_B[95][0] +
                mat_A[99][0] * mat_B[103][0] +
                mat_A[99][1] * mat_B[111][0] +
                mat_A[99][2] * mat_B[119][0] +
                mat_A[99][3] * mat_B[127][0] +
                mat_A[100][0] * mat_B[135][0] +
                mat_A[100][1] * mat_B[143][0] +
                mat_A[100][2] * mat_B[151][0] +
                mat_A[100][3] * mat_B[159][0] +
                mat_A[101][0] * mat_B[167][0] +
                mat_A[101][1] * mat_B[175][0] +
                mat_A[101][2] * mat_B[183][0] +
                mat_A[101][3] * mat_B[191][0] +
                mat_A[102][0] * mat_B[199][0] +
                mat_A[102][1] * mat_B[207][0] +
                mat_A[102][2] * mat_B[215][0] +
                mat_A[102][3] * mat_B[223][0] +
                mat_A[103][0] * mat_B[231][0] +
                mat_A[103][1] * mat_B[239][0] +
                mat_A[103][2] * mat_B[247][0] +
                mat_A[103][3] * mat_B[255][0];
    mat_C[103][1] <=
                mat_A[96][0] * mat_B[7][1] +
                mat_A[96][1] * mat_B[15][1] +
                mat_A[96][2] * mat_B[23][1] +
                mat_A[96][3] * mat_B[31][1] +
                mat_A[97][0] * mat_B[39][1] +
                mat_A[97][1] * mat_B[47][1] +
                mat_A[97][2] * mat_B[55][1] +
                mat_A[97][3] * mat_B[63][1] +
                mat_A[98][0] * mat_B[71][1] +
                mat_A[98][1] * mat_B[79][1] +
                mat_A[98][2] * mat_B[87][1] +
                mat_A[98][3] * mat_B[95][1] +
                mat_A[99][0] * mat_B[103][1] +
                mat_A[99][1] * mat_B[111][1] +
                mat_A[99][2] * mat_B[119][1] +
                mat_A[99][3] * mat_B[127][1] +
                mat_A[100][0] * mat_B[135][1] +
                mat_A[100][1] * mat_B[143][1] +
                mat_A[100][2] * mat_B[151][1] +
                mat_A[100][3] * mat_B[159][1] +
                mat_A[101][0] * mat_B[167][1] +
                mat_A[101][1] * mat_B[175][1] +
                mat_A[101][2] * mat_B[183][1] +
                mat_A[101][3] * mat_B[191][1] +
                mat_A[102][0] * mat_B[199][1] +
                mat_A[102][1] * mat_B[207][1] +
                mat_A[102][2] * mat_B[215][1] +
                mat_A[102][3] * mat_B[223][1] +
                mat_A[103][0] * mat_B[231][1] +
                mat_A[103][1] * mat_B[239][1] +
                mat_A[103][2] * mat_B[247][1] +
                mat_A[103][3] * mat_B[255][1];
    mat_C[103][2] <=
                mat_A[96][0] * mat_B[7][2] +
                mat_A[96][1] * mat_B[15][2] +
                mat_A[96][2] * mat_B[23][2] +
                mat_A[96][3] * mat_B[31][2] +
                mat_A[97][0] * mat_B[39][2] +
                mat_A[97][1] * mat_B[47][2] +
                mat_A[97][2] * mat_B[55][2] +
                mat_A[97][3] * mat_B[63][2] +
                mat_A[98][0] * mat_B[71][2] +
                mat_A[98][1] * mat_B[79][2] +
                mat_A[98][2] * mat_B[87][2] +
                mat_A[98][3] * mat_B[95][2] +
                mat_A[99][0] * mat_B[103][2] +
                mat_A[99][1] * mat_B[111][2] +
                mat_A[99][2] * mat_B[119][2] +
                mat_A[99][3] * mat_B[127][2] +
                mat_A[100][0] * mat_B[135][2] +
                mat_A[100][1] * mat_B[143][2] +
                mat_A[100][2] * mat_B[151][2] +
                mat_A[100][3] * mat_B[159][2] +
                mat_A[101][0] * mat_B[167][2] +
                mat_A[101][1] * mat_B[175][2] +
                mat_A[101][2] * mat_B[183][2] +
                mat_A[101][3] * mat_B[191][2] +
                mat_A[102][0] * mat_B[199][2] +
                mat_A[102][1] * mat_B[207][2] +
                mat_A[102][2] * mat_B[215][2] +
                mat_A[102][3] * mat_B[223][2] +
                mat_A[103][0] * mat_B[231][2] +
                mat_A[103][1] * mat_B[239][2] +
                mat_A[103][2] * mat_B[247][2] +
                mat_A[103][3] * mat_B[255][2];
    mat_C[103][3] <=
                mat_A[96][0] * mat_B[7][3] +
                mat_A[96][1] * mat_B[15][3] +
                mat_A[96][2] * mat_B[23][3] +
                mat_A[96][3] * mat_B[31][3] +
                mat_A[97][0] * mat_B[39][3] +
                mat_A[97][1] * mat_B[47][3] +
                mat_A[97][2] * mat_B[55][3] +
                mat_A[97][3] * mat_B[63][3] +
                mat_A[98][0] * mat_B[71][3] +
                mat_A[98][1] * mat_B[79][3] +
                mat_A[98][2] * mat_B[87][3] +
                mat_A[98][3] * mat_B[95][3] +
                mat_A[99][0] * mat_B[103][3] +
                mat_A[99][1] * mat_B[111][3] +
                mat_A[99][2] * mat_B[119][3] +
                mat_A[99][3] * mat_B[127][3] +
                mat_A[100][0] * mat_B[135][3] +
                mat_A[100][1] * mat_B[143][3] +
                mat_A[100][2] * mat_B[151][3] +
                mat_A[100][3] * mat_B[159][3] +
                mat_A[101][0] * mat_B[167][3] +
                mat_A[101][1] * mat_B[175][3] +
                mat_A[101][2] * mat_B[183][3] +
                mat_A[101][3] * mat_B[191][3] +
                mat_A[102][0] * mat_B[199][3] +
                mat_A[102][1] * mat_B[207][3] +
                mat_A[102][2] * mat_B[215][3] +
                mat_A[102][3] * mat_B[223][3] +
                mat_A[103][0] * mat_B[231][3] +
                mat_A[103][1] * mat_B[239][3] +
                mat_A[103][2] * mat_B[247][3] +
                mat_A[103][3] * mat_B[255][3];
    mat_C[104][0] <=
                mat_A[104][0] * mat_B[0][0] +
                mat_A[104][1] * mat_B[8][0] +
                mat_A[104][2] * mat_B[16][0] +
                mat_A[104][3] * mat_B[24][0] +
                mat_A[105][0] * mat_B[32][0] +
                mat_A[105][1] * mat_B[40][0] +
                mat_A[105][2] * mat_B[48][0] +
                mat_A[105][3] * mat_B[56][0] +
                mat_A[106][0] * mat_B[64][0] +
                mat_A[106][1] * mat_B[72][0] +
                mat_A[106][2] * mat_B[80][0] +
                mat_A[106][3] * mat_B[88][0] +
                mat_A[107][0] * mat_B[96][0] +
                mat_A[107][1] * mat_B[104][0] +
                mat_A[107][2] * mat_B[112][0] +
                mat_A[107][3] * mat_B[120][0] +
                mat_A[108][0] * mat_B[128][0] +
                mat_A[108][1] * mat_B[136][0] +
                mat_A[108][2] * mat_B[144][0] +
                mat_A[108][3] * mat_B[152][0] +
                mat_A[109][0] * mat_B[160][0] +
                mat_A[109][1] * mat_B[168][0] +
                mat_A[109][2] * mat_B[176][0] +
                mat_A[109][3] * mat_B[184][0] +
                mat_A[110][0] * mat_B[192][0] +
                mat_A[110][1] * mat_B[200][0] +
                mat_A[110][2] * mat_B[208][0] +
                mat_A[110][3] * mat_B[216][0] +
                mat_A[111][0] * mat_B[224][0] +
                mat_A[111][1] * mat_B[232][0] +
                mat_A[111][2] * mat_B[240][0] +
                mat_A[111][3] * mat_B[248][0];
    mat_C[104][1] <=
                mat_A[104][0] * mat_B[0][1] +
                mat_A[104][1] * mat_B[8][1] +
                mat_A[104][2] * mat_B[16][1] +
                mat_A[104][3] * mat_B[24][1] +
                mat_A[105][0] * mat_B[32][1] +
                mat_A[105][1] * mat_B[40][1] +
                mat_A[105][2] * mat_B[48][1] +
                mat_A[105][3] * mat_B[56][1] +
                mat_A[106][0] * mat_B[64][1] +
                mat_A[106][1] * mat_B[72][1] +
                mat_A[106][2] * mat_B[80][1] +
                mat_A[106][3] * mat_B[88][1] +
                mat_A[107][0] * mat_B[96][1] +
                mat_A[107][1] * mat_B[104][1] +
                mat_A[107][2] * mat_B[112][1] +
                mat_A[107][3] * mat_B[120][1] +
                mat_A[108][0] * mat_B[128][1] +
                mat_A[108][1] * mat_B[136][1] +
                mat_A[108][2] * mat_B[144][1] +
                mat_A[108][3] * mat_B[152][1] +
                mat_A[109][0] * mat_B[160][1] +
                mat_A[109][1] * mat_B[168][1] +
                mat_A[109][2] * mat_B[176][1] +
                mat_A[109][3] * mat_B[184][1] +
                mat_A[110][0] * mat_B[192][1] +
                mat_A[110][1] * mat_B[200][1] +
                mat_A[110][2] * mat_B[208][1] +
                mat_A[110][3] * mat_B[216][1] +
                mat_A[111][0] * mat_B[224][1] +
                mat_A[111][1] * mat_B[232][1] +
                mat_A[111][2] * mat_B[240][1] +
                mat_A[111][3] * mat_B[248][1];
    mat_C[104][2] <=
                mat_A[104][0] * mat_B[0][2] +
                mat_A[104][1] * mat_B[8][2] +
                mat_A[104][2] * mat_B[16][2] +
                mat_A[104][3] * mat_B[24][2] +
                mat_A[105][0] * mat_B[32][2] +
                mat_A[105][1] * mat_B[40][2] +
                mat_A[105][2] * mat_B[48][2] +
                mat_A[105][3] * mat_B[56][2] +
                mat_A[106][0] * mat_B[64][2] +
                mat_A[106][1] * mat_B[72][2] +
                mat_A[106][2] * mat_B[80][2] +
                mat_A[106][3] * mat_B[88][2] +
                mat_A[107][0] * mat_B[96][2] +
                mat_A[107][1] * mat_B[104][2] +
                mat_A[107][2] * mat_B[112][2] +
                mat_A[107][3] * mat_B[120][2] +
                mat_A[108][0] * mat_B[128][2] +
                mat_A[108][1] * mat_B[136][2] +
                mat_A[108][2] * mat_B[144][2] +
                mat_A[108][3] * mat_B[152][2] +
                mat_A[109][0] * mat_B[160][2] +
                mat_A[109][1] * mat_B[168][2] +
                mat_A[109][2] * mat_B[176][2] +
                mat_A[109][3] * mat_B[184][2] +
                mat_A[110][0] * mat_B[192][2] +
                mat_A[110][1] * mat_B[200][2] +
                mat_A[110][2] * mat_B[208][2] +
                mat_A[110][3] * mat_B[216][2] +
                mat_A[111][0] * mat_B[224][2] +
                mat_A[111][1] * mat_B[232][2] +
                mat_A[111][2] * mat_B[240][2] +
                mat_A[111][3] * mat_B[248][2];
    mat_C[104][3] <=
                mat_A[104][0] * mat_B[0][3] +
                mat_A[104][1] * mat_B[8][3] +
                mat_A[104][2] * mat_B[16][3] +
                mat_A[104][3] * mat_B[24][3] +
                mat_A[105][0] * mat_B[32][3] +
                mat_A[105][1] * mat_B[40][3] +
                mat_A[105][2] * mat_B[48][3] +
                mat_A[105][3] * mat_B[56][3] +
                mat_A[106][0] * mat_B[64][3] +
                mat_A[106][1] * mat_B[72][3] +
                mat_A[106][2] * mat_B[80][3] +
                mat_A[106][3] * mat_B[88][3] +
                mat_A[107][0] * mat_B[96][3] +
                mat_A[107][1] * mat_B[104][3] +
                mat_A[107][2] * mat_B[112][3] +
                mat_A[107][3] * mat_B[120][3] +
                mat_A[108][0] * mat_B[128][3] +
                mat_A[108][1] * mat_B[136][3] +
                mat_A[108][2] * mat_B[144][3] +
                mat_A[108][3] * mat_B[152][3] +
                mat_A[109][0] * mat_B[160][3] +
                mat_A[109][1] * mat_B[168][3] +
                mat_A[109][2] * mat_B[176][3] +
                mat_A[109][3] * mat_B[184][3] +
                mat_A[110][0] * mat_B[192][3] +
                mat_A[110][1] * mat_B[200][3] +
                mat_A[110][2] * mat_B[208][3] +
                mat_A[110][3] * mat_B[216][3] +
                mat_A[111][0] * mat_B[224][3] +
                mat_A[111][1] * mat_B[232][3] +
                mat_A[111][2] * mat_B[240][3] +
                mat_A[111][3] * mat_B[248][3];
    mat_C[105][0] <=
                mat_A[104][0] * mat_B[1][0] +
                mat_A[104][1] * mat_B[9][0] +
                mat_A[104][2] * mat_B[17][0] +
                mat_A[104][3] * mat_B[25][0] +
                mat_A[105][0] * mat_B[33][0] +
                mat_A[105][1] * mat_B[41][0] +
                mat_A[105][2] * mat_B[49][0] +
                mat_A[105][3] * mat_B[57][0] +
                mat_A[106][0] * mat_B[65][0] +
                mat_A[106][1] * mat_B[73][0] +
                mat_A[106][2] * mat_B[81][0] +
                mat_A[106][3] * mat_B[89][0] +
                mat_A[107][0] * mat_B[97][0] +
                mat_A[107][1] * mat_B[105][0] +
                mat_A[107][2] * mat_B[113][0] +
                mat_A[107][3] * mat_B[121][0] +
                mat_A[108][0] * mat_B[129][0] +
                mat_A[108][1] * mat_B[137][0] +
                mat_A[108][2] * mat_B[145][0] +
                mat_A[108][3] * mat_B[153][0] +
                mat_A[109][0] * mat_B[161][0] +
                mat_A[109][1] * mat_B[169][0] +
                mat_A[109][2] * mat_B[177][0] +
                mat_A[109][3] * mat_B[185][0] +
                mat_A[110][0] * mat_B[193][0] +
                mat_A[110][1] * mat_B[201][0] +
                mat_A[110][2] * mat_B[209][0] +
                mat_A[110][3] * mat_B[217][0] +
                mat_A[111][0] * mat_B[225][0] +
                mat_A[111][1] * mat_B[233][0] +
                mat_A[111][2] * mat_B[241][0] +
                mat_A[111][3] * mat_B[249][0];
    mat_C[105][1] <=
                mat_A[104][0] * mat_B[1][1] +
                mat_A[104][1] * mat_B[9][1] +
                mat_A[104][2] * mat_B[17][1] +
                mat_A[104][3] * mat_B[25][1] +
                mat_A[105][0] * mat_B[33][1] +
                mat_A[105][1] * mat_B[41][1] +
                mat_A[105][2] * mat_B[49][1] +
                mat_A[105][3] * mat_B[57][1] +
                mat_A[106][0] * mat_B[65][1] +
                mat_A[106][1] * mat_B[73][1] +
                mat_A[106][2] * mat_B[81][1] +
                mat_A[106][3] * mat_B[89][1] +
                mat_A[107][0] * mat_B[97][1] +
                mat_A[107][1] * mat_B[105][1] +
                mat_A[107][2] * mat_B[113][1] +
                mat_A[107][3] * mat_B[121][1] +
                mat_A[108][0] * mat_B[129][1] +
                mat_A[108][1] * mat_B[137][1] +
                mat_A[108][2] * mat_B[145][1] +
                mat_A[108][3] * mat_B[153][1] +
                mat_A[109][0] * mat_B[161][1] +
                mat_A[109][1] * mat_B[169][1] +
                mat_A[109][2] * mat_B[177][1] +
                mat_A[109][3] * mat_B[185][1] +
                mat_A[110][0] * mat_B[193][1] +
                mat_A[110][1] * mat_B[201][1] +
                mat_A[110][2] * mat_B[209][1] +
                mat_A[110][3] * mat_B[217][1] +
                mat_A[111][0] * mat_B[225][1] +
                mat_A[111][1] * mat_B[233][1] +
                mat_A[111][2] * mat_B[241][1] +
                mat_A[111][3] * mat_B[249][1];
    mat_C[105][2] <=
                mat_A[104][0] * mat_B[1][2] +
                mat_A[104][1] * mat_B[9][2] +
                mat_A[104][2] * mat_B[17][2] +
                mat_A[104][3] * mat_B[25][2] +
                mat_A[105][0] * mat_B[33][2] +
                mat_A[105][1] * mat_B[41][2] +
                mat_A[105][2] * mat_B[49][2] +
                mat_A[105][3] * mat_B[57][2] +
                mat_A[106][0] * mat_B[65][2] +
                mat_A[106][1] * mat_B[73][2] +
                mat_A[106][2] * mat_B[81][2] +
                mat_A[106][3] * mat_B[89][2] +
                mat_A[107][0] * mat_B[97][2] +
                mat_A[107][1] * mat_B[105][2] +
                mat_A[107][2] * mat_B[113][2] +
                mat_A[107][3] * mat_B[121][2] +
                mat_A[108][0] * mat_B[129][2] +
                mat_A[108][1] * mat_B[137][2] +
                mat_A[108][2] * mat_B[145][2] +
                mat_A[108][3] * mat_B[153][2] +
                mat_A[109][0] * mat_B[161][2] +
                mat_A[109][1] * mat_B[169][2] +
                mat_A[109][2] * mat_B[177][2] +
                mat_A[109][3] * mat_B[185][2] +
                mat_A[110][0] * mat_B[193][2] +
                mat_A[110][1] * mat_B[201][2] +
                mat_A[110][2] * mat_B[209][2] +
                mat_A[110][3] * mat_B[217][2] +
                mat_A[111][0] * mat_B[225][2] +
                mat_A[111][1] * mat_B[233][2] +
                mat_A[111][2] * mat_B[241][2] +
                mat_A[111][3] * mat_B[249][2];
    mat_C[105][3] <=
                mat_A[104][0] * mat_B[1][3] +
                mat_A[104][1] * mat_B[9][3] +
                mat_A[104][2] * mat_B[17][3] +
                mat_A[104][3] * mat_B[25][3] +
                mat_A[105][0] * mat_B[33][3] +
                mat_A[105][1] * mat_B[41][3] +
                mat_A[105][2] * mat_B[49][3] +
                mat_A[105][3] * mat_B[57][3] +
                mat_A[106][0] * mat_B[65][3] +
                mat_A[106][1] * mat_B[73][3] +
                mat_A[106][2] * mat_B[81][3] +
                mat_A[106][3] * mat_B[89][3] +
                mat_A[107][0] * mat_B[97][3] +
                mat_A[107][1] * mat_B[105][3] +
                mat_A[107][2] * mat_B[113][3] +
                mat_A[107][3] * mat_B[121][3] +
                mat_A[108][0] * mat_B[129][3] +
                mat_A[108][1] * mat_B[137][3] +
                mat_A[108][2] * mat_B[145][3] +
                mat_A[108][3] * mat_B[153][3] +
                mat_A[109][0] * mat_B[161][3] +
                mat_A[109][1] * mat_B[169][3] +
                mat_A[109][2] * mat_B[177][3] +
                mat_A[109][3] * mat_B[185][3] +
                mat_A[110][0] * mat_B[193][3] +
                mat_A[110][1] * mat_B[201][3] +
                mat_A[110][2] * mat_B[209][3] +
                mat_A[110][3] * mat_B[217][3] +
                mat_A[111][0] * mat_B[225][3] +
                mat_A[111][1] * mat_B[233][3] +
                mat_A[111][2] * mat_B[241][3] +
                mat_A[111][3] * mat_B[249][3];
    mat_C[106][0] <=
                mat_A[104][0] * mat_B[2][0] +
                mat_A[104][1] * mat_B[10][0] +
                mat_A[104][2] * mat_B[18][0] +
                mat_A[104][3] * mat_B[26][0] +
                mat_A[105][0] * mat_B[34][0] +
                mat_A[105][1] * mat_B[42][0] +
                mat_A[105][2] * mat_B[50][0] +
                mat_A[105][3] * mat_B[58][0] +
                mat_A[106][0] * mat_B[66][0] +
                mat_A[106][1] * mat_B[74][0] +
                mat_A[106][2] * mat_B[82][0] +
                mat_A[106][3] * mat_B[90][0] +
                mat_A[107][0] * mat_B[98][0] +
                mat_A[107][1] * mat_B[106][0] +
                mat_A[107][2] * mat_B[114][0] +
                mat_A[107][3] * mat_B[122][0] +
                mat_A[108][0] * mat_B[130][0] +
                mat_A[108][1] * mat_B[138][0] +
                mat_A[108][2] * mat_B[146][0] +
                mat_A[108][3] * mat_B[154][0] +
                mat_A[109][0] * mat_B[162][0] +
                mat_A[109][1] * mat_B[170][0] +
                mat_A[109][2] * mat_B[178][0] +
                mat_A[109][3] * mat_B[186][0] +
                mat_A[110][0] * mat_B[194][0] +
                mat_A[110][1] * mat_B[202][0] +
                mat_A[110][2] * mat_B[210][0] +
                mat_A[110][3] * mat_B[218][0] +
                mat_A[111][0] * mat_B[226][0] +
                mat_A[111][1] * mat_B[234][0] +
                mat_A[111][2] * mat_B[242][0] +
                mat_A[111][3] * mat_B[250][0];
    mat_C[106][1] <=
                mat_A[104][0] * mat_B[2][1] +
                mat_A[104][1] * mat_B[10][1] +
                mat_A[104][2] * mat_B[18][1] +
                mat_A[104][3] * mat_B[26][1] +
                mat_A[105][0] * mat_B[34][1] +
                mat_A[105][1] * mat_B[42][1] +
                mat_A[105][2] * mat_B[50][1] +
                mat_A[105][3] * mat_B[58][1] +
                mat_A[106][0] * mat_B[66][1] +
                mat_A[106][1] * mat_B[74][1] +
                mat_A[106][2] * mat_B[82][1] +
                mat_A[106][3] * mat_B[90][1] +
                mat_A[107][0] * mat_B[98][1] +
                mat_A[107][1] * mat_B[106][1] +
                mat_A[107][2] * mat_B[114][1] +
                mat_A[107][3] * mat_B[122][1] +
                mat_A[108][0] * mat_B[130][1] +
                mat_A[108][1] * mat_B[138][1] +
                mat_A[108][2] * mat_B[146][1] +
                mat_A[108][3] * mat_B[154][1] +
                mat_A[109][0] * mat_B[162][1] +
                mat_A[109][1] * mat_B[170][1] +
                mat_A[109][2] * mat_B[178][1] +
                mat_A[109][3] * mat_B[186][1] +
                mat_A[110][0] * mat_B[194][1] +
                mat_A[110][1] * mat_B[202][1] +
                mat_A[110][2] * mat_B[210][1] +
                mat_A[110][3] * mat_B[218][1] +
                mat_A[111][0] * mat_B[226][1] +
                mat_A[111][1] * mat_B[234][1] +
                mat_A[111][2] * mat_B[242][1] +
                mat_A[111][3] * mat_B[250][1];
    mat_C[106][2] <=
                mat_A[104][0] * mat_B[2][2] +
                mat_A[104][1] * mat_B[10][2] +
                mat_A[104][2] * mat_B[18][2] +
                mat_A[104][3] * mat_B[26][2] +
                mat_A[105][0] * mat_B[34][2] +
                mat_A[105][1] * mat_B[42][2] +
                mat_A[105][2] * mat_B[50][2] +
                mat_A[105][3] * mat_B[58][2] +
                mat_A[106][0] * mat_B[66][2] +
                mat_A[106][1] * mat_B[74][2] +
                mat_A[106][2] * mat_B[82][2] +
                mat_A[106][3] * mat_B[90][2] +
                mat_A[107][0] * mat_B[98][2] +
                mat_A[107][1] * mat_B[106][2] +
                mat_A[107][2] * mat_B[114][2] +
                mat_A[107][3] * mat_B[122][2] +
                mat_A[108][0] * mat_B[130][2] +
                mat_A[108][1] * mat_B[138][2] +
                mat_A[108][2] * mat_B[146][2] +
                mat_A[108][3] * mat_B[154][2] +
                mat_A[109][0] * mat_B[162][2] +
                mat_A[109][1] * mat_B[170][2] +
                mat_A[109][2] * mat_B[178][2] +
                mat_A[109][3] * mat_B[186][2] +
                mat_A[110][0] * mat_B[194][2] +
                mat_A[110][1] * mat_B[202][2] +
                mat_A[110][2] * mat_B[210][2] +
                mat_A[110][3] * mat_B[218][2] +
                mat_A[111][0] * mat_B[226][2] +
                mat_A[111][1] * mat_B[234][2] +
                mat_A[111][2] * mat_B[242][2] +
                mat_A[111][3] * mat_B[250][2];
    mat_C[106][3] <=
                mat_A[104][0] * mat_B[2][3] +
                mat_A[104][1] * mat_B[10][3] +
                mat_A[104][2] * mat_B[18][3] +
                mat_A[104][3] * mat_B[26][3] +
                mat_A[105][0] * mat_B[34][3] +
                mat_A[105][1] * mat_B[42][3] +
                mat_A[105][2] * mat_B[50][3] +
                mat_A[105][3] * mat_B[58][3] +
                mat_A[106][0] * mat_B[66][3] +
                mat_A[106][1] * mat_B[74][3] +
                mat_A[106][2] * mat_B[82][3] +
                mat_A[106][3] * mat_B[90][3] +
                mat_A[107][0] * mat_B[98][3] +
                mat_A[107][1] * mat_B[106][3] +
                mat_A[107][2] * mat_B[114][3] +
                mat_A[107][3] * mat_B[122][3] +
                mat_A[108][0] * mat_B[130][3] +
                mat_A[108][1] * mat_B[138][3] +
                mat_A[108][2] * mat_B[146][3] +
                mat_A[108][3] * mat_B[154][3] +
                mat_A[109][0] * mat_B[162][3] +
                mat_A[109][1] * mat_B[170][3] +
                mat_A[109][2] * mat_B[178][3] +
                mat_A[109][3] * mat_B[186][3] +
                mat_A[110][0] * mat_B[194][3] +
                mat_A[110][1] * mat_B[202][3] +
                mat_A[110][2] * mat_B[210][3] +
                mat_A[110][3] * mat_B[218][3] +
                mat_A[111][0] * mat_B[226][3] +
                mat_A[111][1] * mat_B[234][3] +
                mat_A[111][2] * mat_B[242][3] +
                mat_A[111][3] * mat_B[250][3];
    mat_C[107][0] <=
                mat_A[104][0] * mat_B[3][0] +
                mat_A[104][1] * mat_B[11][0] +
                mat_A[104][2] * mat_B[19][0] +
                mat_A[104][3] * mat_B[27][0] +
                mat_A[105][0] * mat_B[35][0] +
                mat_A[105][1] * mat_B[43][0] +
                mat_A[105][2] * mat_B[51][0] +
                mat_A[105][3] * mat_B[59][0] +
                mat_A[106][0] * mat_B[67][0] +
                mat_A[106][1] * mat_B[75][0] +
                mat_A[106][2] * mat_B[83][0] +
                mat_A[106][3] * mat_B[91][0] +
                mat_A[107][0] * mat_B[99][0] +
                mat_A[107][1] * mat_B[107][0] +
                mat_A[107][2] * mat_B[115][0] +
                mat_A[107][3] * mat_B[123][0] +
                mat_A[108][0] * mat_B[131][0] +
                mat_A[108][1] * mat_B[139][0] +
                mat_A[108][2] * mat_B[147][0] +
                mat_A[108][3] * mat_B[155][0] +
                mat_A[109][0] * mat_B[163][0] +
                mat_A[109][1] * mat_B[171][0] +
                mat_A[109][2] * mat_B[179][0] +
                mat_A[109][3] * mat_B[187][0] +
                mat_A[110][0] * mat_B[195][0] +
                mat_A[110][1] * mat_B[203][0] +
                mat_A[110][2] * mat_B[211][0] +
                mat_A[110][3] * mat_B[219][0] +
                mat_A[111][0] * mat_B[227][0] +
                mat_A[111][1] * mat_B[235][0] +
                mat_A[111][2] * mat_B[243][0] +
                mat_A[111][3] * mat_B[251][0];
    mat_C[107][1] <=
                mat_A[104][0] * mat_B[3][1] +
                mat_A[104][1] * mat_B[11][1] +
                mat_A[104][2] * mat_B[19][1] +
                mat_A[104][3] * mat_B[27][1] +
                mat_A[105][0] * mat_B[35][1] +
                mat_A[105][1] * mat_B[43][1] +
                mat_A[105][2] * mat_B[51][1] +
                mat_A[105][3] * mat_B[59][1] +
                mat_A[106][0] * mat_B[67][1] +
                mat_A[106][1] * mat_B[75][1] +
                mat_A[106][2] * mat_B[83][1] +
                mat_A[106][3] * mat_B[91][1] +
                mat_A[107][0] * mat_B[99][1] +
                mat_A[107][1] * mat_B[107][1] +
                mat_A[107][2] * mat_B[115][1] +
                mat_A[107][3] * mat_B[123][1] +
                mat_A[108][0] * mat_B[131][1] +
                mat_A[108][1] * mat_B[139][1] +
                mat_A[108][2] * mat_B[147][1] +
                mat_A[108][3] * mat_B[155][1] +
                mat_A[109][0] * mat_B[163][1] +
                mat_A[109][1] * mat_B[171][1] +
                mat_A[109][2] * mat_B[179][1] +
                mat_A[109][3] * mat_B[187][1] +
                mat_A[110][0] * mat_B[195][1] +
                mat_A[110][1] * mat_B[203][1] +
                mat_A[110][2] * mat_B[211][1] +
                mat_A[110][3] * mat_B[219][1] +
                mat_A[111][0] * mat_B[227][1] +
                mat_A[111][1] * mat_B[235][1] +
                mat_A[111][2] * mat_B[243][1] +
                mat_A[111][3] * mat_B[251][1];
    mat_C[107][2] <=
                mat_A[104][0] * mat_B[3][2] +
                mat_A[104][1] * mat_B[11][2] +
                mat_A[104][2] * mat_B[19][2] +
                mat_A[104][3] * mat_B[27][2] +
                mat_A[105][0] * mat_B[35][2] +
                mat_A[105][1] * mat_B[43][2] +
                mat_A[105][2] * mat_B[51][2] +
                mat_A[105][3] * mat_B[59][2] +
                mat_A[106][0] * mat_B[67][2] +
                mat_A[106][1] * mat_B[75][2] +
                mat_A[106][2] * mat_B[83][2] +
                mat_A[106][3] * mat_B[91][2] +
                mat_A[107][0] * mat_B[99][2] +
                mat_A[107][1] * mat_B[107][2] +
                mat_A[107][2] * mat_B[115][2] +
                mat_A[107][3] * mat_B[123][2] +
                mat_A[108][0] * mat_B[131][2] +
                mat_A[108][1] * mat_B[139][2] +
                mat_A[108][2] * mat_B[147][2] +
                mat_A[108][3] * mat_B[155][2] +
                mat_A[109][0] * mat_B[163][2] +
                mat_A[109][1] * mat_B[171][2] +
                mat_A[109][2] * mat_B[179][2] +
                mat_A[109][3] * mat_B[187][2] +
                mat_A[110][0] * mat_B[195][2] +
                mat_A[110][1] * mat_B[203][2] +
                mat_A[110][2] * mat_B[211][2] +
                mat_A[110][3] * mat_B[219][2] +
                mat_A[111][0] * mat_B[227][2] +
                mat_A[111][1] * mat_B[235][2] +
                mat_A[111][2] * mat_B[243][2] +
                mat_A[111][3] * mat_B[251][2];
    mat_C[107][3] <=
                mat_A[104][0] * mat_B[3][3] +
                mat_A[104][1] * mat_B[11][3] +
                mat_A[104][2] * mat_B[19][3] +
                mat_A[104][3] * mat_B[27][3] +
                mat_A[105][0] * mat_B[35][3] +
                mat_A[105][1] * mat_B[43][3] +
                mat_A[105][2] * mat_B[51][3] +
                mat_A[105][3] * mat_B[59][3] +
                mat_A[106][0] * mat_B[67][3] +
                mat_A[106][1] * mat_B[75][3] +
                mat_A[106][2] * mat_B[83][3] +
                mat_A[106][3] * mat_B[91][3] +
                mat_A[107][0] * mat_B[99][3] +
                mat_A[107][1] * mat_B[107][3] +
                mat_A[107][2] * mat_B[115][3] +
                mat_A[107][3] * mat_B[123][3] +
                mat_A[108][0] * mat_B[131][3] +
                mat_A[108][1] * mat_B[139][3] +
                mat_A[108][2] * mat_B[147][3] +
                mat_A[108][3] * mat_B[155][3] +
                mat_A[109][0] * mat_B[163][3] +
                mat_A[109][1] * mat_B[171][3] +
                mat_A[109][2] * mat_B[179][3] +
                mat_A[109][3] * mat_B[187][3] +
                mat_A[110][0] * mat_B[195][3] +
                mat_A[110][1] * mat_B[203][3] +
                mat_A[110][2] * mat_B[211][3] +
                mat_A[110][3] * mat_B[219][3] +
                mat_A[111][0] * mat_B[227][3] +
                mat_A[111][1] * mat_B[235][3] +
                mat_A[111][2] * mat_B[243][3] +
                mat_A[111][3] * mat_B[251][3];
    mat_C[108][0] <=
                mat_A[104][0] * mat_B[4][0] +
                mat_A[104][1] * mat_B[12][0] +
                mat_A[104][2] * mat_B[20][0] +
                mat_A[104][3] * mat_B[28][0] +
                mat_A[105][0] * mat_B[36][0] +
                mat_A[105][1] * mat_B[44][0] +
                mat_A[105][2] * mat_B[52][0] +
                mat_A[105][3] * mat_B[60][0] +
                mat_A[106][0] * mat_B[68][0] +
                mat_A[106][1] * mat_B[76][0] +
                mat_A[106][2] * mat_B[84][0] +
                mat_A[106][3] * mat_B[92][0] +
                mat_A[107][0] * mat_B[100][0] +
                mat_A[107][1] * mat_B[108][0] +
                mat_A[107][2] * mat_B[116][0] +
                mat_A[107][3] * mat_B[124][0] +
                mat_A[108][0] * mat_B[132][0] +
                mat_A[108][1] * mat_B[140][0] +
                mat_A[108][2] * mat_B[148][0] +
                mat_A[108][3] * mat_B[156][0] +
                mat_A[109][0] * mat_B[164][0] +
                mat_A[109][1] * mat_B[172][0] +
                mat_A[109][2] * mat_B[180][0] +
                mat_A[109][3] * mat_B[188][0] +
                mat_A[110][0] * mat_B[196][0] +
                mat_A[110][1] * mat_B[204][0] +
                mat_A[110][2] * mat_B[212][0] +
                mat_A[110][3] * mat_B[220][0] +
                mat_A[111][0] * mat_B[228][0] +
                mat_A[111][1] * mat_B[236][0] +
                mat_A[111][2] * mat_B[244][0] +
                mat_A[111][3] * mat_B[252][0];
    mat_C[108][1] <=
                mat_A[104][0] * mat_B[4][1] +
                mat_A[104][1] * mat_B[12][1] +
                mat_A[104][2] * mat_B[20][1] +
                mat_A[104][3] * mat_B[28][1] +
                mat_A[105][0] * mat_B[36][1] +
                mat_A[105][1] * mat_B[44][1] +
                mat_A[105][2] * mat_B[52][1] +
                mat_A[105][3] * mat_B[60][1] +
                mat_A[106][0] * mat_B[68][1] +
                mat_A[106][1] * mat_B[76][1] +
                mat_A[106][2] * mat_B[84][1] +
                mat_A[106][3] * mat_B[92][1] +
                mat_A[107][0] * mat_B[100][1] +
                mat_A[107][1] * mat_B[108][1] +
                mat_A[107][2] * mat_B[116][1] +
                mat_A[107][3] * mat_B[124][1] +
                mat_A[108][0] * mat_B[132][1] +
                mat_A[108][1] * mat_B[140][1] +
                mat_A[108][2] * mat_B[148][1] +
                mat_A[108][3] * mat_B[156][1] +
                mat_A[109][0] * mat_B[164][1] +
                mat_A[109][1] * mat_B[172][1] +
                mat_A[109][2] * mat_B[180][1] +
                mat_A[109][3] * mat_B[188][1] +
                mat_A[110][0] * mat_B[196][1] +
                mat_A[110][1] * mat_B[204][1] +
                mat_A[110][2] * mat_B[212][1] +
                mat_A[110][3] * mat_B[220][1] +
                mat_A[111][0] * mat_B[228][1] +
                mat_A[111][1] * mat_B[236][1] +
                mat_A[111][2] * mat_B[244][1] +
                mat_A[111][3] * mat_B[252][1];
    mat_C[108][2] <=
                mat_A[104][0] * mat_B[4][2] +
                mat_A[104][1] * mat_B[12][2] +
                mat_A[104][2] * mat_B[20][2] +
                mat_A[104][3] * mat_B[28][2] +
                mat_A[105][0] * mat_B[36][2] +
                mat_A[105][1] * mat_B[44][2] +
                mat_A[105][2] * mat_B[52][2] +
                mat_A[105][3] * mat_B[60][2] +
                mat_A[106][0] * mat_B[68][2] +
                mat_A[106][1] * mat_B[76][2] +
                mat_A[106][2] * mat_B[84][2] +
                mat_A[106][3] * mat_B[92][2] +
                mat_A[107][0] * mat_B[100][2] +
                mat_A[107][1] * mat_B[108][2] +
                mat_A[107][2] * mat_B[116][2] +
                mat_A[107][3] * mat_B[124][2] +
                mat_A[108][0] * mat_B[132][2] +
                mat_A[108][1] * mat_B[140][2] +
                mat_A[108][2] * mat_B[148][2] +
                mat_A[108][3] * mat_B[156][2] +
                mat_A[109][0] * mat_B[164][2] +
                mat_A[109][1] * mat_B[172][2] +
                mat_A[109][2] * mat_B[180][2] +
                mat_A[109][3] * mat_B[188][2] +
                mat_A[110][0] * mat_B[196][2] +
                mat_A[110][1] * mat_B[204][2] +
                mat_A[110][2] * mat_B[212][2] +
                mat_A[110][3] * mat_B[220][2] +
                mat_A[111][0] * mat_B[228][2] +
                mat_A[111][1] * mat_B[236][2] +
                mat_A[111][2] * mat_B[244][2] +
                mat_A[111][3] * mat_B[252][2];
    mat_C[108][3] <=
                mat_A[104][0] * mat_B[4][3] +
                mat_A[104][1] * mat_B[12][3] +
                mat_A[104][2] * mat_B[20][3] +
                mat_A[104][3] * mat_B[28][3] +
                mat_A[105][0] * mat_B[36][3] +
                mat_A[105][1] * mat_B[44][3] +
                mat_A[105][2] * mat_B[52][3] +
                mat_A[105][3] * mat_B[60][3] +
                mat_A[106][0] * mat_B[68][3] +
                mat_A[106][1] * mat_B[76][3] +
                mat_A[106][2] * mat_B[84][3] +
                mat_A[106][3] * mat_B[92][3] +
                mat_A[107][0] * mat_B[100][3] +
                mat_A[107][1] * mat_B[108][3] +
                mat_A[107][2] * mat_B[116][3] +
                mat_A[107][3] * mat_B[124][3] +
                mat_A[108][0] * mat_B[132][3] +
                mat_A[108][1] * mat_B[140][3] +
                mat_A[108][2] * mat_B[148][3] +
                mat_A[108][3] * mat_B[156][3] +
                mat_A[109][0] * mat_B[164][3] +
                mat_A[109][1] * mat_B[172][3] +
                mat_A[109][2] * mat_B[180][3] +
                mat_A[109][3] * mat_B[188][3] +
                mat_A[110][0] * mat_B[196][3] +
                mat_A[110][1] * mat_B[204][3] +
                mat_A[110][2] * mat_B[212][3] +
                mat_A[110][3] * mat_B[220][3] +
                mat_A[111][0] * mat_B[228][3] +
                mat_A[111][1] * mat_B[236][3] +
                mat_A[111][2] * mat_B[244][3] +
                mat_A[111][3] * mat_B[252][3];
    mat_C[109][0] <=
                mat_A[104][0] * mat_B[5][0] +
                mat_A[104][1] * mat_B[13][0] +
                mat_A[104][2] * mat_B[21][0] +
                mat_A[104][3] * mat_B[29][0] +
                mat_A[105][0] * mat_B[37][0] +
                mat_A[105][1] * mat_B[45][0] +
                mat_A[105][2] * mat_B[53][0] +
                mat_A[105][3] * mat_B[61][0] +
                mat_A[106][0] * mat_B[69][0] +
                mat_A[106][1] * mat_B[77][0] +
                mat_A[106][2] * mat_B[85][0] +
                mat_A[106][3] * mat_B[93][0] +
                mat_A[107][0] * mat_B[101][0] +
                mat_A[107][1] * mat_B[109][0] +
                mat_A[107][2] * mat_B[117][0] +
                mat_A[107][3] * mat_B[125][0] +
                mat_A[108][0] * mat_B[133][0] +
                mat_A[108][1] * mat_B[141][0] +
                mat_A[108][2] * mat_B[149][0] +
                mat_A[108][3] * mat_B[157][0] +
                mat_A[109][0] * mat_B[165][0] +
                mat_A[109][1] * mat_B[173][0] +
                mat_A[109][2] * mat_B[181][0] +
                mat_A[109][3] * mat_B[189][0] +
                mat_A[110][0] * mat_B[197][0] +
                mat_A[110][1] * mat_B[205][0] +
                mat_A[110][2] * mat_B[213][0] +
                mat_A[110][3] * mat_B[221][0] +
                mat_A[111][0] * mat_B[229][0] +
                mat_A[111][1] * mat_B[237][0] +
                mat_A[111][2] * mat_B[245][0] +
                mat_A[111][3] * mat_B[253][0];
    mat_C[109][1] <=
                mat_A[104][0] * mat_B[5][1] +
                mat_A[104][1] * mat_B[13][1] +
                mat_A[104][2] * mat_B[21][1] +
                mat_A[104][3] * mat_B[29][1] +
                mat_A[105][0] * mat_B[37][1] +
                mat_A[105][1] * mat_B[45][1] +
                mat_A[105][2] * mat_B[53][1] +
                mat_A[105][3] * mat_B[61][1] +
                mat_A[106][0] * mat_B[69][1] +
                mat_A[106][1] * mat_B[77][1] +
                mat_A[106][2] * mat_B[85][1] +
                mat_A[106][3] * mat_B[93][1] +
                mat_A[107][0] * mat_B[101][1] +
                mat_A[107][1] * mat_B[109][1] +
                mat_A[107][2] * mat_B[117][1] +
                mat_A[107][3] * mat_B[125][1] +
                mat_A[108][0] * mat_B[133][1] +
                mat_A[108][1] * mat_B[141][1] +
                mat_A[108][2] * mat_B[149][1] +
                mat_A[108][3] * mat_B[157][1] +
                mat_A[109][0] * mat_B[165][1] +
                mat_A[109][1] * mat_B[173][1] +
                mat_A[109][2] * mat_B[181][1] +
                mat_A[109][3] * mat_B[189][1] +
                mat_A[110][0] * mat_B[197][1] +
                mat_A[110][1] * mat_B[205][1] +
                mat_A[110][2] * mat_B[213][1] +
                mat_A[110][3] * mat_B[221][1] +
                mat_A[111][0] * mat_B[229][1] +
                mat_A[111][1] * mat_B[237][1] +
                mat_A[111][2] * mat_B[245][1] +
                mat_A[111][3] * mat_B[253][1];
    mat_C[109][2] <=
                mat_A[104][0] * mat_B[5][2] +
                mat_A[104][1] * mat_B[13][2] +
                mat_A[104][2] * mat_B[21][2] +
                mat_A[104][3] * mat_B[29][2] +
                mat_A[105][0] * mat_B[37][2] +
                mat_A[105][1] * mat_B[45][2] +
                mat_A[105][2] * mat_B[53][2] +
                mat_A[105][3] * mat_B[61][2] +
                mat_A[106][0] * mat_B[69][2] +
                mat_A[106][1] * mat_B[77][2] +
                mat_A[106][2] * mat_B[85][2] +
                mat_A[106][3] * mat_B[93][2] +
                mat_A[107][0] * mat_B[101][2] +
                mat_A[107][1] * mat_B[109][2] +
                mat_A[107][2] * mat_B[117][2] +
                mat_A[107][3] * mat_B[125][2] +
                mat_A[108][0] * mat_B[133][2] +
                mat_A[108][1] * mat_B[141][2] +
                mat_A[108][2] * mat_B[149][2] +
                mat_A[108][3] * mat_B[157][2] +
                mat_A[109][0] * mat_B[165][2] +
                mat_A[109][1] * mat_B[173][2] +
                mat_A[109][2] * mat_B[181][2] +
                mat_A[109][3] * mat_B[189][2] +
                mat_A[110][0] * mat_B[197][2] +
                mat_A[110][1] * mat_B[205][2] +
                mat_A[110][2] * mat_B[213][2] +
                mat_A[110][3] * mat_B[221][2] +
                mat_A[111][0] * mat_B[229][2] +
                mat_A[111][1] * mat_B[237][2] +
                mat_A[111][2] * mat_B[245][2] +
                mat_A[111][3] * mat_B[253][2];
    mat_C[109][3] <=
                mat_A[104][0] * mat_B[5][3] +
                mat_A[104][1] * mat_B[13][3] +
                mat_A[104][2] * mat_B[21][3] +
                mat_A[104][3] * mat_B[29][3] +
                mat_A[105][0] * mat_B[37][3] +
                mat_A[105][1] * mat_B[45][3] +
                mat_A[105][2] * mat_B[53][3] +
                mat_A[105][3] * mat_B[61][3] +
                mat_A[106][0] * mat_B[69][3] +
                mat_A[106][1] * mat_B[77][3] +
                mat_A[106][2] * mat_B[85][3] +
                mat_A[106][3] * mat_B[93][3] +
                mat_A[107][0] * mat_B[101][3] +
                mat_A[107][1] * mat_B[109][3] +
                mat_A[107][2] * mat_B[117][3] +
                mat_A[107][3] * mat_B[125][3] +
                mat_A[108][0] * mat_B[133][3] +
                mat_A[108][1] * mat_B[141][3] +
                mat_A[108][2] * mat_B[149][3] +
                mat_A[108][3] * mat_B[157][3] +
                mat_A[109][0] * mat_B[165][3] +
                mat_A[109][1] * mat_B[173][3] +
                mat_A[109][2] * mat_B[181][3] +
                mat_A[109][3] * mat_B[189][3] +
                mat_A[110][0] * mat_B[197][3] +
                mat_A[110][1] * mat_B[205][3] +
                mat_A[110][2] * mat_B[213][3] +
                mat_A[110][3] * mat_B[221][3] +
                mat_A[111][0] * mat_B[229][3] +
                mat_A[111][1] * mat_B[237][3] +
                mat_A[111][2] * mat_B[245][3] +
                mat_A[111][3] * mat_B[253][3];
    mat_C[110][0] <=
                mat_A[104][0] * mat_B[6][0] +
                mat_A[104][1] * mat_B[14][0] +
                mat_A[104][2] * mat_B[22][0] +
                mat_A[104][3] * mat_B[30][0] +
                mat_A[105][0] * mat_B[38][0] +
                mat_A[105][1] * mat_B[46][0] +
                mat_A[105][2] * mat_B[54][0] +
                mat_A[105][3] * mat_B[62][0] +
                mat_A[106][0] * mat_B[70][0] +
                mat_A[106][1] * mat_B[78][0] +
                mat_A[106][2] * mat_B[86][0] +
                mat_A[106][3] * mat_B[94][0] +
                mat_A[107][0] * mat_B[102][0] +
                mat_A[107][1] * mat_B[110][0] +
                mat_A[107][2] * mat_B[118][0] +
                mat_A[107][3] * mat_B[126][0] +
                mat_A[108][0] * mat_B[134][0] +
                mat_A[108][1] * mat_B[142][0] +
                mat_A[108][2] * mat_B[150][0] +
                mat_A[108][3] * mat_B[158][0] +
                mat_A[109][0] * mat_B[166][0] +
                mat_A[109][1] * mat_B[174][0] +
                mat_A[109][2] * mat_B[182][0] +
                mat_A[109][3] * mat_B[190][0] +
                mat_A[110][0] * mat_B[198][0] +
                mat_A[110][1] * mat_B[206][0] +
                mat_A[110][2] * mat_B[214][0] +
                mat_A[110][3] * mat_B[222][0] +
                mat_A[111][0] * mat_B[230][0] +
                mat_A[111][1] * mat_B[238][0] +
                mat_A[111][2] * mat_B[246][0] +
                mat_A[111][3] * mat_B[254][0];
    mat_C[110][1] <=
                mat_A[104][0] * mat_B[6][1] +
                mat_A[104][1] * mat_B[14][1] +
                mat_A[104][2] * mat_B[22][1] +
                mat_A[104][3] * mat_B[30][1] +
                mat_A[105][0] * mat_B[38][1] +
                mat_A[105][1] * mat_B[46][1] +
                mat_A[105][2] * mat_B[54][1] +
                mat_A[105][3] * mat_B[62][1] +
                mat_A[106][0] * mat_B[70][1] +
                mat_A[106][1] * mat_B[78][1] +
                mat_A[106][2] * mat_B[86][1] +
                mat_A[106][3] * mat_B[94][1] +
                mat_A[107][0] * mat_B[102][1] +
                mat_A[107][1] * mat_B[110][1] +
                mat_A[107][2] * mat_B[118][1] +
                mat_A[107][3] * mat_B[126][1] +
                mat_A[108][0] * mat_B[134][1] +
                mat_A[108][1] * mat_B[142][1] +
                mat_A[108][2] * mat_B[150][1] +
                mat_A[108][3] * mat_B[158][1] +
                mat_A[109][0] * mat_B[166][1] +
                mat_A[109][1] * mat_B[174][1] +
                mat_A[109][2] * mat_B[182][1] +
                mat_A[109][3] * mat_B[190][1] +
                mat_A[110][0] * mat_B[198][1] +
                mat_A[110][1] * mat_B[206][1] +
                mat_A[110][2] * mat_B[214][1] +
                mat_A[110][3] * mat_B[222][1] +
                mat_A[111][0] * mat_B[230][1] +
                mat_A[111][1] * mat_B[238][1] +
                mat_A[111][2] * mat_B[246][1] +
                mat_A[111][3] * mat_B[254][1];
    mat_C[110][2] <=
                mat_A[104][0] * mat_B[6][2] +
                mat_A[104][1] * mat_B[14][2] +
                mat_A[104][2] * mat_B[22][2] +
                mat_A[104][3] * mat_B[30][2] +
                mat_A[105][0] * mat_B[38][2] +
                mat_A[105][1] * mat_B[46][2] +
                mat_A[105][2] * mat_B[54][2] +
                mat_A[105][3] * mat_B[62][2] +
                mat_A[106][0] * mat_B[70][2] +
                mat_A[106][1] * mat_B[78][2] +
                mat_A[106][2] * mat_B[86][2] +
                mat_A[106][3] * mat_B[94][2] +
                mat_A[107][0] * mat_B[102][2] +
                mat_A[107][1] * mat_B[110][2] +
                mat_A[107][2] * mat_B[118][2] +
                mat_A[107][3] * mat_B[126][2] +
                mat_A[108][0] * mat_B[134][2] +
                mat_A[108][1] * mat_B[142][2] +
                mat_A[108][2] * mat_B[150][2] +
                mat_A[108][3] * mat_B[158][2] +
                mat_A[109][0] * mat_B[166][2] +
                mat_A[109][1] * mat_B[174][2] +
                mat_A[109][2] * mat_B[182][2] +
                mat_A[109][3] * mat_B[190][2] +
                mat_A[110][0] * mat_B[198][2] +
                mat_A[110][1] * mat_B[206][2] +
                mat_A[110][2] * mat_B[214][2] +
                mat_A[110][3] * mat_B[222][2] +
                mat_A[111][0] * mat_B[230][2] +
                mat_A[111][1] * mat_B[238][2] +
                mat_A[111][2] * mat_B[246][2] +
                mat_A[111][3] * mat_B[254][2];
    mat_C[110][3] <=
                mat_A[104][0] * mat_B[6][3] +
                mat_A[104][1] * mat_B[14][3] +
                mat_A[104][2] * mat_B[22][3] +
                mat_A[104][3] * mat_B[30][3] +
                mat_A[105][0] * mat_B[38][3] +
                mat_A[105][1] * mat_B[46][3] +
                mat_A[105][2] * mat_B[54][3] +
                mat_A[105][3] * mat_B[62][3] +
                mat_A[106][0] * mat_B[70][3] +
                mat_A[106][1] * mat_B[78][3] +
                mat_A[106][2] * mat_B[86][3] +
                mat_A[106][3] * mat_B[94][3] +
                mat_A[107][0] * mat_B[102][3] +
                mat_A[107][1] * mat_B[110][3] +
                mat_A[107][2] * mat_B[118][3] +
                mat_A[107][3] * mat_B[126][3] +
                mat_A[108][0] * mat_B[134][3] +
                mat_A[108][1] * mat_B[142][3] +
                mat_A[108][2] * mat_B[150][3] +
                mat_A[108][3] * mat_B[158][3] +
                mat_A[109][0] * mat_B[166][3] +
                mat_A[109][1] * mat_B[174][3] +
                mat_A[109][2] * mat_B[182][3] +
                mat_A[109][3] * mat_B[190][3] +
                mat_A[110][0] * mat_B[198][3] +
                mat_A[110][1] * mat_B[206][3] +
                mat_A[110][2] * mat_B[214][3] +
                mat_A[110][3] * mat_B[222][3] +
                mat_A[111][0] * mat_B[230][3] +
                mat_A[111][1] * mat_B[238][3] +
                mat_A[111][2] * mat_B[246][3] +
                mat_A[111][3] * mat_B[254][3];
    mat_C[111][0] <=
                mat_A[104][0] * mat_B[7][0] +
                mat_A[104][1] * mat_B[15][0] +
                mat_A[104][2] * mat_B[23][0] +
                mat_A[104][3] * mat_B[31][0] +
                mat_A[105][0] * mat_B[39][0] +
                mat_A[105][1] * mat_B[47][0] +
                mat_A[105][2] * mat_B[55][0] +
                mat_A[105][3] * mat_B[63][0] +
                mat_A[106][0] * mat_B[71][0] +
                mat_A[106][1] * mat_B[79][0] +
                mat_A[106][2] * mat_B[87][0] +
                mat_A[106][3] * mat_B[95][0] +
                mat_A[107][0] * mat_B[103][0] +
                mat_A[107][1] * mat_B[111][0] +
                mat_A[107][2] * mat_B[119][0] +
                mat_A[107][3] * mat_B[127][0] +
                mat_A[108][0] * mat_B[135][0] +
                mat_A[108][1] * mat_B[143][0] +
                mat_A[108][2] * mat_B[151][0] +
                mat_A[108][3] * mat_B[159][0] +
                mat_A[109][0] * mat_B[167][0] +
                mat_A[109][1] * mat_B[175][0] +
                mat_A[109][2] * mat_B[183][0] +
                mat_A[109][3] * mat_B[191][0] +
                mat_A[110][0] * mat_B[199][0] +
                mat_A[110][1] * mat_B[207][0] +
                mat_A[110][2] * mat_B[215][0] +
                mat_A[110][3] * mat_B[223][0] +
                mat_A[111][0] * mat_B[231][0] +
                mat_A[111][1] * mat_B[239][0] +
                mat_A[111][2] * mat_B[247][0] +
                mat_A[111][3] * mat_B[255][0];
    mat_C[111][1] <=
                mat_A[104][0] * mat_B[7][1] +
                mat_A[104][1] * mat_B[15][1] +
                mat_A[104][2] * mat_B[23][1] +
                mat_A[104][3] * mat_B[31][1] +
                mat_A[105][0] * mat_B[39][1] +
                mat_A[105][1] * mat_B[47][1] +
                mat_A[105][2] * mat_B[55][1] +
                mat_A[105][3] * mat_B[63][1] +
                mat_A[106][0] * mat_B[71][1] +
                mat_A[106][1] * mat_B[79][1] +
                mat_A[106][2] * mat_B[87][1] +
                mat_A[106][3] * mat_B[95][1] +
                mat_A[107][0] * mat_B[103][1] +
                mat_A[107][1] * mat_B[111][1] +
                mat_A[107][2] * mat_B[119][1] +
                mat_A[107][3] * mat_B[127][1] +
                mat_A[108][0] * mat_B[135][1] +
                mat_A[108][1] * mat_B[143][1] +
                mat_A[108][2] * mat_B[151][1] +
                mat_A[108][3] * mat_B[159][1] +
                mat_A[109][0] * mat_B[167][1] +
                mat_A[109][1] * mat_B[175][1] +
                mat_A[109][2] * mat_B[183][1] +
                mat_A[109][3] * mat_B[191][1] +
                mat_A[110][0] * mat_B[199][1] +
                mat_A[110][1] * mat_B[207][1] +
                mat_A[110][2] * mat_B[215][1] +
                mat_A[110][3] * mat_B[223][1] +
                mat_A[111][0] * mat_B[231][1] +
                mat_A[111][1] * mat_B[239][1] +
                mat_A[111][2] * mat_B[247][1] +
                mat_A[111][3] * mat_B[255][1];
    mat_C[111][2] <=
                mat_A[104][0] * mat_B[7][2] +
                mat_A[104][1] * mat_B[15][2] +
                mat_A[104][2] * mat_B[23][2] +
                mat_A[104][3] * mat_B[31][2] +
                mat_A[105][0] * mat_B[39][2] +
                mat_A[105][1] * mat_B[47][2] +
                mat_A[105][2] * mat_B[55][2] +
                mat_A[105][3] * mat_B[63][2] +
                mat_A[106][0] * mat_B[71][2] +
                mat_A[106][1] * mat_B[79][2] +
                mat_A[106][2] * mat_B[87][2] +
                mat_A[106][3] * mat_B[95][2] +
                mat_A[107][0] * mat_B[103][2] +
                mat_A[107][1] * mat_B[111][2] +
                mat_A[107][2] * mat_B[119][2] +
                mat_A[107][3] * mat_B[127][2] +
                mat_A[108][0] * mat_B[135][2] +
                mat_A[108][1] * mat_B[143][2] +
                mat_A[108][2] * mat_B[151][2] +
                mat_A[108][3] * mat_B[159][2] +
                mat_A[109][0] * mat_B[167][2] +
                mat_A[109][1] * mat_B[175][2] +
                mat_A[109][2] * mat_B[183][2] +
                mat_A[109][3] * mat_B[191][2] +
                mat_A[110][0] * mat_B[199][2] +
                mat_A[110][1] * mat_B[207][2] +
                mat_A[110][2] * mat_B[215][2] +
                mat_A[110][3] * mat_B[223][2] +
                mat_A[111][0] * mat_B[231][2] +
                mat_A[111][1] * mat_B[239][2] +
                mat_A[111][2] * mat_B[247][2] +
                mat_A[111][3] * mat_B[255][2];
    mat_C[111][3] <=
                mat_A[104][0] * mat_B[7][3] +
                mat_A[104][1] * mat_B[15][3] +
                mat_A[104][2] * mat_B[23][3] +
                mat_A[104][3] * mat_B[31][3] +
                mat_A[105][0] * mat_B[39][3] +
                mat_A[105][1] * mat_B[47][3] +
                mat_A[105][2] * mat_B[55][3] +
                mat_A[105][3] * mat_B[63][3] +
                mat_A[106][0] * mat_B[71][3] +
                mat_A[106][1] * mat_B[79][3] +
                mat_A[106][2] * mat_B[87][3] +
                mat_A[106][3] * mat_B[95][3] +
                mat_A[107][0] * mat_B[103][3] +
                mat_A[107][1] * mat_B[111][3] +
                mat_A[107][2] * mat_B[119][3] +
                mat_A[107][3] * mat_B[127][3] +
                mat_A[108][0] * mat_B[135][3] +
                mat_A[108][1] * mat_B[143][3] +
                mat_A[108][2] * mat_B[151][3] +
                mat_A[108][3] * mat_B[159][3] +
                mat_A[109][0] * mat_B[167][3] +
                mat_A[109][1] * mat_B[175][3] +
                mat_A[109][2] * mat_B[183][3] +
                mat_A[109][3] * mat_B[191][3] +
                mat_A[110][0] * mat_B[199][3] +
                mat_A[110][1] * mat_B[207][3] +
                mat_A[110][2] * mat_B[215][3] +
                mat_A[110][3] * mat_B[223][3] +
                mat_A[111][0] * mat_B[231][3] +
                mat_A[111][1] * mat_B[239][3] +
                mat_A[111][2] * mat_B[247][3] +
                mat_A[111][3] * mat_B[255][3];
    mat_C[112][0] <=
                mat_A[112][0] * mat_B[0][0] +
                mat_A[112][1] * mat_B[8][0] +
                mat_A[112][2] * mat_B[16][0] +
                mat_A[112][3] * mat_B[24][0] +
                mat_A[113][0] * mat_B[32][0] +
                mat_A[113][1] * mat_B[40][0] +
                mat_A[113][2] * mat_B[48][0] +
                mat_A[113][3] * mat_B[56][0] +
                mat_A[114][0] * mat_B[64][0] +
                mat_A[114][1] * mat_B[72][0] +
                mat_A[114][2] * mat_B[80][0] +
                mat_A[114][3] * mat_B[88][0] +
                mat_A[115][0] * mat_B[96][0] +
                mat_A[115][1] * mat_B[104][0] +
                mat_A[115][2] * mat_B[112][0] +
                mat_A[115][3] * mat_B[120][0] +
                mat_A[116][0] * mat_B[128][0] +
                mat_A[116][1] * mat_B[136][0] +
                mat_A[116][2] * mat_B[144][0] +
                mat_A[116][3] * mat_B[152][0] +
                mat_A[117][0] * mat_B[160][0] +
                mat_A[117][1] * mat_B[168][0] +
                mat_A[117][2] * mat_B[176][0] +
                mat_A[117][3] * mat_B[184][0] +
                mat_A[118][0] * mat_B[192][0] +
                mat_A[118][1] * mat_B[200][0] +
                mat_A[118][2] * mat_B[208][0] +
                mat_A[118][3] * mat_B[216][0] +
                mat_A[119][0] * mat_B[224][0] +
                mat_A[119][1] * mat_B[232][0] +
                mat_A[119][2] * mat_B[240][0] +
                mat_A[119][3] * mat_B[248][0];
    mat_C[112][1] <=
                mat_A[112][0] * mat_B[0][1] +
                mat_A[112][1] * mat_B[8][1] +
                mat_A[112][2] * mat_B[16][1] +
                mat_A[112][3] * mat_B[24][1] +
                mat_A[113][0] * mat_B[32][1] +
                mat_A[113][1] * mat_B[40][1] +
                mat_A[113][2] * mat_B[48][1] +
                mat_A[113][3] * mat_B[56][1] +
                mat_A[114][0] * mat_B[64][1] +
                mat_A[114][1] * mat_B[72][1] +
                mat_A[114][2] * mat_B[80][1] +
                mat_A[114][3] * mat_B[88][1] +
                mat_A[115][0] * mat_B[96][1] +
                mat_A[115][1] * mat_B[104][1] +
                mat_A[115][2] * mat_B[112][1] +
                mat_A[115][3] * mat_B[120][1] +
                mat_A[116][0] * mat_B[128][1] +
                mat_A[116][1] * mat_B[136][1] +
                mat_A[116][2] * mat_B[144][1] +
                mat_A[116][3] * mat_B[152][1] +
                mat_A[117][0] * mat_B[160][1] +
                mat_A[117][1] * mat_B[168][1] +
                mat_A[117][2] * mat_B[176][1] +
                mat_A[117][3] * mat_B[184][1] +
                mat_A[118][0] * mat_B[192][1] +
                mat_A[118][1] * mat_B[200][1] +
                mat_A[118][2] * mat_B[208][1] +
                mat_A[118][3] * mat_B[216][1] +
                mat_A[119][0] * mat_B[224][1] +
                mat_A[119][1] * mat_B[232][1] +
                mat_A[119][2] * mat_B[240][1] +
                mat_A[119][3] * mat_B[248][1];
    mat_C[112][2] <=
                mat_A[112][0] * mat_B[0][2] +
                mat_A[112][1] * mat_B[8][2] +
                mat_A[112][2] * mat_B[16][2] +
                mat_A[112][3] * mat_B[24][2] +
                mat_A[113][0] * mat_B[32][2] +
                mat_A[113][1] * mat_B[40][2] +
                mat_A[113][2] * mat_B[48][2] +
                mat_A[113][3] * mat_B[56][2] +
                mat_A[114][0] * mat_B[64][2] +
                mat_A[114][1] * mat_B[72][2] +
                mat_A[114][2] * mat_B[80][2] +
                mat_A[114][3] * mat_B[88][2] +
                mat_A[115][0] * mat_B[96][2] +
                mat_A[115][1] * mat_B[104][2] +
                mat_A[115][2] * mat_B[112][2] +
                mat_A[115][3] * mat_B[120][2] +
                mat_A[116][0] * mat_B[128][2] +
                mat_A[116][1] * mat_B[136][2] +
                mat_A[116][2] * mat_B[144][2] +
                mat_A[116][3] * mat_B[152][2] +
                mat_A[117][0] * mat_B[160][2] +
                mat_A[117][1] * mat_B[168][2] +
                mat_A[117][2] * mat_B[176][2] +
                mat_A[117][3] * mat_B[184][2] +
                mat_A[118][0] * mat_B[192][2] +
                mat_A[118][1] * mat_B[200][2] +
                mat_A[118][2] * mat_B[208][2] +
                mat_A[118][3] * mat_B[216][2] +
                mat_A[119][0] * mat_B[224][2] +
                mat_A[119][1] * mat_B[232][2] +
                mat_A[119][2] * mat_B[240][2] +
                mat_A[119][3] * mat_B[248][2];
    mat_C[112][3] <=
                mat_A[112][0] * mat_B[0][3] +
                mat_A[112][1] * mat_B[8][3] +
                mat_A[112][2] * mat_B[16][3] +
                mat_A[112][3] * mat_B[24][3] +
                mat_A[113][0] * mat_B[32][3] +
                mat_A[113][1] * mat_B[40][3] +
                mat_A[113][2] * mat_B[48][3] +
                mat_A[113][3] * mat_B[56][3] +
                mat_A[114][0] * mat_B[64][3] +
                mat_A[114][1] * mat_B[72][3] +
                mat_A[114][2] * mat_B[80][3] +
                mat_A[114][3] * mat_B[88][3] +
                mat_A[115][0] * mat_B[96][3] +
                mat_A[115][1] * mat_B[104][3] +
                mat_A[115][2] * mat_B[112][3] +
                mat_A[115][3] * mat_B[120][3] +
                mat_A[116][0] * mat_B[128][3] +
                mat_A[116][1] * mat_B[136][3] +
                mat_A[116][2] * mat_B[144][3] +
                mat_A[116][3] * mat_B[152][3] +
                mat_A[117][0] * mat_B[160][3] +
                mat_A[117][1] * mat_B[168][3] +
                mat_A[117][2] * mat_B[176][3] +
                mat_A[117][3] * mat_B[184][3] +
                mat_A[118][0] * mat_B[192][3] +
                mat_A[118][1] * mat_B[200][3] +
                mat_A[118][2] * mat_B[208][3] +
                mat_A[118][3] * mat_B[216][3] +
                mat_A[119][0] * mat_B[224][3] +
                mat_A[119][1] * mat_B[232][3] +
                mat_A[119][2] * mat_B[240][3] +
                mat_A[119][3] * mat_B[248][3];
    mat_C[113][0] <=
                mat_A[112][0] * mat_B[1][0] +
                mat_A[112][1] * mat_B[9][0] +
                mat_A[112][2] * mat_B[17][0] +
                mat_A[112][3] * mat_B[25][0] +
                mat_A[113][0] * mat_B[33][0] +
                mat_A[113][1] * mat_B[41][0] +
                mat_A[113][2] * mat_B[49][0] +
                mat_A[113][3] * mat_B[57][0] +
                mat_A[114][0] * mat_B[65][0] +
                mat_A[114][1] * mat_B[73][0] +
                mat_A[114][2] * mat_B[81][0] +
                mat_A[114][3] * mat_B[89][0] +
                mat_A[115][0] * mat_B[97][0] +
                mat_A[115][1] * mat_B[105][0] +
                mat_A[115][2] * mat_B[113][0] +
                mat_A[115][3] * mat_B[121][0] +
                mat_A[116][0] * mat_B[129][0] +
                mat_A[116][1] * mat_B[137][0] +
                mat_A[116][2] * mat_B[145][0] +
                mat_A[116][3] * mat_B[153][0] +
                mat_A[117][0] * mat_B[161][0] +
                mat_A[117][1] * mat_B[169][0] +
                mat_A[117][2] * mat_B[177][0] +
                mat_A[117][3] * mat_B[185][0] +
                mat_A[118][0] * mat_B[193][0] +
                mat_A[118][1] * mat_B[201][0] +
                mat_A[118][2] * mat_B[209][0] +
                mat_A[118][3] * mat_B[217][0] +
                mat_A[119][0] * mat_B[225][0] +
                mat_A[119][1] * mat_B[233][0] +
                mat_A[119][2] * mat_B[241][0] +
                mat_A[119][3] * mat_B[249][0];
    mat_C[113][1] <=
                mat_A[112][0] * mat_B[1][1] +
                mat_A[112][1] * mat_B[9][1] +
                mat_A[112][2] * mat_B[17][1] +
                mat_A[112][3] * mat_B[25][1] +
                mat_A[113][0] * mat_B[33][1] +
                mat_A[113][1] * mat_B[41][1] +
                mat_A[113][2] * mat_B[49][1] +
                mat_A[113][3] * mat_B[57][1] +
                mat_A[114][0] * mat_B[65][1] +
                mat_A[114][1] * mat_B[73][1] +
                mat_A[114][2] * mat_B[81][1] +
                mat_A[114][3] * mat_B[89][1] +
                mat_A[115][0] * mat_B[97][1] +
                mat_A[115][1] * mat_B[105][1] +
                mat_A[115][2] * mat_B[113][1] +
                mat_A[115][3] * mat_B[121][1] +
                mat_A[116][0] * mat_B[129][1] +
                mat_A[116][1] * mat_B[137][1] +
                mat_A[116][2] * mat_B[145][1] +
                mat_A[116][3] * mat_B[153][1] +
                mat_A[117][0] * mat_B[161][1] +
                mat_A[117][1] * mat_B[169][1] +
                mat_A[117][2] * mat_B[177][1] +
                mat_A[117][3] * mat_B[185][1] +
                mat_A[118][0] * mat_B[193][1] +
                mat_A[118][1] * mat_B[201][1] +
                mat_A[118][2] * mat_B[209][1] +
                mat_A[118][3] * mat_B[217][1] +
                mat_A[119][0] * mat_B[225][1] +
                mat_A[119][1] * mat_B[233][1] +
                mat_A[119][2] * mat_B[241][1] +
                mat_A[119][3] * mat_B[249][1];
    mat_C[113][2] <=
                mat_A[112][0] * mat_B[1][2] +
                mat_A[112][1] * mat_B[9][2] +
                mat_A[112][2] * mat_B[17][2] +
                mat_A[112][3] * mat_B[25][2] +
                mat_A[113][0] * mat_B[33][2] +
                mat_A[113][1] * mat_B[41][2] +
                mat_A[113][2] * mat_B[49][2] +
                mat_A[113][3] * mat_B[57][2] +
                mat_A[114][0] * mat_B[65][2] +
                mat_A[114][1] * mat_B[73][2] +
                mat_A[114][2] * mat_B[81][2] +
                mat_A[114][3] * mat_B[89][2] +
                mat_A[115][0] * mat_B[97][2] +
                mat_A[115][1] * mat_B[105][2] +
                mat_A[115][2] * mat_B[113][2] +
                mat_A[115][3] * mat_B[121][2] +
                mat_A[116][0] * mat_B[129][2] +
                mat_A[116][1] * mat_B[137][2] +
                mat_A[116][2] * mat_B[145][2] +
                mat_A[116][3] * mat_B[153][2] +
                mat_A[117][0] * mat_B[161][2] +
                mat_A[117][1] * mat_B[169][2] +
                mat_A[117][2] * mat_B[177][2] +
                mat_A[117][3] * mat_B[185][2] +
                mat_A[118][0] * mat_B[193][2] +
                mat_A[118][1] * mat_B[201][2] +
                mat_A[118][2] * mat_B[209][2] +
                mat_A[118][3] * mat_B[217][2] +
                mat_A[119][0] * mat_B[225][2] +
                mat_A[119][1] * mat_B[233][2] +
                mat_A[119][2] * mat_B[241][2] +
                mat_A[119][3] * mat_B[249][2];
    mat_C[113][3] <=
                mat_A[112][0] * mat_B[1][3] +
                mat_A[112][1] * mat_B[9][3] +
                mat_A[112][2] * mat_B[17][3] +
                mat_A[112][3] * mat_B[25][3] +
                mat_A[113][0] * mat_B[33][3] +
                mat_A[113][1] * mat_B[41][3] +
                mat_A[113][2] * mat_B[49][3] +
                mat_A[113][3] * mat_B[57][3] +
                mat_A[114][0] * mat_B[65][3] +
                mat_A[114][1] * mat_B[73][3] +
                mat_A[114][2] * mat_B[81][3] +
                mat_A[114][3] * mat_B[89][3] +
                mat_A[115][0] * mat_B[97][3] +
                mat_A[115][1] * mat_B[105][3] +
                mat_A[115][2] * mat_B[113][3] +
                mat_A[115][3] * mat_B[121][3] +
                mat_A[116][0] * mat_B[129][3] +
                mat_A[116][1] * mat_B[137][3] +
                mat_A[116][2] * mat_B[145][3] +
                mat_A[116][3] * mat_B[153][3] +
                mat_A[117][0] * mat_B[161][3] +
                mat_A[117][1] * mat_B[169][3] +
                mat_A[117][2] * mat_B[177][3] +
                mat_A[117][3] * mat_B[185][3] +
                mat_A[118][0] * mat_B[193][3] +
                mat_A[118][1] * mat_B[201][3] +
                mat_A[118][2] * mat_B[209][3] +
                mat_A[118][3] * mat_B[217][3] +
                mat_A[119][0] * mat_B[225][3] +
                mat_A[119][1] * mat_B[233][3] +
                mat_A[119][2] * mat_B[241][3] +
                mat_A[119][3] * mat_B[249][3];
    mat_C[114][0] <=
                mat_A[112][0] * mat_B[2][0] +
                mat_A[112][1] * mat_B[10][0] +
                mat_A[112][2] * mat_B[18][0] +
                mat_A[112][3] * mat_B[26][0] +
                mat_A[113][0] * mat_B[34][0] +
                mat_A[113][1] * mat_B[42][0] +
                mat_A[113][2] * mat_B[50][0] +
                mat_A[113][3] * mat_B[58][0] +
                mat_A[114][0] * mat_B[66][0] +
                mat_A[114][1] * mat_B[74][0] +
                mat_A[114][2] * mat_B[82][0] +
                mat_A[114][3] * mat_B[90][0] +
                mat_A[115][0] * mat_B[98][0] +
                mat_A[115][1] * mat_B[106][0] +
                mat_A[115][2] * mat_B[114][0] +
                mat_A[115][3] * mat_B[122][0] +
                mat_A[116][0] * mat_B[130][0] +
                mat_A[116][1] * mat_B[138][0] +
                mat_A[116][2] * mat_B[146][0] +
                mat_A[116][3] * mat_B[154][0] +
                mat_A[117][0] * mat_B[162][0] +
                mat_A[117][1] * mat_B[170][0] +
                mat_A[117][2] * mat_B[178][0] +
                mat_A[117][3] * mat_B[186][0] +
                mat_A[118][0] * mat_B[194][0] +
                mat_A[118][1] * mat_B[202][0] +
                mat_A[118][2] * mat_B[210][0] +
                mat_A[118][3] * mat_B[218][0] +
                mat_A[119][0] * mat_B[226][0] +
                mat_A[119][1] * mat_B[234][0] +
                mat_A[119][2] * mat_B[242][0] +
                mat_A[119][3] * mat_B[250][0];
    mat_C[114][1] <=
                mat_A[112][0] * mat_B[2][1] +
                mat_A[112][1] * mat_B[10][1] +
                mat_A[112][2] * mat_B[18][1] +
                mat_A[112][3] * mat_B[26][1] +
                mat_A[113][0] * mat_B[34][1] +
                mat_A[113][1] * mat_B[42][1] +
                mat_A[113][2] * mat_B[50][1] +
                mat_A[113][3] * mat_B[58][1] +
                mat_A[114][0] * mat_B[66][1] +
                mat_A[114][1] * mat_B[74][1] +
                mat_A[114][2] * mat_B[82][1] +
                mat_A[114][3] * mat_B[90][1] +
                mat_A[115][0] * mat_B[98][1] +
                mat_A[115][1] * mat_B[106][1] +
                mat_A[115][2] * mat_B[114][1] +
                mat_A[115][3] * mat_B[122][1] +
                mat_A[116][0] * mat_B[130][1] +
                mat_A[116][1] * mat_B[138][1] +
                mat_A[116][2] * mat_B[146][1] +
                mat_A[116][3] * mat_B[154][1] +
                mat_A[117][0] * mat_B[162][1] +
                mat_A[117][1] * mat_B[170][1] +
                mat_A[117][2] * mat_B[178][1] +
                mat_A[117][3] * mat_B[186][1] +
                mat_A[118][0] * mat_B[194][1] +
                mat_A[118][1] * mat_B[202][1] +
                mat_A[118][2] * mat_B[210][1] +
                mat_A[118][3] * mat_B[218][1] +
                mat_A[119][0] * mat_B[226][1] +
                mat_A[119][1] * mat_B[234][1] +
                mat_A[119][2] * mat_B[242][1] +
                mat_A[119][3] * mat_B[250][1];
    mat_C[114][2] <=
                mat_A[112][0] * mat_B[2][2] +
                mat_A[112][1] * mat_B[10][2] +
                mat_A[112][2] * mat_B[18][2] +
                mat_A[112][3] * mat_B[26][2] +
                mat_A[113][0] * mat_B[34][2] +
                mat_A[113][1] * mat_B[42][2] +
                mat_A[113][2] * mat_B[50][2] +
                mat_A[113][3] * mat_B[58][2] +
                mat_A[114][0] * mat_B[66][2] +
                mat_A[114][1] * mat_B[74][2] +
                mat_A[114][2] * mat_B[82][2] +
                mat_A[114][3] * mat_B[90][2] +
                mat_A[115][0] * mat_B[98][2] +
                mat_A[115][1] * mat_B[106][2] +
                mat_A[115][2] * mat_B[114][2] +
                mat_A[115][3] * mat_B[122][2] +
                mat_A[116][0] * mat_B[130][2] +
                mat_A[116][1] * mat_B[138][2] +
                mat_A[116][2] * mat_B[146][2] +
                mat_A[116][3] * mat_B[154][2] +
                mat_A[117][0] * mat_B[162][2] +
                mat_A[117][1] * mat_B[170][2] +
                mat_A[117][2] * mat_B[178][2] +
                mat_A[117][3] * mat_B[186][2] +
                mat_A[118][0] * mat_B[194][2] +
                mat_A[118][1] * mat_B[202][2] +
                mat_A[118][2] * mat_B[210][2] +
                mat_A[118][3] * mat_B[218][2] +
                mat_A[119][0] * mat_B[226][2] +
                mat_A[119][1] * mat_B[234][2] +
                mat_A[119][2] * mat_B[242][2] +
                mat_A[119][3] * mat_B[250][2];
    mat_C[114][3] <=
                mat_A[112][0] * mat_B[2][3] +
                mat_A[112][1] * mat_B[10][3] +
                mat_A[112][2] * mat_B[18][3] +
                mat_A[112][3] * mat_B[26][3] +
                mat_A[113][0] * mat_B[34][3] +
                mat_A[113][1] * mat_B[42][3] +
                mat_A[113][2] * mat_B[50][3] +
                mat_A[113][3] * mat_B[58][3] +
                mat_A[114][0] * mat_B[66][3] +
                mat_A[114][1] * mat_B[74][3] +
                mat_A[114][2] * mat_B[82][3] +
                mat_A[114][3] * mat_B[90][3] +
                mat_A[115][0] * mat_B[98][3] +
                mat_A[115][1] * mat_B[106][3] +
                mat_A[115][2] * mat_B[114][3] +
                mat_A[115][3] * mat_B[122][3] +
                mat_A[116][0] * mat_B[130][3] +
                mat_A[116][1] * mat_B[138][3] +
                mat_A[116][2] * mat_B[146][3] +
                mat_A[116][3] * mat_B[154][3] +
                mat_A[117][0] * mat_B[162][3] +
                mat_A[117][1] * mat_B[170][3] +
                mat_A[117][2] * mat_B[178][3] +
                mat_A[117][3] * mat_B[186][3] +
                mat_A[118][0] * mat_B[194][3] +
                mat_A[118][1] * mat_B[202][3] +
                mat_A[118][2] * mat_B[210][3] +
                mat_A[118][3] * mat_B[218][3] +
                mat_A[119][0] * mat_B[226][3] +
                mat_A[119][1] * mat_B[234][3] +
                mat_A[119][2] * mat_B[242][3] +
                mat_A[119][3] * mat_B[250][3];
    mat_C[115][0] <=
                mat_A[112][0] * mat_B[3][0] +
                mat_A[112][1] * mat_B[11][0] +
                mat_A[112][2] * mat_B[19][0] +
                mat_A[112][3] * mat_B[27][0] +
                mat_A[113][0] * mat_B[35][0] +
                mat_A[113][1] * mat_B[43][0] +
                mat_A[113][2] * mat_B[51][0] +
                mat_A[113][3] * mat_B[59][0] +
                mat_A[114][0] * mat_B[67][0] +
                mat_A[114][1] * mat_B[75][0] +
                mat_A[114][2] * mat_B[83][0] +
                mat_A[114][3] * mat_B[91][0] +
                mat_A[115][0] * mat_B[99][0] +
                mat_A[115][1] * mat_B[107][0] +
                mat_A[115][2] * mat_B[115][0] +
                mat_A[115][3] * mat_B[123][0] +
                mat_A[116][0] * mat_B[131][0] +
                mat_A[116][1] * mat_B[139][0] +
                mat_A[116][2] * mat_B[147][0] +
                mat_A[116][3] * mat_B[155][0] +
                mat_A[117][0] * mat_B[163][0] +
                mat_A[117][1] * mat_B[171][0] +
                mat_A[117][2] * mat_B[179][0] +
                mat_A[117][3] * mat_B[187][0] +
                mat_A[118][0] * mat_B[195][0] +
                mat_A[118][1] * mat_B[203][0] +
                mat_A[118][2] * mat_B[211][0] +
                mat_A[118][3] * mat_B[219][0] +
                mat_A[119][0] * mat_B[227][0] +
                mat_A[119][1] * mat_B[235][0] +
                mat_A[119][2] * mat_B[243][0] +
                mat_A[119][3] * mat_B[251][0];
    mat_C[115][1] <=
                mat_A[112][0] * mat_B[3][1] +
                mat_A[112][1] * mat_B[11][1] +
                mat_A[112][2] * mat_B[19][1] +
                mat_A[112][3] * mat_B[27][1] +
                mat_A[113][0] * mat_B[35][1] +
                mat_A[113][1] * mat_B[43][1] +
                mat_A[113][2] * mat_B[51][1] +
                mat_A[113][3] * mat_B[59][1] +
                mat_A[114][0] * mat_B[67][1] +
                mat_A[114][1] * mat_B[75][1] +
                mat_A[114][2] * mat_B[83][1] +
                mat_A[114][3] * mat_B[91][1] +
                mat_A[115][0] * mat_B[99][1] +
                mat_A[115][1] * mat_B[107][1] +
                mat_A[115][2] * mat_B[115][1] +
                mat_A[115][3] * mat_B[123][1] +
                mat_A[116][0] * mat_B[131][1] +
                mat_A[116][1] * mat_B[139][1] +
                mat_A[116][2] * mat_B[147][1] +
                mat_A[116][3] * mat_B[155][1] +
                mat_A[117][0] * mat_B[163][1] +
                mat_A[117][1] * mat_B[171][1] +
                mat_A[117][2] * mat_B[179][1] +
                mat_A[117][3] * mat_B[187][1] +
                mat_A[118][0] * mat_B[195][1] +
                mat_A[118][1] * mat_B[203][1] +
                mat_A[118][2] * mat_B[211][1] +
                mat_A[118][3] * mat_B[219][1] +
                mat_A[119][0] * mat_B[227][1] +
                mat_A[119][1] * mat_B[235][1] +
                mat_A[119][2] * mat_B[243][1] +
                mat_A[119][3] * mat_B[251][1];
    mat_C[115][2] <=
                mat_A[112][0] * mat_B[3][2] +
                mat_A[112][1] * mat_B[11][2] +
                mat_A[112][2] * mat_B[19][2] +
                mat_A[112][3] * mat_B[27][2] +
                mat_A[113][0] * mat_B[35][2] +
                mat_A[113][1] * mat_B[43][2] +
                mat_A[113][2] * mat_B[51][2] +
                mat_A[113][3] * mat_B[59][2] +
                mat_A[114][0] * mat_B[67][2] +
                mat_A[114][1] * mat_B[75][2] +
                mat_A[114][2] * mat_B[83][2] +
                mat_A[114][3] * mat_B[91][2] +
                mat_A[115][0] * mat_B[99][2] +
                mat_A[115][1] * mat_B[107][2] +
                mat_A[115][2] * mat_B[115][2] +
                mat_A[115][3] * mat_B[123][2] +
                mat_A[116][0] * mat_B[131][2] +
                mat_A[116][1] * mat_B[139][2] +
                mat_A[116][2] * mat_B[147][2] +
                mat_A[116][3] * mat_B[155][2] +
                mat_A[117][0] * mat_B[163][2] +
                mat_A[117][1] * mat_B[171][2] +
                mat_A[117][2] * mat_B[179][2] +
                mat_A[117][3] * mat_B[187][2] +
                mat_A[118][0] * mat_B[195][2] +
                mat_A[118][1] * mat_B[203][2] +
                mat_A[118][2] * mat_B[211][2] +
                mat_A[118][3] * mat_B[219][2] +
                mat_A[119][0] * mat_B[227][2] +
                mat_A[119][1] * mat_B[235][2] +
                mat_A[119][2] * mat_B[243][2] +
                mat_A[119][3] * mat_B[251][2];
    mat_C[115][3] <=
                mat_A[112][0] * mat_B[3][3] +
                mat_A[112][1] * mat_B[11][3] +
                mat_A[112][2] * mat_B[19][3] +
                mat_A[112][3] * mat_B[27][3] +
                mat_A[113][0] * mat_B[35][3] +
                mat_A[113][1] * mat_B[43][3] +
                mat_A[113][2] * mat_B[51][3] +
                mat_A[113][3] * mat_B[59][3] +
                mat_A[114][0] * mat_B[67][3] +
                mat_A[114][1] * mat_B[75][3] +
                mat_A[114][2] * mat_B[83][3] +
                mat_A[114][3] * mat_B[91][3] +
                mat_A[115][0] * mat_B[99][3] +
                mat_A[115][1] * mat_B[107][3] +
                mat_A[115][2] * mat_B[115][3] +
                mat_A[115][3] * mat_B[123][3] +
                mat_A[116][0] * mat_B[131][3] +
                mat_A[116][1] * mat_B[139][3] +
                mat_A[116][2] * mat_B[147][3] +
                mat_A[116][3] * mat_B[155][3] +
                mat_A[117][0] * mat_B[163][3] +
                mat_A[117][1] * mat_B[171][3] +
                mat_A[117][2] * mat_B[179][3] +
                mat_A[117][3] * mat_B[187][3] +
                mat_A[118][0] * mat_B[195][3] +
                mat_A[118][1] * mat_B[203][3] +
                mat_A[118][2] * mat_B[211][3] +
                mat_A[118][3] * mat_B[219][3] +
                mat_A[119][0] * mat_B[227][3] +
                mat_A[119][1] * mat_B[235][3] +
                mat_A[119][2] * mat_B[243][3] +
                mat_A[119][3] * mat_B[251][3];
    mat_C[116][0] <=
                mat_A[112][0] * mat_B[4][0] +
                mat_A[112][1] * mat_B[12][0] +
                mat_A[112][2] * mat_B[20][0] +
                mat_A[112][3] * mat_B[28][0] +
                mat_A[113][0] * mat_B[36][0] +
                mat_A[113][1] * mat_B[44][0] +
                mat_A[113][2] * mat_B[52][0] +
                mat_A[113][3] * mat_B[60][0] +
                mat_A[114][0] * mat_B[68][0] +
                mat_A[114][1] * mat_B[76][0] +
                mat_A[114][2] * mat_B[84][0] +
                mat_A[114][3] * mat_B[92][0] +
                mat_A[115][0] * mat_B[100][0] +
                mat_A[115][1] * mat_B[108][0] +
                mat_A[115][2] * mat_B[116][0] +
                mat_A[115][3] * mat_B[124][0] +
                mat_A[116][0] * mat_B[132][0] +
                mat_A[116][1] * mat_B[140][0] +
                mat_A[116][2] * mat_B[148][0] +
                mat_A[116][3] * mat_B[156][0] +
                mat_A[117][0] * mat_B[164][0] +
                mat_A[117][1] * mat_B[172][0] +
                mat_A[117][2] * mat_B[180][0] +
                mat_A[117][3] * mat_B[188][0] +
                mat_A[118][0] * mat_B[196][0] +
                mat_A[118][1] * mat_B[204][0] +
                mat_A[118][2] * mat_B[212][0] +
                mat_A[118][3] * mat_B[220][0] +
                mat_A[119][0] * mat_B[228][0] +
                mat_A[119][1] * mat_B[236][0] +
                mat_A[119][2] * mat_B[244][0] +
                mat_A[119][3] * mat_B[252][0];
    mat_C[116][1] <=
                mat_A[112][0] * mat_B[4][1] +
                mat_A[112][1] * mat_B[12][1] +
                mat_A[112][2] * mat_B[20][1] +
                mat_A[112][3] * mat_B[28][1] +
                mat_A[113][0] * mat_B[36][1] +
                mat_A[113][1] * mat_B[44][1] +
                mat_A[113][2] * mat_B[52][1] +
                mat_A[113][3] * mat_B[60][1] +
                mat_A[114][0] * mat_B[68][1] +
                mat_A[114][1] * mat_B[76][1] +
                mat_A[114][2] * mat_B[84][1] +
                mat_A[114][3] * mat_B[92][1] +
                mat_A[115][0] * mat_B[100][1] +
                mat_A[115][1] * mat_B[108][1] +
                mat_A[115][2] * mat_B[116][1] +
                mat_A[115][3] * mat_B[124][1] +
                mat_A[116][0] * mat_B[132][1] +
                mat_A[116][1] * mat_B[140][1] +
                mat_A[116][2] * mat_B[148][1] +
                mat_A[116][3] * mat_B[156][1] +
                mat_A[117][0] * mat_B[164][1] +
                mat_A[117][1] * mat_B[172][1] +
                mat_A[117][2] * mat_B[180][1] +
                mat_A[117][3] * mat_B[188][1] +
                mat_A[118][0] * mat_B[196][1] +
                mat_A[118][1] * mat_B[204][1] +
                mat_A[118][2] * mat_B[212][1] +
                mat_A[118][3] * mat_B[220][1] +
                mat_A[119][0] * mat_B[228][1] +
                mat_A[119][1] * mat_B[236][1] +
                mat_A[119][2] * mat_B[244][1] +
                mat_A[119][3] * mat_B[252][1];
    mat_C[116][2] <=
                mat_A[112][0] * mat_B[4][2] +
                mat_A[112][1] * mat_B[12][2] +
                mat_A[112][2] * mat_B[20][2] +
                mat_A[112][3] * mat_B[28][2] +
                mat_A[113][0] * mat_B[36][2] +
                mat_A[113][1] * mat_B[44][2] +
                mat_A[113][2] * mat_B[52][2] +
                mat_A[113][3] * mat_B[60][2] +
                mat_A[114][0] * mat_B[68][2] +
                mat_A[114][1] * mat_B[76][2] +
                mat_A[114][2] * mat_B[84][2] +
                mat_A[114][3] * mat_B[92][2] +
                mat_A[115][0] * mat_B[100][2] +
                mat_A[115][1] * mat_B[108][2] +
                mat_A[115][2] * mat_B[116][2] +
                mat_A[115][3] * mat_B[124][2] +
                mat_A[116][0] * mat_B[132][2] +
                mat_A[116][1] * mat_B[140][2] +
                mat_A[116][2] * mat_B[148][2] +
                mat_A[116][3] * mat_B[156][2] +
                mat_A[117][0] * mat_B[164][2] +
                mat_A[117][1] * mat_B[172][2] +
                mat_A[117][2] * mat_B[180][2] +
                mat_A[117][3] * mat_B[188][2] +
                mat_A[118][0] * mat_B[196][2] +
                mat_A[118][1] * mat_B[204][2] +
                mat_A[118][2] * mat_B[212][2] +
                mat_A[118][3] * mat_B[220][2] +
                mat_A[119][0] * mat_B[228][2] +
                mat_A[119][1] * mat_B[236][2] +
                mat_A[119][2] * mat_B[244][2] +
                mat_A[119][3] * mat_B[252][2];
    mat_C[116][3] <=
                mat_A[112][0] * mat_B[4][3] +
                mat_A[112][1] * mat_B[12][3] +
                mat_A[112][2] * mat_B[20][3] +
                mat_A[112][3] * mat_B[28][3] +
                mat_A[113][0] * mat_B[36][3] +
                mat_A[113][1] * mat_B[44][3] +
                mat_A[113][2] * mat_B[52][3] +
                mat_A[113][3] * mat_B[60][3] +
                mat_A[114][0] * mat_B[68][3] +
                mat_A[114][1] * mat_B[76][3] +
                mat_A[114][2] * mat_B[84][3] +
                mat_A[114][3] * mat_B[92][3] +
                mat_A[115][0] * mat_B[100][3] +
                mat_A[115][1] * mat_B[108][3] +
                mat_A[115][2] * mat_B[116][3] +
                mat_A[115][3] * mat_B[124][3] +
                mat_A[116][0] * mat_B[132][3] +
                mat_A[116][1] * mat_B[140][3] +
                mat_A[116][2] * mat_B[148][3] +
                mat_A[116][3] * mat_B[156][3] +
                mat_A[117][0] * mat_B[164][3] +
                mat_A[117][1] * mat_B[172][3] +
                mat_A[117][2] * mat_B[180][3] +
                mat_A[117][3] * mat_B[188][3] +
                mat_A[118][0] * mat_B[196][3] +
                mat_A[118][1] * mat_B[204][3] +
                mat_A[118][2] * mat_B[212][3] +
                mat_A[118][3] * mat_B[220][3] +
                mat_A[119][0] * mat_B[228][3] +
                mat_A[119][1] * mat_B[236][3] +
                mat_A[119][2] * mat_B[244][3] +
                mat_A[119][3] * mat_B[252][3];
    mat_C[117][0] <=
                mat_A[112][0] * mat_B[5][0] +
                mat_A[112][1] * mat_B[13][0] +
                mat_A[112][2] * mat_B[21][0] +
                mat_A[112][3] * mat_B[29][0] +
                mat_A[113][0] * mat_B[37][0] +
                mat_A[113][1] * mat_B[45][0] +
                mat_A[113][2] * mat_B[53][0] +
                mat_A[113][3] * mat_B[61][0] +
                mat_A[114][0] * mat_B[69][0] +
                mat_A[114][1] * mat_B[77][0] +
                mat_A[114][2] * mat_B[85][0] +
                mat_A[114][3] * mat_B[93][0] +
                mat_A[115][0] * mat_B[101][0] +
                mat_A[115][1] * mat_B[109][0] +
                mat_A[115][2] * mat_B[117][0] +
                mat_A[115][3] * mat_B[125][0] +
                mat_A[116][0] * mat_B[133][0] +
                mat_A[116][1] * mat_B[141][0] +
                mat_A[116][2] * mat_B[149][0] +
                mat_A[116][3] * mat_B[157][0] +
                mat_A[117][0] * mat_B[165][0] +
                mat_A[117][1] * mat_B[173][0] +
                mat_A[117][2] * mat_B[181][0] +
                mat_A[117][3] * mat_B[189][0] +
                mat_A[118][0] * mat_B[197][0] +
                mat_A[118][1] * mat_B[205][0] +
                mat_A[118][2] * mat_B[213][0] +
                mat_A[118][3] * mat_B[221][0] +
                mat_A[119][0] * mat_B[229][0] +
                mat_A[119][1] * mat_B[237][0] +
                mat_A[119][2] * mat_B[245][0] +
                mat_A[119][3] * mat_B[253][0];
    mat_C[117][1] <=
                mat_A[112][0] * mat_B[5][1] +
                mat_A[112][1] * mat_B[13][1] +
                mat_A[112][2] * mat_B[21][1] +
                mat_A[112][3] * mat_B[29][1] +
                mat_A[113][0] * mat_B[37][1] +
                mat_A[113][1] * mat_B[45][1] +
                mat_A[113][2] * mat_B[53][1] +
                mat_A[113][3] * mat_B[61][1] +
                mat_A[114][0] * mat_B[69][1] +
                mat_A[114][1] * mat_B[77][1] +
                mat_A[114][2] * mat_B[85][1] +
                mat_A[114][3] * mat_B[93][1] +
                mat_A[115][0] * mat_B[101][1] +
                mat_A[115][1] * mat_B[109][1] +
                mat_A[115][2] * mat_B[117][1] +
                mat_A[115][3] * mat_B[125][1] +
                mat_A[116][0] * mat_B[133][1] +
                mat_A[116][1] * mat_B[141][1] +
                mat_A[116][2] * mat_B[149][1] +
                mat_A[116][3] * mat_B[157][1] +
                mat_A[117][0] * mat_B[165][1] +
                mat_A[117][1] * mat_B[173][1] +
                mat_A[117][2] * mat_B[181][1] +
                mat_A[117][3] * mat_B[189][1] +
                mat_A[118][0] * mat_B[197][1] +
                mat_A[118][1] * mat_B[205][1] +
                mat_A[118][2] * mat_B[213][1] +
                mat_A[118][3] * mat_B[221][1] +
                mat_A[119][0] * mat_B[229][1] +
                mat_A[119][1] * mat_B[237][1] +
                mat_A[119][2] * mat_B[245][1] +
                mat_A[119][3] * mat_B[253][1];
    mat_C[117][2] <=
                mat_A[112][0] * mat_B[5][2] +
                mat_A[112][1] * mat_B[13][2] +
                mat_A[112][2] * mat_B[21][2] +
                mat_A[112][3] * mat_B[29][2] +
                mat_A[113][0] * mat_B[37][2] +
                mat_A[113][1] * mat_B[45][2] +
                mat_A[113][2] * mat_B[53][2] +
                mat_A[113][3] * mat_B[61][2] +
                mat_A[114][0] * mat_B[69][2] +
                mat_A[114][1] * mat_B[77][2] +
                mat_A[114][2] * mat_B[85][2] +
                mat_A[114][3] * mat_B[93][2] +
                mat_A[115][0] * mat_B[101][2] +
                mat_A[115][1] * mat_B[109][2] +
                mat_A[115][2] * mat_B[117][2] +
                mat_A[115][3] * mat_B[125][2] +
                mat_A[116][0] * mat_B[133][2] +
                mat_A[116][1] * mat_B[141][2] +
                mat_A[116][2] * mat_B[149][2] +
                mat_A[116][3] * mat_B[157][2] +
                mat_A[117][0] * mat_B[165][2] +
                mat_A[117][1] * mat_B[173][2] +
                mat_A[117][2] * mat_B[181][2] +
                mat_A[117][3] * mat_B[189][2] +
                mat_A[118][0] * mat_B[197][2] +
                mat_A[118][1] * mat_B[205][2] +
                mat_A[118][2] * mat_B[213][2] +
                mat_A[118][3] * mat_B[221][2] +
                mat_A[119][0] * mat_B[229][2] +
                mat_A[119][1] * mat_B[237][2] +
                mat_A[119][2] * mat_B[245][2] +
                mat_A[119][3] * mat_B[253][2];
    mat_C[117][3] <=
                mat_A[112][0] * mat_B[5][3] +
                mat_A[112][1] * mat_B[13][3] +
                mat_A[112][2] * mat_B[21][3] +
                mat_A[112][3] * mat_B[29][3] +
                mat_A[113][0] * mat_B[37][3] +
                mat_A[113][1] * mat_B[45][3] +
                mat_A[113][2] * mat_B[53][3] +
                mat_A[113][3] * mat_B[61][3] +
                mat_A[114][0] * mat_B[69][3] +
                mat_A[114][1] * mat_B[77][3] +
                mat_A[114][2] * mat_B[85][3] +
                mat_A[114][3] * mat_B[93][3] +
                mat_A[115][0] * mat_B[101][3] +
                mat_A[115][1] * mat_B[109][3] +
                mat_A[115][2] * mat_B[117][3] +
                mat_A[115][3] * mat_B[125][3] +
                mat_A[116][0] * mat_B[133][3] +
                mat_A[116][1] * mat_B[141][3] +
                mat_A[116][2] * mat_B[149][3] +
                mat_A[116][3] * mat_B[157][3] +
                mat_A[117][0] * mat_B[165][3] +
                mat_A[117][1] * mat_B[173][3] +
                mat_A[117][2] * mat_B[181][3] +
                mat_A[117][3] * mat_B[189][3] +
                mat_A[118][0] * mat_B[197][3] +
                mat_A[118][1] * mat_B[205][3] +
                mat_A[118][2] * mat_B[213][3] +
                mat_A[118][3] * mat_B[221][3] +
                mat_A[119][0] * mat_B[229][3] +
                mat_A[119][1] * mat_B[237][3] +
                mat_A[119][2] * mat_B[245][3] +
                mat_A[119][3] * mat_B[253][3];
    mat_C[118][0] <=
                mat_A[112][0] * mat_B[6][0] +
                mat_A[112][1] * mat_B[14][0] +
                mat_A[112][2] * mat_B[22][0] +
                mat_A[112][3] * mat_B[30][0] +
                mat_A[113][0] * mat_B[38][0] +
                mat_A[113][1] * mat_B[46][0] +
                mat_A[113][2] * mat_B[54][0] +
                mat_A[113][3] * mat_B[62][0] +
                mat_A[114][0] * mat_B[70][0] +
                mat_A[114][1] * mat_B[78][0] +
                mat_A[114][2] * mat_B[86][0] +
                mat_A[114][3] * mat_B[94][0] +
                mat_A[115][0] * mat_B[102][0] +
                mat_A[115][1] * mat_B[110][0] +
                mat_A[115][2] * mat_B[118][0] +
                mat_A[115][3] * mat_B[126][0] +
                mat_A[116][0] * mat_B[134][0] +
                mat_A[116][1] * mat_B[142][0] +
                mat_A[116][2] * mat_B[150][0] +
                mat_A[116][3] * mat_B[158][0] +
                mat_A[117][0] * mat_B[166][0] +
                mat_A[117][1] * mat_B[174][0] +
                mat_A[117][2] * mat_B[182][0] +
                mat_A[117][3] * mat_B[190][0] +
                mat_A[118][0] * mat_B[198][0] +
                mat_A[118][1] * mat_B[206][0] +
                mat_A[118][2] * mat_B[214][0] +
                mat_A[118][3] * mat_B[222][0] +
                mat_A[119][0] * mat_B[230][0] +
                mat_A[119][1] * mat_B[238][0] +
                mat_A[119][2] * mat_B[246][0] +
                mat_A[119][3] * mat_B[254][0];
    mat_C[118][1] <=
                mat_A[112][0] * mat_B[6][1] +
                mat_A[112][1] * mat_B[14][1] +
                mat_A[112][2] * mat_B[22][1] +
                mat_A[112][3] * mat_B[30][1] +
                mat_A[113][0] * mat_B[38][1] +
                mat_A[113][1] * mat_B[46][1] +
                mat_A[113][2] * mat_B[54][1] +
                mat_A[113][3] * mat_B[62][1] +
                mat_A[114][0] * mat_B[70][1] +
                mat_A[114][1] * mat_B[78][1] +
                mat_A[114][2] * mat_B[86][1] +
                mat_A[114][3] * mat_B[94][1] +
                mat_A[115][0] * mat_B[102][1] +
                mat_A[115][1] * mat_B[110][1] +
                mat_A[115][2] * mat_B[118][1] +
                mat_A[115][3] * mat_B[126][1] +
                mat_A[116][0] * mat_B[134][1] +
                mat_A[116][1] * mat_B[142][1] +
                mat_A[116][2] * mat_B[150][1] +
                mat_A[116][3] * mat_B[158][1] +
                mat_A[117][0] * mat_B[166][1] +
                mat_A[117][1] * mat_B[174][1] +
                mat_A[117][2] * mat_B[182][1] +
                mat_A[117][3] * mat_B[190][1] +
                mat_A[118][0] * mat_B[198][1] +
                mat_A[118][1] * mat_B[206][1] +
                mat_A[118][2] * mat_B[214][1] +
                mat_A[118][3] * mat_B[222][1] +
                mat_A[119][0] * mat_B[230][1] +
                mat_A[119][1] * mat_B[238][1] +
                mat_A[119][2] * mat_B[246][1] +
                mat_A[119][3] * mat_B[254][1];
    mat_C[118][2] <=
                mat_A[112][0] * mat_B[6][2] +
                mat_A[112][1] * mat_B[14][2] +
                mat_A[112][2] * mat_B[22][2] +
                mat_A[112][3] * mat_B[30][2] +
                mat_A[113][0] * mat_B[38][2] +
                mat_A[113][1] * mat_B[46][2] +
                mat_A[113][2] * mat_B[54][2] +
                mat_A[113][3] * mat_B[62][2] +
                mat_A[114][0] * mat_B[70][2] +
                mat_A[114][1] * mat_B[78][2] +
                mat_A[114][2] * mat_B[86][2] +
                mat_A[114][3] * mat_B[94][2] +
                mat_A[115][0] * mat_B[102][2] +
                mat_A[115][1] * mat_B[110][2] +
                mat_A[115][2] * mat_B[118][2] +
                mat_A[115][3] * mat_B[126][2] +
                mat_A[116][0] * mat_B[134][2] +
                mat_A[116][1] * mat_B[142][2] +
                mat_A[116][2] * mat_B[150][2] +
                mat_A[116][3] * mat_B[158][2] +
                mat_A[117][0] * mat_B[166][2] +
                mat_A[117][1] * mat_B[174][2] +
                mat_A[117][2] * mat_B[182][2] +
                mat_A[117][3] * mat_B[190][2] +
                mat_A[118][0] * mat_B[198][2] +
                mat_A[118][1] * mat_B[206][2] +
                mat_A[118][2] * mat_B[214][2] +
                mat_A[118][3] * mat_B[222][2] +
                mat_A[119][0] * mat_B[230][2] +
                mat_A[119][1] * mat_B[238][2] +
                mat_A[119][2] * mat_B[246][2] +
                mat_A[119][3] * mat_B[254][2];
    mat_C[118][3] <=
                mat_A[112][0] * mat_B[6][3] +
                mat_A[112][1] * mat_B[14][3] +
                mat_A[112][2] * mat_B[22][3] +
                mat_A[112][3] * mat_B[30][3] +
                mat_A[113][0] * mat_B[38][3] +
                mat_A[113][1] * mat_B[46][3] +
                mat_A[113][2] * mat_B[54][3] +
                mat_A[113][3] * mat_B[62][3] +
                mat_A[114][0] * mat_B[70][3] +
                mat_A[114][1] * mat_B[78][3] +
                mat_A[114][2] * mat_B[86][3] +
                mat_A[114][3] * mat_B[94][3] +
                mat_A[115][0] * mat_B[102][3] +
                mat_A[115][1] * mat_B[110][3] +
                mat_A[115][2] * mat_B[118][3] +
                mat_A[115][3] * mat_B[126][3] +
                mat_A[116][0] * mat_B[134][3] +
                mat_A[116][1] * mat_B[142][3] +
                mat_A[116][2] * mat_B[150][3] +
                mat_A[116][3] * mat_B[158][3] +
                mat_A[117][0] * mat_B[166][3] +
                mat_A[117][1] * mat_B[174][3] +
                mat_A[117][2] * mat_B[182][3] +
                mat_A[117][3] * mat_B[190][3] +
                mat_A[118][0] * mat_B[198][3] +
                mat_A[118][1] * mat_B[206][3] +
                mat_A[118][2] * mat_B[214][3] +
                mat_A[118][3] * mat_B[222][3] +
                mat_A[119][0] * mat_B[230][3] +
                mat_A[119][1] * mat_B[238][3] +
                mat_A[119][2] * mat_B[246][3] +
                mat_A[119][3] * mat_B[254][3];
    mat_C[119][0] <=
                mat_A[112][0] * mat_B[7][0] +
                mat_A[112][1] * mat_B[15][0] +
                mat_A[112][2] * mat_B[23][0] +
                mat_A[112][3] * mat_B[31][0] +
                mat_A[113][0] * mat_B[39][0] +
                mat_A[113][1] * mat_B[47][0] +
                mat_A[113][2] * mat_B[55][0] +
                mat_A[113][3] * mat_B[63][0] +
                mat_A[114][0] * mat_B[71][0] +
                mat_A[114][1] * mat_B[79][0] +
                mat_A[114][2] * mat_B[87][0] +
                mat_A[114][3] * mat_B[95][0] +
                mat_A[115][0] * mat_B[103][0] +
                mat_A[115][1] * mat_B[111][0] +
                mat_A[115][2] * mat_B[119][0] +
                mat_A[115][3] * mat_B[127][0] +
                mat_A[116][0] * mat_B[135][0] +
                mat_A[116][1] * mat_B[143][0] +
                mat_A[116][2] * mat_B[151][0] +
                mat_A[116][3] * mat_B[159][0] +
                mat_A[117][0] * mat_B[167][0] +
                mat_A[117][1] * mat_B[175][0] +
                mat_A[117][2] * mat_B[183][0] +
                mat_A[117][3] * mat_B[191][0] +
                mat_A[118][0] * mat_B[199][0] +
                mat_A[118][1] * mat_B[207][0] +
                mat_A[118][2] * mat_B[215][0] +
                mat_A[118][3] * mat_B[223][0] +
                mat_A[119][0] * mat_B[231][0] +
                mat_A[119][1] * mat_B[239][0] +
                mat_A[119][2] * mat_B[247][0] +
                mat_A[119][3] * mat_B[255][0];
    mat_C[119][1] <=
                mat_A[112][0] * mat_B[7][1] +
                mat_A[112][1] * mat_B[15][1] +
                mat_A[112][2] * mat_B[23][1] +
                mat_A[112][3] * mat_B[31][1] +
                mat_A[113][0] * mat_B[39][1] +
                mat_A[113][1] * mat_B[47][1] +
                mat_A[113][2] * mat_B[55][1] +
                mat_A[113][3] * mat_B[63][1] +
                mat_A[114][0] * mat_B[71][1] +
                mat_A[114][1] * mat_B[79][1] +
                mat_A[114][2] * mat_B[87][1] +
                mat_A[114][3] * mat_B[95][1] +
                mat_A[115][0] * mat_B[103][1] +
                mat_A[115][1] * mat_B[111][1] +
                mat_A[115][2] * mat_B[119][1] +
                mat_A[115][3] * mat_B[127][1] +
                mat_A[116][0] * mat_B[135][1] +
                mat_A[116][1] * mat_B[143][1] +
                mat_A[116][2] * mat_B[151][1] +
                mat_A[116][3] * mat_B[159][1] +
                mat_A[117][0] * mat_B[167][1] +
                mat_A[117][1] * mat_B[175][1] +
                mat_A[117][2] * mat_B[183][1] +
                mat_A[117][3] * mat_B[191][1] +
                mat_A[118][0] * mat_B[199][1] +
                mat_A[118][1] * mat_B[207][1] +
                mat_A[118][2] * mat_B[215][1] +
                mat_A[118][3] * mat_B[223][1] +
                mat_A[119][0] * mat_B[231][1] +
                mat_A[119][1] * mat_B[239][1] +
                mat_A[119][2] * mat_B[247][1] +
                mat_A[119][3] * mat_B[255][1];
    mat_C[119][2] <=
                mat_A[112][0] * mat_B[7][2] +
                mat_A[112][1] * mat_B[15][2] +
                mat_A[112][2] * mat_B[23][2] +
                mat_A[112][3] * mat_B[31][2] +
                mat_A[113][0] * mat_B[39][2] +
                mat_A[113][1] * mat_B[47][2] +
                mat_A[113][2] * mat_B[55][2] +
                mat_A[113][3] * mat_B[63][2] +
                mat_A[114][0] * mat_B[71][2] +
                mat_A[114][1] * mat_B[79][2] +
                mat_A[114][2] * mat_B[87][2] +
                mat_A[114][3] * mat_B[95][2] +
                mat_A[115][0] * mat_B[103][2] +
                mat_A[115][1] * mat_B[111][2] +
                mat_A[115][2] * mat_B[119][2] +
                mat_A[115][3] * mat_B[127][2] +
                mat_A[116][0] * mat_B[135][2] +
                mat_A[116][1] * mat_B[143][2] +
                mat_A[116][2] * mat_B[151][2] +
                mat_A[116][3] * mat_B[159][2] +
                mat_A[117][0] * mat_B[167][2] +
                mat_A[117][1] * mat_B[175][2] +
                mat_A[117][2] * mat_B[183][2] +
                mat_A[117][3] * mat_B[191][2] +
                mat_A[118][0] * mat_B[199][2] +
                mat_A[118][1] * mat_B[207][2] +
                mat_A[118][2] * mat_B[215][2] +
                mat_A[118][3] * mat_B[223][2] +
                mat_A[119][0] * mat_B[231][2] +
                mat_A[119][1] * mat_B[239][2] +
                mat_A[119][2] * mat_B[247][2] +
                mat_A[119][3] * mat_B[255][2];
    mat_C[119][3] <=
                mat_A[112][0] * mat_B[7][3] +
                mat_A[112][1] * mat_B[15][3] +
                mat_A[112][2] * mat_B[23][3] +
                mat_A[112][3] * mat_B[31][3] +
                mat_A[113][0] * mat_B[39][3] +
                mat_A[113][1] * mat_B[47][3] +
                mat_A[113][2] * mat_B[55][3] +
                mat_A[113][3] * mat_B[63][3] +
                mat_A[114][0] * mat_B[71][3] +
                mat_A[114][1] * mat_B[79][3] +
                mat_A[114][2] * mat_B[87][3] +
                mat_A[114][3] * mat_B[95][3] +
                mat_A[115][0] * mat_B[103][3] +
                mat_A[115][1] * mat_B[111][3] +
                mat_A[115][2] * mat_B[119][3] +
                mat_A[115][3] * mat_B[127][3] +
                mat_A[116][0] * mat_B[135][3] +
                mat_A[116][1] * mat_B[143][3] +
                mat_A[116][2] * mat_B[151][3] +
                mat_A[116][3] * mat_B[159][3] +
                mat_A[117][0] * mat_B[167][3] +
                mat_A[117][1] * mat_B[175][3] +
                mat_A[117][2] * mat_B[183][3] +
                mat_A[117][3] * mat_B[191][3] +
                mat_A[118][0] * mat_B[199][3] +
                mat_A[118][1] * mat_B[207][3] +
                mat_A[118][2] * mat_B[215][3] +
                mat_A[118][3] * mat_B[223][3] +
                mat_A[119][0] * mat_B[231][3] +
                mat_A[119][1] * mat_B[239][3] +
                mat_A[119][2] * mat_B[247][3] +
                mat_A[119][3] * mat_B[255][3];
    mat_C[120][0] <=
                mat_A[120][0] * mat_B[0][0] +
                mat_A[120][1] * mat_B[8][0] +
                mat_A[120][2] * mat_B[16][0] +
                mat_A[120][3] * mat_B[24][0] +
                mat_A[121][0] * mat_B[32][0] +
                mat_A[121][1] * mat_B[40][0] +
                mat_A[121][2] * mat_B[48][0] +
                mat_A[121][3] * mat_B[56][0] +
                mat_A[122][0] * mat_B[64][0] +
                mat_A[122][1] * mat_B[72][0] +
                mat_A[122][2] * mat_B[80][0] +
                mat_A[122][3] * mat_B[88][0] +
                mat_A[123][0] * mat_B[96][0] +
                mat_A[123][1] * mat_B[104][0] +
                mat_A[123][2] * mat_B[112][0] +
                mat_A[123][3] * mat_B[120][0] +
                mat_A[124][0] * mat_B[128][0] +
                mat_A[124][1] * mat_B[136][0] +
                mat_A[124][2] * mat_B[144][0] +
                mat_A[124][3] * mat_B[152][0] +
                mat_A[125][0] * mat_B[160][0] +
                mat_A[125][1] * mat_B[168][0] +
                mat_A[125][2] * mat_B[176][0] +
                mat_A[125][3] * mat_B[184][0] +
                mat_A[126][0] * mat_B[192][0] +
                mat_A[126][1] * mat_B[200][0] +
                mat_A[126][2] * mat_B[208][0] +
                mat_A[126][3] * mat_B[216][0] +
                mat_A[127][0] * mat_B[224][0] +
                mat_A[127][1] * mat_B[232][0] +
                mat_A[127][2] * mat_B[240][0] +
                mat_A[127][3] * mat_B[248][0];
    mat_C[120][1] <=
                mat_A[120][0] * mat_B[0][1] +
                mat_A[120][1] * mat_B[8][1] +
                mat_A[120][2] * mat_B[16][1] +
                mat_A[120][3] * mat_B[24][1] +
                mat_A[121][0] * mat_B[32][1] +
                mat_A[121][1] * mat_B[40][1] +
                mat_A[121][2] * mat_B[48][1] +
                mat_A[121][3] * mat_B[56][1] +
                mat_A[122][0] * mat_B[64][1] +
                mat_A[122][1] * mat_B[72][1] +
                mat_A[122][2] * mat_B[80][1] +
                mat_A[122][3] * mat_B[88][1] +
                mat_A[123][0] * mat_B[96][1] +
                mat_A[123][1] * mat_B[104][1] +
                mat_A[123][2] * mat_B[112][1] +
                mat_A[123][3] * mat_B[120][1] +
                mat_A[124][0] * mat_B[128][1] +
                mat_A[124][1] * mat_B[136][1] +
                mat_A[124][2] * mat_B[144][1] +
                mat_A[124][3] * mat_B[152][1] +
                mat_A[125][0] * mat_B[160][1] +
                mat_A[125][1] * mat_B[168][1] +
                mat_A[125][2] * mat_B[176][1] +
                mat_A[125][3] * mat_B[184][1] +
                mat_A[126][0] * mat_B[192][1] +
                mat_A[126][1] * mat_B[200][1] +
                mat_A[126][2] * mat_B[208][1] +
                mat_A[126][3] * mat_B[216][1] +
                mat_A[127][0] * mat_B[224][1] +
                mat_A[127][1] * mat_B[232][1] +
                mat_A[127][2] * mat_B[240][1] +
                mat_A[127][3] * mat_B[248][1];
    mat_C[120][2] <=
                mat_A[120][0] * mat_B[0][2] +
                mat_A[120][1] * mat_B[8][2] +
                mat_A[120][2] * mat_B[16][2] +
                mat_A[120][3] * mat_B[24][2] +
                mat_A[121][0] * mat_B[32][2] +
                mat_A[121][1] * mat_B[40][2] +
                mat_A[121][2] * mat_B[48][2] +
                mat_A[121][3] * mat_B[56][2] +
                mat_A[122][0] * mat_B[64][2] +
                mat_A[122][1] * mat_B[72][2] +
                mat_A[122][2] * mat_B[80][2] +
                mat_A[122][3] * mat_B[88][2] +
                mat_A[123][0] * mat_B[96][2] +
                mat_A[123][1] * mat_B[104][2] +
                mat_A[123][2] * mat_B[112][2] +
                mat_A[123][3] * mat_B[120][2] +
                mat_A[124][0] * mat_B[128][2] +
                mat_A[124][1] * mat_B[136][2] +
                mat_A[124][2] * mat_B[144][2] +
                mat_A[124][3] * mat_B[152][2] +
                mat_A[125][0] * mat_B[160][2] +
                mat_A[125][1] * mat_B[168][2] +
                mat_A[125][2] * mat_B[176][2] +
                mat_A[125][3] * mat_B[184][2] +
                mat_A[126][0] * mat_B[192][2] +
                mat_A[126][1] * mat_B[200][2] +
                mat_A[126][2] * mat_B[208][2] +
                mat_A[126][3] * mat_B[216][2] +
                mat_A[127][0] * mat_B[224][2] +
                mat_A[127][1] * mat_B[232][2] +
                mat_A[127][2] * mat_B[240][2] +
                mat_A[127][3] * mat_B[248][2];
    mat_C[120][3] <=
                mat_A[120][0] * mat_B[0][3] +
                mat_A[120][1] * mat_B[8][3] +
                mat_A[120][2] * mat_B[16][3] +
                mat_A[120][3] * mat_B[24][3] +
                mat_A[121][0] * mat_B[32][3] +
                mat_A[121][1] * mat_B[40][3] +
                mat_A[121][2] * mat_B[48][3] +
                mat_A[121][3] * mat_B[56][3] +
                mat_A[122][0] * mat_B[64][3] +
                mat_A[122][1] * mat_B[72][3] +
                mat_A[122][2] * mat_B[80][3] +
                mat_A[122][3] * mat_B[88][3] +
                mat_A[123][0] * mat_B[96][3] +
                mat_A[123][1] * mat_B[104][3] +
                mat_A[123][2] * mat_B[112][3] +
                mat_A[123][3] * mat_B[120][3] +
                mat_A[124][0] * mat_B[128][3] +
                mat_A[124][1] * mat_B[136][3] +
                mat_A[124][2] * mat_B[144][3] +
                mat_A[124][3] * mat_B[152][3] +
                mat_A[125][0] * mat_B[160][3] +
                mat_A[125][1] * mat_B[168][3] +
                mat_A[125][2] * mat_B[176][3] +
                mat_A[125][3] * mat_B[184][3] +
                mat_A[126][0] * mat_B[192][3] +
                mat_A[126][1] * mat_B[200][3] +
                mat_A[126][2] * mat_B[208][3] +
                mat_A[126][3] * mat_B[216][3] +
                mat_A[127][0] * mat_B[224][3] +
                mat_A[127][1] * mat_B[232][3] +
                mat_A[127][2] * mat_B[240][3] +
                mat_A[127][3] * mat_B[248][3];
    mat_C[121][0] <=
                mat_A[120][0] * mat_B[1][0] +
                mat_A[120][1] * mat_B[9][0] +
                mat_A[120][2] * mat_B[17][0] +
                mat_A[120][3] * mat_B[25][0] +
                mat_A[121][0] * mat_B[33][0] +
                mat_A[121][1] * mat_B[41][0] +
                mat_A[121][2] * mat_B[49][0] +
                mat_A[121][3] * mat_B[57][0] +
                mat_A[122][0] * mat_B[65][0] +
                mat_A[122][1] * mat_B[73][0] +
                mat_A[122][2] * mat_B[81][0] +
                mat_A[122][3] * mat_B[89][0] +
                mat_A[123][0] * mat_B[97][0] +
                mat_A[123][1] * mat_B[105][0] +
                mat_A[123][2] * mat_B[113][0] +
                mat_A[123][3] * mat_B[121][0] +
                mat_A[124][0] * mat_B[129][0] +
                mat_A[124][1] * mat_B[137][0] +
                mat_A[124][2] * mat_B[145][0] +
                mat_A[124][3] * mat_B[153][0] +
                mat_A[125][0] * mat_B[161][0] +
                mat_A[125][1] * mat_B[169][0] +
                mat_A[125][2] * mat_B[177][0] +
                mat_A[125][3] * mat_B[185][0] +
                mat_A[126][0] * mat_B[193][0] +
                mat_A[126][1] * mat_B[201][0] +
                mat_A[126][2] * mat_B[209][0] +
                mat_A[126][3] * mat_B[217][0] +
                mat_A[127][0] * mat_B[225][0] +
                mat_A[127][1] * mat_B[233][0] +
                mat_A[127][2] * mat_B[241][0] +
                mat_A[127][3] * mat_B[249][0];
    mat_C[121][1] <=
                mat_A[120][0] * mat_B[1][1] +
                mat_A[120][1] * mat_B[9][1] +
                mat_A[120][2] * mat_B[17][1] +
                mat_A[120][3] * mat_B[25][1] +
                mat_A[121][0] * mat_B[33][1] +
                mat_A[121][1] * mat_B[41][1] +
                mat_A[121][2] * mat_B[49][1] +
                mat_A[121][3] * mat_B[57][1] +
                mat_A[122][0] * mat_B[65][1] +
                mat_A[122][1] * mat_B[73][1] +
                mat_A[122][2] * mat_B[81][1] +
                mat_A[122][3] * mat_B[89][1] +
                mat_A[123][0] * mat_B[97][1] +
                mat_A[123][1] * mat_B[105][1] +
                mat_A[123][2] * mat_B[113][1] +
                mat_A[123][3] * mat_B[121][1] +
                mat_A[124][0] * mat_B[129][1] +
                mat_A[124][1] * mat_B[137][1] +
                mat_A[124][2] * mat_B[145][1] +
                mat_A[124][3] * mat_B[153][1] +
                mat_A[125][0] * mat_B[161][1] +
                mat_A[125][1] * mat_B[169][1] +
                mat_A[125][2] * mat_B[177][1] +
                mat_A[125][3] * mat_B[185][1] +
                mat_A[126][0] * mat_B[193][1] +
                mat_A[126][1] * mat_B[201][1] +
                mat_A[126][2] * mat_B[209][1] +
                mat_A[126][3] * mat_B[217][1] +
                mat_A[127][0] * mat_B[225][1] +
                mat_A[127][1] * mat_B[233][1] +
                mat_A[127][2] * mat_B[241][1] +
                mat_A[127][3] * mat_B[249][1];
    mat_C[121][2] <=
                mat_A[120][0] * mat_B[1][2] +
                mat_A[120][1] * mat_B[9][2] +
                mat_A[120][2] * mat_B[17][2] +
                mat_A[120][3] * mat_B[25][2] +
                mat_A[121][0] * mat_B[33][2] +
                mat_A[121][1] * mat_B[41][2] +
                mat_A[121][2] * mat_B[49][2] +
                mat_A[121][3] * mat_B[57][2] +
                mat_A[122][0] * mat_B[65][2] +
                mat_A[122][1] * mat_B[73][2] +
                mat_A[122][2] * mat_B[81][2] +
                mat_A[122][3] * mat_B[89][2] +
                mat_A[123][0] * mat_B[97][2] +
                mat_A[123][1] * mat_B[105][2] +
                mat_A[123][2] * mat_B[113][2] +
                mat_A[123][3] * mat_B[121][2] +
                mat_A[124][0] * mat_B[129][2] +
                mat_A[124][1] * mat_B[137][2] +
                mat_A[124][2] * mat_B[145][2] +
                mat_A[124][3] * mat_B[153][2] +
                mat_A[125][0] * mat_B[161][2] +
                mat_A[125][1] * mat_B[169][2] +
                mat_A[125][2] * mat_B[177][2] +
                mat_A[125][3] * mat_B[185][2] +
                mat_A[126][0] * mat_B[193][2] +
                mat_A[126][1] * mat_B[201][2] +
                mat_A[126][2] * mat_B[209][2] +
                mat_A[126][3] * mat_B[217][2] +
                mat_A[127][0] * mat_B[225][2] +
                mat_A[127][1] * mat_B[233][2] +
                mat_A[127][2] * mat_B[241][2] +
                mat_A[127][3] * mat_B[249][2];
    mat_C[121][3] <=
                mat_A[120][0] * mat_B[1][3] +
                mat_A[120][1] * mat_B[9][3] +
                mat_A[120][2] * mat_B[17][3] +
                mat_A[120][3] * mat_B[25][3] +
                mat_A[121][0] * mat_B[33][3] +
                mat_A[121][1] * mat_B[41][3] +
                mat_A[121][2] * mat_B[49][3] +
                mat_A[121][3] * mat_B[57][3] +
                mat_A[122][0] * mat_B[65][3] +
                mat_A[122][1] * mat_B[73][3] +
                mat_A[122][2] * mat_B[81][3] +
                mat_A[122][3] * mat_B[89][3] +
                mat_A[123][0] * mat_B[97][3] +
                mat_A[123][1] * mat_B[105][3] +
                mat_A[123][2] * mat_B[113][3] +
                mat_A[123][3] * mat_B[121][3] +
                mat_A[124][0] * mat_B[129][3] +
                mat_A[124][1] * mat_B[137][3] +
                mat_A[124][2] * mat_B[145][3] +
                mat_A[124][3] * mat_B[153][3] +
                mat_A[125][0] * mat_B[161][3] +
                mat_A[125][1] * mat_B[169][3] +
                mat_A[125][2] * mat_B[177][3] +
                mat_A[125][3] * mat_B[185][3] +
                mat_A[126][0] * mat_B[193][3] +
                mat_A[126][1] * mat_B[201][3] +
                mat_A[126][2] * mat_B[209][3] +
                mat_A[126][3] * mat_B[217][3] +
                mat_A[127][0] * mat_B[225][3] +
                mat_A[127][1] * mat_B[233][3] +
                mat_A[127][2] * mat_B[241][3] +
                mat_A[127][3] * mat_B[249][3];
    mat_C[122][0] <=
                mat_A[120][0] * mat_B[2][0] +
                mat_A[120][1] * mat_B[10][0] +
                mat_A[120][2] * mat_B[18][0] +
                mat_A[120][3] * mat_B[26][0] +
                mat_A[121][0] * mat_B[34][0] +
                mat_A[121][1] * mat_B[42][0] +
                mat_A[121][2] * mat_B[50][0] +
                mat_A[121][3] * mat_B[58][0] +
                mat_A[122][0] * mat_B[66][0] +
                mat_A[122][1] * mat_B[74][0] +
                mat_A[122][2] * mat_B[82][0] +
                mat_A[122][3] * mat_B[90][0] +
                mat_A[123][0] * mat_B[98][0] +
                mat_A[123][1] * mat_B[106][0] +
                mat_A[123][2] * mat_B[114][0] +
                mat_A[123][3] * mat_B[122][0] +
                mat_A[124][0] * mat_B[130][0] +
                mat_A[124][1] * mat_B[138][0] +
                mat_A[124][2] * mat_B[146][0] +
                mat_A[124][3] * mat_B[154][0] +
                mat_A[125][0] * mat_B[162][0] +
                mat_A[125][1] * mat_B[170][0] +
                mat_A[125][2] * mat_B[178][0] +
                mat_A[125][3] * mat_B[186][0] +
                mat_A[126][0] * mat_B[194][0] +
                mat_A[126][1] * mat_B[202][0] +
                mat_A[126][2] * mat_B[210][0] +
                mat_A[126][3] * mat_B[218][0] +
                mat_A[127][0] * mat_B[226][0] +
                mat_A[127][1] * mat_B[234][0] +
                mat_A[127][2] * mat_B[242][0] +
                mat_A[127][3] * mat_B[250][0];
    mat_C[122][1] <=
                mat_A[120][0] * mat_B[2][1] +
                mat_A[120][1] * mat_B[10][1] +
                mat_A[120][2] * mat_B[18][1] +
                mat_A[120][3] * mat_B[26][1] +
                mat_A[121][0] * mat_B[34][1] +
                mat_A[121][1] * mat_B[42][1] +
                mat_A[121][2] * mat_B[50][1] +
                mat_A[121][3] * mat_B[58][1] +
                mat_A[122][0] * mat_B[66][1] +
                mat_A[122][1] * mat_B[74][1] +
                mat_A[122][2] * mat_B[82][1] +
                mat_A[122][3] * mat_B[90][1] +
                mat_A[123][0] * mat_B[98][1] +
                mat_A[123][1] * mat_B[106][1] +
                mat_A[123][2] * mat_B[114][1] +
                mat_A[123][3] * mat_B[122][1] +
                mat_A[124][0] * mat_B[130][1] +
                mat_A[124][1] * mat_B[138][1] +
                mat_A[124][2] * mat_B[146][1] +
                mat_A[124][3] * mat_B[154][1] +
                mat_A[125][0] * mat_B[162][1] +
                mat_A[125][1] * mat_B[170][1] +
                mat_A[125][2] * mat_B[178][1] +
                mat_A[125][3] * mat_B[186][1] +
                mat_A[126][0] * mat_B[194][1] +
                mat_A[126][1] * mat_B[202][1] +
                mat_A[126][2] * mat_B[210][1] +
                mat_A[126][3] * mat_B[218][1] +
                mat_A[127][0] * mat_B[226][1] +
                mat_A[127][1] * mat_B[234][1] +
                mat_A[127][2] * mat_B[242][1] +
                mat_A[127][3] * mat_B[250][1];
    mat_C[122][2] <=
                mat_A[120][0] * mat_B[2][2] +
                mat_A[120][1] * mat_B[10][2] +
                mat_A[120][2] * mat_B[18][2] +
                mat_A[120][3] * mat_B[26][2] +
                mat_A[121][0] * mat_B[34][2] +
                mat_A[121][1] * mat_B[42][2] +
                mat_A[121][2] * mat_B[50][2] +
                mat_A[121][3] * mat_B[58][2] +
                mat_A[122][0] * mat_B[66][2] +
                mat_A[122][1] * mat_B[74][2] +
                mat_A[122][2] * mat_B[82][2] +
                mat_A[122][3] * mat_B[90][2] +
                mat_A[123][0] * mat_B[98][2] +
                mat_A[123][1] * mat_B[106][2] +
                mat_A[123][2] * mat_B[114][2] +
                mat_A[123][3] * mat_B[122][2] +
                mat_A[124][0] * mat_B[130][2] +
                mat_A[124][1] * mat_B[138][2] +
                mat_A[124][2] * mat_B[146][2] +
                mat_A[124][3] * mat_B[154][2] +
                mat_A[125][0] * mat_B[162][2] +
                mat_A[125][1] * mat_B[170][2] +
                mat_A[125][2] * mat_B[178][2] +
                mat_A[125][3] * mat_B[186][2] +
                mat_A[126][0] * mat_B[194][2] +
                mat_A[126][1] * mat_B[202][2] +
                mat_A[126][2] * mat_B[210][2] +
                mat_A[126][3] * mat_B[218][2] +
                mat_A[127][0] * mat_B[226][2] +
                mat_A[127][1] * mat_B[234][2] +
                mat_A[127][2] * mat_B[242][2] +
                mat_A[127][3] * mat_B[250][2];
    mat_C[122][3] <=
                mat_A[120][0] * mat_B[2][3] +
                mat_A[120][1] * mat_B[10][3] +
                mat_A[120][2] * mat_B[18][3] +
                mat_A[120][3] * mat_B[26][3] +
                mat_A[121][0] * mat_B[34][3] +
                mat_A[121][1] * mat_B[42][3] +
                mat_A[121][2] * mat_B[50][3] +
                mat_A[121][3] * mat_B[58][3] +
                mat_A[122][0] * mat_B[66][3] +
                mat_A[122][1] * mat_B[74][3] +
                mat_A[122][2] * mat_B[82][3] +
                mat_A[122][3] * mat_B[90][3] +
                mat_A[123][0] * mat_B[98][3] +
                mat_A[123][1] * mat_B[106][3] +
                mat_A[123][2] * mat_B[114][3] +
                mat_A[123][3] * mat_B[122][3] +
                mat_A[124][0] * mat_B[130][3] +
                mat_A[124][1] * mat_B[138][3] +
                mat_A[124][2] * mat_B[146][3] +
                mat_A[124][3] * mat_B[154][3] +
                mat_A[125][0] * mat_B[162][3] +
                mat_A[125][1] * mat_B[170][3] +
                mat_A[125][2] * mat_B[178][3] +
                mat_A[125][3] * mat_B[186][3] +
                mat_A[126][0] * mat_B[194][3] +
                mat_A[126][1] * mat_B[202][3] +
                mat_A[126][2] * mat_B[210][3] +
                mat_A[126][3] * mat_B[218][3] +
                mat_A[127][0] * mat_B[226][3] +
                mat_A[127][1] * mat_B[234][3] +
                mat_A[127][2] * mat_B[242][3] +
                mat_A[127][3] * mat_B[250][3];
    mat_C[123][0] <=
                mat_A[120][0] * mat_B[3][0] +
                mat_A[120][1] * mat_B[11][0] +
                mat_A[120][2] * mat_B[19][0] +
                mat_A[120][3] * mat_B[27][0] +
                mat_A[121][0] * mat_B[35][0] +
                mat_A[121][1] * mat_B[43][0] +
                mat_A[121][2] * mat_B[51][0] +
                mat_A[121][3] * mat_B[59][0] +
                mat_A[122][0] * mat_B[67][0] +
                mat_A[122][1] * mat_B[75][0] +
                mat_A[122][2] * mat_B[83][0] +
                mat_A[122][3] * mat_B[91][0] +
                mat_A[123][0] * mat_B[99][0] +
                mat_A[123][1] * mat_B[107][0] +
                mat_A[123][2] * mat_B[115][0] +
                mat_A[123][3] * mat_B[123][0] +
                mat_A[124][0] * mat_B[131][0] +
                mat_A[124][1] * mat_B[139][0] +
                mat_A[124][2] * mat_B[147][0] +
                mat_A[124][3] * mat_B[155][0] +
                mat_A[125][0] * mat_B[163][0] +
                mat_A[125][1] * mat_B[171][0] +
                mat_A[125][2] * mat_B[179][0] +
                mat_A[125][3] * mat_B[187][0] +
                mat_A[126][0] * mat_B[195][0] +
                mat_A[126][1] * mat_B[203][0] +
                mat_A[126][2] * mat_B[211][0] +
                mat_A[126][3] * mat_B[219][0] +
                mat_A[127][0] * mat_B[227][0] +
                mat_A[127][1] * mat_B[235][0] +
                mat_A[127][2] * mat_B[243][0] +
                mat_A[127][3] * mat_B[251][0];
    mat_C[123][1] <=
                mat_A[120][0] * mat_B[3][1] +
                mat_A[120][1] * mat_B[11][1] +
                mat_A[120][2] * mat_B[19][1] +
                mat_A[120][3] * mat_B[27][1] +
                mat_A[121][0] * mat_B[35][1] +
                mat_A[121][1] * mat_B[43][1] +
                mat_A[121][2] * mat_B[51][1] +
                mat_A[121][3] * mat_B[59][1] +
                mat_A[122][0] * mat_B[67][1] +
                mat_A[122][1] * mat_B[75][1] +
                mat_A[122][2] * mat_B[83][1] +
                mat_A[122][3] * mat_B[91][1] +
                mat_A[123][0] * mat_B[99][1] +
                mat_A[123][1] * mat_B[107][1] +
                mat_A[123][2] * mat_B[115][1] +
                mat_A[123][3] * mat_B[123][1] +
                mat_A[124][0] * mat_B[131][1] +
                mat_A[124][1] * mat_B[139][1] +
                mat_A[124][2] * mat_B[147][1] +
                mat_A[124][3] * mat_B[155][1] +
                mat_A[125][0] * mat_B[163][1] +
                mat_A[125][1] * mat_B[171][1] +
                mat_A[125][2] * mat_B[179][1] +
                mat_A[125][3] * mat_B[187][1] +
                mat_A[126][0] * mat_B[195][1] +
                mat_A[126][1] * mat_B[203][1] +
                mat_A[126][2] * mat_B[211][1] +
                mat_A[126][3] * mat_B[219][1] +
                mat_A[127][0] * mat_B[227][1] +
                mat_A[127][1] * mat_B[235][1] +
                mat_A[127][2] * mat_B[243][1] +
                mat_A[127][3] * mat_B[251][1];
    mat_C[123][2] <=
                mat_A[120][0] * mat_B[3][2] +
                mat_A[120][1] * mat_B[11][2] +
                mat_A[120][2] * mat_B[19][2] +
                mat_A[120][3] * mat_B[27][2] +
                mat_A[121][0] * mat_B[35][2] +
                mat_A[121][1] * mat_B[43][2] +
                mat_A[121][2] * mat_B[51][2] +
                mat_A[121][3] * mat_B[59][2] +
                mat_A[122][0] * mat_B[67][2] +
                mat_A[122][1] * mat_B[75][2] +
                mat_A[122][2] * mat_B[83][2] +
                mat_A[122][3] * mat_B[91][2] +
                mat_A[123][0] * mat_B[99][2] +
                mat_A[123][1] * mat_B[107][2] +
                mat_A[123][2] * mat_B[115][2] +
                mat_A[123][3] * mat_B[123][2] +
                mat_A[124][0] * mat_B[131][2] +
                mat_A[124][1] * mat_B[139][2] +
                mat_A[124][2] * mat_B[147][2] +
                mat_A[124][3] * mat_B[155][2] +
                mat_A[125][0] * mat_B[163][2] +
                mat_A[125][1] * mat_B[171][2] +
                mat_A[125][2] * mat_B[179][2] +
                mat_A[125][3] * mat_B[187][2] +
                mat_A[126][0] * mat_B[195][2] +
                mat_A[126][1] * mat_B[203][2] +
                mat_A[126][2] * mat_B[211][2] +
                mat_A[126][3] * mat_B[219][2] +
                mat_A[127][0] * mat_B[227][2] +
                mat_A[127][1] * mat_B[235][2] +
                mat_A[127][2] * mat_B[243][2] +
                mat_A[127][3] * mat_B[251][2];
    mat_C[123][3] <=
                mat_A[120][0] * mat_B[3][3] +
                mat_A[120][1] * mat_B[11][3] +
                mat_A[120][2] * mat_B[19][3] +
                mat_A[120][3] * mat_B[27][3] +
                mat_A[121][0] * mat_B[35][3] +
                mat_A[121][1] * mat_B[43][3] +
                mat_A[121][2] * mat_B[51][3] +
                mat_A[121][3] * mat_B[59][3] +
                mat_A[122][0] * mat_B[67][3] +
                mat_A[122][1] * mat_B[75][3] +
                mat_A[122][2] * mat_B[83][3] +
                mat_A[122][3] * mat_B[91][3] +
                mat_A[123][0] * mat_B[99][3] +
                mat_A[123][1] * mat_B[107][3] +
                mat_A[123][2] * mat_B[115][3] +
                mat_A[123][3] * mat_B[123][3] +
                mat_A[124][0] * mat_B[131][3] +
                mat_A[124][1] * mat_B[139][3] +
                mat_A[124][2] * mat_B[147][3] +
                mat_A[124][3] * mat_B[155][3] +
                mat_A[125][0] * mat_B[163][3] +
                mat_A[125][1] * mat_B[171][3] +
                mat_A[125][2] * mat_B[179][3] +
                mat_A[125][3] * mat_B[187][3] +
                mat_A[126][0] * mat_B[195][3] +
                mat_A[126][1] * mat_B[203][3] +
                mat_A[126][2] * mat_B[211][3] +
                mat_A[126][3] * mat_B[219][3] +
                mat_A[127][0] * mat_B[227][3] +
                mat_A[127][1] * mat_B[235][3] +
                mat_A[127][2] * mat_B[243][3] +
                mat_A[127][3] * mat_B[251][3];
    mat_C[124][0] <=
                mat_A[120][0] * mat_B[4][0] +
                mat_A[120][1] * mat_B[12][0] +
                mat_A[120][2] * mat_B[20][0] +
                mat_A[120][3] * mat_B[28][0] +
                mat_A[121][0] * mat_B[36][0] +
                mat_A[121][1] * mat_B[44][0] +
                mat_A[121][2] * mat_B[52][0] +
                mat_A[121][3] * mat_B[60][0] +
                mat_A[122][0] * mat_B[68][0] +
                mat_A[122][1] * mat_B[76][0] +
                mat_A[122][2] * mat_B[84][0] +
                mat_A[122][3] * mat_B[92][0] +
                mat_A[123][0] * mat_B[100][0] +
                mat_A[123][1] * mat_B[108][0] +
                mat_A[123][2] * mat_B[116][0] +
                mat_A[123][3] * mat_B[124][0] +
                mat_A[124][0] * mat_B[132][0] +
                mat_A[124][1] * mat_B[140][0] +
                mat_A[124][2] * mat_B[148][0] +
                mat_A[124][3] * mat_B[156][0] +
                mat_A[125][0] * mat_B[164][0] +
                mat_A[125][1] * mat_B[172][0] +
                mat_A[125][2] * mat_B[180][0] +
                mat_A[125][3] * mat_B[188][0] +
                mat_A[126][0] * mat_B[196][0] +
                mat_A[126][1] * mat_B[204][0] +
                mat_A[126][2] * mat_B[212][0] +
                mat_A[126][3] * mat_B[220][0] +
                mat_A[127][0] * mat_B[228][0] +
                mat_A[127][1] * mat_B[236][0] +
                mat_A[127][2] * mat_B[244][0] +
                mat_A[127][3] * mat_B[252][0];
    mat_C[124][1] <=
                mat_A[120][0] * mat_B[4][1] +
                mat_A[120][1] * mat_B[12][1] +
                mat_A[120][2] * mat_B[20][1] +
                mat_A[120][3] * mat_B[28][1] +
                mat_A[121][0] * mat_B[36][1] +
                mat_A[121][1] * mat_B[44][1] +
                mat_A[121][2] * mat_B[52][1] +
                mat_A[121][3] * mat_B[60][1] +
                mat_A[122][0] * mat_B[68][1] +
                mat_A[122][1] * mat_B[76][1] +
                mat_A[122][2] * mat_B[84][1] +
                mat_A[122][3] * mat_B[92][1] +
                mat_A[123][0] * mat_B[100][1] +
                mat_A[123][1] * mat_B[108][1] +
                mat_A[123][2] * mat_B[116][1] +
                mat_A[123][3] * mat_B[124][1] +
                mat_A[124][0] * mat_B[132][1] +
                mat_A[124][1] * mat_B[140][1] +
                mat_A[124][2] * mat_B[148][1] +
                mat_A[124][3] * mat_B[156][1] +
                mat_A[125][0] * mat_B[164][1] +
                mat_A[125][1] * mat_B[172][1] +
                mat_A[125][2] * mat_B[180][1] +
                mat_A[125][3] * mat_B[188][1] +
                mat_A[126][0] * mat_B[196][1] +
                mat_A[126][1] * mat_B[204][1] +
                mat_A[126][2] * mat_B[212][1] +
                mat_A[126][3] * mat_B[220][1] +
                mat_A[127][0] * mat_B[228][1] +
                mat_A[127][1] * mat_B[236][1] +
                mat_A[127][2] * mat_B[244][1] +
                mat_A[127][3] * mat_B[252][1];
    mat_C[124][2] <=
                mat_A[120][0] * mat_B[4][2] +
                mat_A[120][1] * mat_B[12][2] +
                mat_A[120][2] * mat_B[20][2] +
                mat_A[120][3] * mat_B[28][2] +
                mat_A[121][0] * mat_B[36][2] +
                mat_A[121][1] * mat_B[44][2] +
                mat_A[121][2] * mat_B[52][2] +
                mat_A[121][3] * mat_B[60][2] +
                mat_A[122][0] * mat_B[68][2] +
                mat_A[122][1] * mat_B[76][2] +
                mat_A[122][2] * mat_B[84][2] +
                mat_A[122][3] * mat_B[92][2] +
                mat_A[123][0] * mat_B[100][2] +
                mat_A[123][1] * mat_B[108][2] +
                mat_A[123][2] * mat_B[116][2] +
                mat_A[123][3] * mat_B[124][2] +
                mat_A[124][0] * mat_B[132][2] +
                mat_A[124][1] * mat_B[140][2] +
                mat_A[124][2] * mat_B[148][2] +
                mat_A[124][3] * mat_B[156][2] +
                mat_A[125][0] * mat_B[164][2] +
                mat_A[125][1] * mat_B[172][2] +
                mat_A[125][2] * mat_B[180][2] +
                mat_A[125][3] * mat_B[188][2] +
                mat_A[126][0] * mat_B[196][2] +
                mat_A[126][1] * mat_B[204][2] +
                mat_A[126][2] * mat_B[212][2] +
                mat_A[126][3] * mat_B[220][2] +
                mat_A[127][0] * mat_B[228][2] +
                mat_A[127][1] * mat_B[236][2] +
                mat_A[127][2] * mat_B[244][2] +
                mat_A[127][3] * mat_B[252][2];
    mat_C[124][3] <=
                mat_A[120][0] * mat_B[4][3] +
                mat_A[120][1] * mat_B[12][3] +
                mat_A[120][2] * mat_B[20][3] +
                mat_A[120][3] * mat_B[28][3] +
                mat_A[121][0] * mat_B[36][3] +
                mat_A[121][1] * mat_B[44][3] +
                mat_A[121][2] * mat_B[52][3] +
                mat_A[121][3] * mat_B[60][3] +
                mat_A[122][0] * mat_B[68][3] +
                mat_A[122][1] * mat_B[76][3] +
                mat_A[122][2] * mat_B[84][3] +
                mat_A[122][3] * mat_B[92][3] +
                mat_A[123][0] * mat_B[100][3] +
                mat_A[123][1] * mat_B[108][3] +
                mat_A[123][2] * mat_B[116][3] +
                mat_A[123][3] * mat_B[124][3] +
                mat_A[124][0] * mat_B[132][3] +
                mat_A[124][1] * mat_B[140][3] +
                mat_A[124][2] * mat_B[148][3] +
                mat_A[124][3] * mat_B[156][3] +
                mat_A[125][0] * mat_B[164][3] +
                mat_A[125][1] * mat_B[172][3] +
                mat_A[125][2] * mat_B[180][3] +
                mat_A[125][3] * mat_B[188][3] +
                mat_A[126][0] * mat_B[196][3] +
                mat_A[126][1] * mat_B[204][3] +
                mat_A[126][2] * mat_B[212][3] +
                mat_A[126][3] * mat_B[220][3] +
                mat_A[127][0] * mat_B[228][3] +
                mat_A[127][1] * mat_B[236][3] +
                mat_A[127][2] * mat_B[244][3] +
                mat_A[127][3] * mat_B[252][3];
    mat_C[125][0] <=
                mat_A[120][0] * mat_B[5][0] +
                mat_A[120][1] * mat_B[13][0] +
                mat_A[120][2] * mat_B[21][0] +
                mat_A[120][3] * mat_B[29][0] +
                mat_A[121][0] * mat_B[37][0] +
                mat_A[121][1] * mat_B[45][0] +
                mat_A[121][2] * mat_B[53][0] +
                mat_A[121][3] * mat_B[61][0] +
                mat_A[122][0] * mat_B[69][0] +
                mat_A[122][1] * mat_B[77][0] +
                mat_A[122][2] * mat_B[85][0] +
                mat_A[122][3] * mat_B[93][0] +
                mat_A[123][0] * mat_B[101][0] +
                mat_A[123][1] * mat_B[109][0] +
                mat_A[123][2] * mat_B[117][0] +
                mat_A[123][3] * mat_B[125][0] +
                mat_A[124][0] * mat_B[133][0] +
                mat_A[124][1] * mat_B[141][0] +
                mat_A[124][2] * mat_B[149][0] +
                mat_A[124][3] * mat_B[157][0] +
                mat_A[125][0] * mat_B[165][0] +
                mat_A[125][1] * mat_B[173][0] +
                mat_A[125][2] * mat_B[181][0] +
                mat_A[125][3] * mat_B[189][0] +
                mat_A[126][0] * mat_B[197][0] +
                mat_A[126][1] * mat_B[205][0] +
                mat_A[126][2] * mat_B[213][0] +
                mat_A[126][3] * mat_B[221][0] +
                mat_A[127][0] * mat_B[229][0] +
                mat_A[127][1] * mat_B[237][0] +
                mat_A[127][2] * mat_B[245][0] +
                mat_A[127][3] * mat_B[253][0];
    mat_C[125][1] <=
                mat_A[120][0] * mat_B[5][1] +
                mat_A[120][1] * mat_B[13][1] +
                mat_A[120][2] * mat_B[21][1] +
                mat_A[120][3] * mat_B[29][1] +
                mat_A[121][0] * mat_B[37][1] +
                mat_A[121][1] * mat_B[45][1] +
                mat_A[121][2] * mat_B[53][1] +
                mat_A[121][3] * mat_B[61][1] +
                mat_A[122][0] * mat_B[69][1] +
                mat_A[122][1] * mat_B[77][1] +
                mat_A[122][2] * mat_B[85][1] +
                mat_A[122][3] * mat_B[93][1] +
                mat_A[123][0] * mat_B[101][1] +
                mat_A[123][1] * mat_B[109][1] +
                mat_A[123][2] * mat_B[117][1] +
                mat_A[123][3] * mat_B[125][1] +
                mat_A[124][0] * mat_B[133][1] +
                mat_A[124][1] * mat_B[141][1] +
                mat_A[124][2] * mat_B[149][1] +
                mat_A[124][3] * mat_B[157][1] +
                mat_A[125][0] * mat_B[165][1] +
                mat_A[125][1] * mat_B[173][1] +
                mat_A[125][2] * mat_B[181][1] +
                mat_A[125][3] * mat_B[189][1] +
                mat_A[126][0] * mat_B[197][1] +
                mat_A[126][1] * mat_B[205][1] +
                mat_A[126][2] * mat_B[213][1] +
                mat_A[126][3] * mat_B[221][1] +
                mat_A[127][0] * mat_B[229][1] +
                mat_A[127][1] * mat_B[237][1] +
                mat_A[127][2] * mat_B[245][1] +
                mat_A[127][3] * mat_B[253][1];
    mat_C[125][2] <=
                mat_A[120][0] * mat_B[5][2] +
                mat_A[120][1] * mat_B[13][2] +
                mat_A[120][2] * mat_B[21][2] +
                mat_A[120][3] * mat_B[29][2] +
                mat_A[121][0] * mat_B[37][2] +
                mat_A[121][1] * mat_B[45][2] +
                mat_A[121][2] * mat_B[53][2] +
                mat_A[121][3] * mat_B[61][2] +
                mat_A[122][0] * mat_B[69][2] +
                mat_A[122][1] * mat_B[77][2] +
                mat_A[122][2] * mat_B[85][2] +
                mat_A[122][3] * mat_B[93][2] +
                mat_A[123][0] * mat_B[101][2] +
                mat_A[123][1] * mat_B[109][2] +
                mat_A[123][2] * mat_B[117][2] +
                mat_A[123][3] * mat_B[125][2] +
                mat_A[124][0] * mat_B[133][2] +
                mat_A[124][1] * mat_B[141][2] +
                mat_A[124][2] * mat_B[149][2] +
                mat_A[124][3] * mat_B[157][2] +
                mat_A[125][0] * mat_B[165][2] +
                mat_A[125][1] * mat_B[173][2] +
                mat_A[125][2] * mat_B[181][2] +
                mat_A[125][3] * mat_B[189][2] +
                mat_A[126][0] * mat_B[197][2] +
                mat_A[126][1] * mat_B[205][2] +
                mat_A[126][2] * mat_B[213][2] +
                mat_A[126][3] * mat_B[221][2] +
                mat_A[127][0] * mat_B[229][2] +
                mat_A[127][1] * mat_B[237][2] +
                mat_A[127][2] * mat_B[245][2] +
                mat_A[127][3] * mat_B[253][2];
    mat_C[125][3] <=
                mat_A[120][0] * mat_B[5][3] +
                mat_A[120][1] * mat_B[13][3] +
                mat_A[120][2] * mat_B[21][3] +
                mat_A[120][3] * mat_B[29][3] +
                mat_A[121][0] * mat_B[37][3] +
                mat_A[121][1] * mat_B[45][3] +
                mat_A[121][2] * mat_B[53][3] +
                mat_A[121][3] * mat_B[61][3] +
                mat_A[122][0] * mat_B[69][3] +
                mat_A[122][1] * mat_B[77][3] +
                mat_A[122][2] * mat_B[85][3] +
                mat_A[122][3] * mat_B[93][3] +
                mat_A[123][0] * mat_B[101][3] +
                mat_A[123][1] * mat_B[109][3] +
                mat_A[123][2] * mat_B[117][3] +
                mat_A[123][3] * mat_B[125][3] +
                mat_A[124][0] * mat_B[133][3] +
                mat_A[124][1] * mat_B[141][3] +
                mat_A[124][2] * mat_B[149][3] +
                mat_A[124][3] * mat_B[157][3] +
                mat_A[125][0] * mat_B[165][3] +
                mat_A[125][1] * mat_B[173][3] +
                mat_A[125][2] * mat_B[181][3] +
                mat_A[125][3] * mat_B[189][3] +
                mat_A[126][0] * mat_B[197][3] +
                mat_A[126][1] * mat_B[205][3] +
                mat_A[126][2] * mat_B[213][3] +
                mat_A[126][3] * mat_B[221][3] +
                mat_A[127][0] * mat_B[229][3] +
                mat_A[127][1] * mat_B[237][3] +
                mat_A[127][2] * mat_B[245][3] +
                mat_A[127][3] * mat_B[253][3];
    mat_C[126][0] <=
                mat_A[120][0] * mat_B[6][0] +
                mat_A[120][1] * mat_B[14][0] +
                mat_A[120][2] * mat_B[22][0] +
                mat_A[120][3] * mat_B[30][0] +
                mat_A[121][0] * mat_B[38][0] +
                mat_A[121][1] * mat_B[46][0] +
                mat_A[121][2] * mat_B[54][0] +
                mat_A[121][3] * mat_B[62][0] +
                mat_A[122][0] * mat_B[70][0] +
                mat_A[122][1] * mat_B[78][0] +
                mat_A[122][2] * mat_B[86][0] +
                mat_A[122][3] * mat_B[94][0] +
                mat_A[123][0] * mat_B[102][0] +
                mat_A[123][1] * mat_B[110][0] +
                mat_A[123][2] * mat_B[118][0] +
                mat_A[123][3] * mat_B[126][0] +
                mat_A[124][0] * mat_B[134][0] +
                mat_A[124][1] * mat_B[142][0] +
                mat_A[124][2] * mat_B[150][0] +
                mat_A[124][3] * mat_B[158][0] +
                mat_A[125][0] * mat_B[166][0] +
                mat_A[125][1] * mat_B[174][0] +
                mat_A[125][2] * mat_B[182][0] +
                mat_A[125][3] * mat_B[190][0] +
                mat_A[126][0] * mat_B[198][0] +
                mat_A[126][1] * mat_B[206][0] +
                mat_A[126][2] * mat_B[214][0] +
                mat_A[126][3] * mat_B[222][0] +
                mat_A[127][0] * mat_B[230][0] +
                mat_A[127][1] * mat_B[238][0] +
                mat_A[127][2] * mat_B[246][0] +
                mat_A[127][3] * mat_B[254][0];
    mat_C[126][1] <=
                mat_A[120][0] * mat_B[6][1] +
                mat_A[120][1] * mat_B[14][1] +
                mat_A[120][2] * mat_B[22][1] +
                mat_A[120][3] * mat_B[30][1] +
                mat_A[121][0] * mat_B[38][1] +
                mat_A[121][1] * mat_B[46][1] +
                mat_A[121][2] * mat_B[54][1] +
                mat_A[121][3] * mat_B[62][1] +
                mat_A[122][0] * mat_B[70][1] +
                mat_A[122][1] * mat_B[78][1] +
                mat_A[122][2] * mat_B[86][1] +
                mat_A[122][3] * mat_B[94][1] +
                mat_A[123][0] * mat_B[102][1] +
                mat_A[123][1] * mat_B[110][1] +
                mat_A[123][2] * mat_B[118][1] +
                mat_A[123][3] * mat_B[126][1] +
                mat_A[124][0] * mat_B[134][1] +
                mat_A[124][1] * mat_B[142][1] +
                mat_A[124][2] * mat_B[150][1] +
                mat_A[124][3] * mat_B[158][1] +
                mat_A[125][0] * mat_B[166][1] +
                mat_A[125][1] * mat_B[174][1] +
                mat_A[125][2] * mat_B[182][1] +
                mat_A[125][3] * mat_B[190][1] +
                mat_A[126][0] * mat_B[198][1] +
                mat_A[126][1] * mat_B[206][1] +
                mat_A[126][2] * mat_B[214][1] +
                mat_A[126][3] * mat_B[222][1] +
                mat_A[127][0] * mat_B[230][1] +
                mat_A[127][1] * mat_B[238][1] +
                mat_A[127][2] * mat_B[246][1] +
                mat_A[127][3] * mat_B[254][1];
    mat_C[126][2] <=
                mat_A[120][0] * mat_B[6][2] +
                mat_A[120][1] * mat_B[14][2] +
                mat_A[120][2] * mat_B[22][2] +
                mat_A[120][3] * mat_B[30][2] +
                mat_A[121][0] * mat_B[38][2] +
                mat_A[121][1] * mat_B[46][2] +
                mat_A[121][2] * mat_B[54][2] +
                mat_A[121][3] * mat_B[62][2] +
                mat_A[122][0] * mat_B[70][2] +
                mat_A[122][1] * mat_B[78][2] +
                mat_A[122][2] * mat_B[86][2] +
                mat_A[122][3] * mat_B[94][2] +
                mat_A[123][0] * mat_B[102][2] +
                mat_A[123][1] * mat_B[110][2] +
                mat_A[123][2] * mat_B[118][2] +
                mat_A[123][3] * mat_B[126][2] +
                mat_A[124][0] * mat_B[134][2] +
                mat_A[124][1] * mat_B[142][2] +
                mat_A[124][2] * mat_B[150][2] +
                mat_A[124][3] * mat_B[158][2] +
                mat_A[125][0] * mat_B[166][2] +
                mat_A[125][1] * mat_B[174][2] +
                mat_A[125][2] * mat_B[182][2] +
                mat_A[125][3] * mat_B[190][2] +
                mat_A[126][0] * mat_B[198][2] +
                mat_A[126][1] * mat_B[206][2] +
                mat_A[126][2] * mat_B[214][2] +
                mat_A[126][3] * mat_B[222][2] +
                mat_A[127][0] * mat_B[230][2] +
                mat_A[127][1] * mat_B[238][2] +
                mat_A[127][2] * mat_B[246][2] +
                mat_A[127][3] * mat_B[254][2];
    mat_C[126][3] <=
                mat_A[120][0] * mat_B[6][3] +
                mat_A[120][1] * mat_B[14][3] +
                mat_A[120][2] * mat_B[22][3] +
                mat_A[120][3] * mat_B[30][3] +
                mat_A[121][0] * mat_B[38][3] +
                mat_A[121][1] * mat_B[46][3] +
                mat_A[121][2] * mat_B[54][3] +
                mat_A[121][3] * mat_B[62][3] +
                mat_A[122][0] * mat_B[70][3] +
                mat_A[122][1] * mat_B[78][3] +
                mat_A[122][2] * mat_B[86][3] +
                mat_A[122][3] * mat_B[94][3] +
                mat_A[123][0] * mat_B[102][3] +
                mat_A[123][1] * mat_B[110][3] +
                mat_A[123][2] * mat_B[118][3] +
                mat_A[123][3] * mat_B[126][3] +
                mat_A[124][0] * mat_B[134][3] +
                mat_A[124][1] * mat_B[142][3] +
                mat_A[124][2] * mat_B[150][3] +
                mat_A[124][3] * mat_B[158][3] +
                mat_A[125][0] * mat_B[166][3] +
                mat_A[125][1] * mat_B[174][3] +
                mat_A[125][2] * mat_B[182][3] +
                mat_A[125][3] * mat_B[190][3] +
                mat_A[126][0] * mat_B[198][3] +
                mat_A[126][1] * mat_B[206][3] +
                mat_A[126][2] * mat_B[214][3] +
                mat_A[126][3] * mat_B[222][3] +
                mat_A[127][0] * mat_B[230][3] +
                mat_A[127][1] * mat_B[238][3] +
                mat_A[127][2] * mat_B[246][3] +
                mat_A[127][3] * mat_B[254][3];
    mat_C[127][0] <=
                mat_A[120][0] * mat_B[7][0] +
                mat_A[120][1] * mat_B[15][0] +
                mat_A[120][2] * mat_B[23][0] +
                mat_A[120][3] * mat_B[31][0] +
                mat_A[121][0] * mat_B[39][0] +
                mat_A[121][1] * mat_B[47][0] +
                mat_A[121][2] * mat_B[55][0] +
                mat_A[121][3] * mat_B[63][0] +
                mat_A[122][0] * mat_B[71][0] +
                mat_A[122][1] * mat_B[79][0] +
                mat_A[122][2] * mat_B[87][0] +
                mat_A[122][3] * mat_B[95][0] +
                mat_A[123][0] * mat_B[103][0] +
                mat_A[123][1] * mat_B[111][0] +
                mat_A[123][2] * mat_B[119][0] +
                mat_A[123][3] * mat_B[127][0] +
                mat_A[124][0] * mat_B[135][0] +
                mat_A[124][1] * mat_B[143][0] +
                mat_A[124][2] * mat_B[151][0] +
                mat_A[124][3] * mat_B[159][0] +
                mat_A[125][0] * mat_B[167][0] +
                mat_A[125][1] * mat_B[175][0] +
                mat_A[125][2] * mat_B[183][0] +
                mat_A[125][3] * mat_B[191][0] +
                mat_A[126][0] * mat_B[199][0] +
                mat_A[126][1] * mat_B[207][0] +
                mat_A[126][2] * mat_B[215][0] +
                mat_A[126][3] * mat_B[223][0] +
                mat_A[127][0] * mat_B[231][0] +
                mat_A[127][1] * mat_B[239][0] +
                mat_A[127][2] * mat_B[247][0] +
                mat_A[127][3] * mat_B[255][0];
    mat_C[127][1] <=
                mat_A[120][0] * mat_B[7][1] +
                mat_A[120][1] * mat_B[15][1] +
                mat_A[120][2] * mat_B[23][1] +
                mat_A[120][3] * mat_B[31][1] +
                mat_A[121][0] * mat_B[39][1] +
                mat_A[121][1] * mat_B[47][1] +
                mat_A[121][2] * mat_B[55][1] +
                mat_A[121][3] * mat_B[63][1] +
                mat_A[122][0] * mat_B[71][1] +
                mat_A[122][1] * mat_B[79][1] +
                mat_A[122][2] * mat_B[87][1] +
                mat_A[122][3] * mat_B[95][1] +
                mat_A[123][0] * mat_B[103][1] +
                mat_A[123][1] * mat_B[111][1] +
                mat_A[123][2] * mat_B[119][1] +
                mat_A[123][3] * mat_B[127][1] +
                mat_A[124][0] * mat_B[135][1] +
                mat_A[124][1] * mat_B[143][1] +
                mat_A[124][2] * mat_B[151][1] +
                mat_A[124][3] * mat_B[159][1] +
                mat_A[125][0] * mat_B[167][1] +
                mat_A[125][1] * mat_B[175][1] +
                mat_A[125][2] * mat_B[183][1] +
                mat_A[125][3] * mat_B[191][1] +
                mat_A[126][0] * mat_B[199][1] +
                mat_A[126][1] * mat_B[207][1] +
                mat_A[126][2] * mat_B[215][1] +
                mat_A[126][3] * mat_B[223][1] +
                mat_A[127][0] * mat_B[231][1] +
                mat_A[127][1] * mat_B[239][1] +
                mat_A[127][2] * mat_B[247][1] +
                mat_A[127][3] * mat_B[255][1];
    mat_C[127][2] <=
                mat_A[120][0] * mat_B[7][2] +
                mat_A[120][1] * mat_B[15][2] +
                mat_A[120][2] * mat_B[23][2] +
                mat_A[120][3] * mat_B[31][2] +
                mat_A[121][0] * mat_B[39][2] +
                mat_A[121][1] * mat_B[47][2] +
                mat_A[121][2] * mat_B[55][2] +
                mat_A[121][3] * mat_B[63][2] +
                mat_A[122][0] * mat_B[71][2] +
                mat_A[122][1] * mat_B[79][2] +
                mat_A[122][2] * mat_B[87][2] +
                mat_A[122][3] * mat_B[95][2] +
                mat_A[123][0] * mat_B[103][2] +
                mat_A[123][1] * mat_B[111][2] +
                mat_A[123][2] * mat_B[119][2] +
                mat_A[123][3] * mat_B[127][2] +
                mat_A[124][0] * mat_B[135][2] +
                mat_A[124][1] * mat_B[143][2] +
                mat_A[124][2] * mat_B[151][2] +
                mat_A[124][3] * mat_B[159][2] +
                mat_A[125][0] * mat_B[167][2] +
                mat_A[125][1] * mat_B[175][2] +
                mat_A[125][2] * mat_B[183][2] +
                mat_A[125][3] * mat_B[191][2] +
                mat_A[126][0] * mat_B[199][2] +
                mat_A[126][1] * mat_B[207][2] +
                mat_A[126][2] * mat_B[215][2] +
                mat_A[126][3] * mat_B[223][2] +
                mat_A[127][0] * mat_B[231][2] +
                mat_A[127][1] * mat_B[239][2] +
                mat_A[127][2] * mat_B[247][2] +
                mat_A[127][3] * mat_B[255][2];
    mat_C[127][3] <=
                mat_A[120][0] * mat_B[7][3] +
                mat_A[120][1] * mat_B[15][3] +
                mat_A[120][2] * mat_B[23][3] +
                mat_A[120][3] * mat_B[31][3] +
                mat_A[121][0] * mat_B[39][3] +
                mat_A[121][1] * mat_B[47][3] +
                mat_A[121][2] * mat_B[55][3] +
                mat_A[121][3] * mat_B[63][3] +
                mat_A[122][0] * mat_B[71][3] +
                mat_A[122][1] * mat_B[79][3] +
                mat_A[122][2] * mat_B[87][3] +
                mat_A[122][3] * mat_B[95][3] +
                mat_A[123][0] * mat_B[103][3] +
                mat_A[123][1] * mat_B[111][3] +
                mat_A[123][2] * mat_B[119][3] +
                mat_A[123][3] * mat_B[127][3] +
                mat_A[124][0] * mat_B[135][3] +
                mat_A[124][1] * mat_B[143][3] +
                mat_A[124][2] * mat_B[151][3] +
                mat_A[124][3] * mat_B[159][3] +
                mat_A[125][0] * mat_B[167][3] +
                mat_A[125][1] * mat_B[175][3] +
                mat_A[125][2] * mat_B[183][3] +
                mat_A[125][3] * mat_B[191][3] +
                mat_A[126][0] * mat_B[199][3] +
                mat_A[126][1] * mat_B[207][3] +
                mat_A[126][2] * mat_B[215][3] +
                mat_A[126][3] * mat_B[223][3] +
                mat_A[127][0] * mat_B[231][3] +
                mat_A[127][1] * mat_B[239][3] +
                mat_A[127][2] * mat_B[247][3] +
                mat_A[127][3] * mat_B[255][3];
    mat_C[128][0] <=
                mat_A[128][0] * mat_B[0][0] +
                mat_A[128][1] * mat_B[8][0] +
                mat_A[128][2] * mat_B[16][0] +
                mat_A[128][3] * mat_B[24][0] +
                mat_A[129][0] * mat_B[32][0] +
                mat_A[129][1] * mat_B[40][0] +
                mat_A[129][2] * mat_B[48][0] +
                mat_A[129][3] * mat_B[56][0] +
                mat_A[130][0] * mat_B[64][0] +
                mat_A[130][1] * mat_B[72][0] +
                mat_A[130][2] * mat_B[80][0] +
                mat_A[130][3] * mat_B[88][0] +
                mat_A[131][0] * mat_B[96][0] +
                mat_A[131][1] * mat_B[104][0] +
                mat_A[131][2] * mat_B[112][0] +
                mat_A[131][3] * mat_B[120][0] +
                mat_A[132][0] * mat_B[128][0] +
                mat_A[132][1] * mat_B[136][0] +
                mat_A[132][2] * mat_B[144][0] +
                mat_A[132][3] * mat_B[152][0] +
                mat_A[133][0] * mat_B[160][0] +
                mat_A[133][1] * mat_B[168][0] +
                mat_A[133][2] * mat_B[176][0] +
                mat_A[133][3] * mat_B[184][0] +
                mat_A[134][0] * mat_B[192][0] +
                mat_A[134][1] * mat_B[200][0] +
                mat_A[134][2] * mat_B[208][0] +
                mat_A[134][3] * mat_B[216][0] +
                mat_A[135][0] * mat_B[224][0] +
                mat_A[135][1] * mat_B[232][0] +
                mat_A[135][2] * mat_B[240][0] +
                mat_A[135][3] * mat_B[248][0];
    mat_C[128][1] <=
                mat_A[128][0] * mat_B[0][1] +
                mat_A[128][1] * mat_B[8][1] +
                mat_A[128][2] * mat_B[16][1] +
                mat_A[128][3] * mat_B[24][1] +
                mat_A[129][0] * mat_B[32][1] +
                mat_A[129][1] * mat_B[40][1] +
                mat_A[129][2] * mat_B[48][1] +
                mat_A[129][3] * mat_B[56][1] +
                mat_A[130][0] * mat_B[64][1] +
                mat_A[130][1] * mat_B[72][1] +
                mat_A[130][2] * mat_B[80][1] +
                mat_A[130][3] * mat_B[88][1] +
                mat_A[131][0] * mat_B[96][1] +
                mat_A[131][1] * mat_B[104][1] +
                mat_A[131][2] * mat_B[112][1] +
                mat_A[131][3] * mat_B[120][1] +
                mat_A[132][0] * mat_B[128][1] +
                mat_A[132][1] * mat_B[136][1] +
                mat_A[132][2] * mat_B[144][1] +
                mat_A[132][3] * mat_B[152][1] +
                mat_A[133][0] * mat_B[160][1] +
                mat_A[133][1] * mat_B[168][1] +
                mat_A[133][2] * mat_B[176][1] +
                mat_A[133][3] * mat_B[184][1] +
                mat_A[134][0] * mat_B[192][1] +
                mat_A[134][1] * mat_B[200][1] +
                mat_A[134][2] * mat_B[208][1] +
                mat_A[134][3] * mat_B[216][1] +
                mat_A[135][0] * mat_B[224][1] +
                mat_A[135][1] * mat_B[232][1] +
                mat_A[135][2] * mat_B[240][1] +
                mat_A[135][3] * mat_B[248][1];
    mat_C[128][2] <=
                mat_A[128][0] * mat_B[0][2] +
                mat_A[128][1] * mat_B[8][2] +
                mat_A[128][2] * mat_B[16][2] +
                mat_A[128][3] * mat_B[24][2] +
                mat_A[129][0] * mat_B[32][2] +
                mat_A[129][1] * mat_B[40][2] +
                mat_A[129][2] * mat_B[48][2] +
                mat_A[129][3] * mat_B[56][2] +
                mat_A[130][0] * mat_B[64][2] +
                mat_A[130][1] * mat_B[72][2] +
                mat_A[130][2] * mat_B[80][2] +
                mat_A[130][3] * mat_B[88][2] +
                mat_A[131][0] * mat_B[96][2] +
                mat_A[131][1] * mat_B[104][2] +
                mat_A[131][2] * mat_B[112][2] +
                mat_A[131][3] * mat_B[120][2] +
                mat_A[132][0] * mat_B[128][2] +
                mat_A[132][1] * mat_B[136][2] +
                mat_A[132][2] * mat_B[144][2] +
                mat_A[132][3] * mat_B[152][2] +
                mat_A[133][0] * mat_B[160][2] +
                mat_A[133][1] * mat_B[168][2] +
                mat_A[133][2] * mat_B[176][2] +
                mat_A[133][3] * mat_B[184][2] +
                mat_A[134][0] * mat_B[192][2] +
                mat_A[134][1] * mat_B[200][2] +
                mat_A[134][2] * mat_B[208][2] +
                mat_A[134][3] * mat_B[216][2] +
                mat_A[135][0] * mat_B[224][2] +
                mat_A[135][1] * mat_B[232][2] +
                mat_A[135][2] * mat_B[240][2] +
                mat_A[135][3] * mat_B[248][2];
    mat_C[128][3] <=
                mat_A[128][0] * mat_B[0][3] +
                mat_A[128][1] * mat_B[8][3] +
                mat_A[128][2] * mat_B[16][3] +
                mat_A[128][3] * mat_B[24][3] +
                mat_A[129][0] * mat_B[32][3] +
                mat_A[129][1] * mat_B[40][3] +
                mat_A[129][2] * mat_B[48][3] +
                mat_A[129][3] * mat_B[56][3] +
                mat_A[130][0] * mat_B[64][3] +
                mat_A[130][1] * mat_B[72][3] +
                mat_A[130][2] * mat_B[80][3] +
                mat_A[130][3] * mat_B[88][3] +
                mat_A[131][0] * mat_B[96][3] +
                mat_A[131][1] * mat_B[104][3] +
                mat_A[131][2] * mat_B[112][3] +
                mat_A[131][3] * mat_B[120][3] +
                mat_A[132][0] * mat_B[128][3] +
                mat_A[132][1] * mat_B[136][3] +
                mat_A[132][2] * mat_B[144][3] +
                mat_A[132][3] * mat_B[152][3] +
                mat_A[133][0] * mat_B[160][3] +
                mat_A[133][1] * mat_B[168][3] +
                mat_A[133][2] * mat_B[176][3] +
                mat_A[133][3] * mat_B[184][3] +
                mat_A[134][0] * mat_B[192][3] +
                mat_A[134][1] * mat_B[200][3] +
                mat_A[134][2] * mat_B[208][3] +
                mat_A[134][3] * mat_B[216][3] +
                mat_A[135][0] * mat_B[224][3] +
                mat_A[135][1] * mat_B[232][3] +
                mat_A[135][2] * mat_B[240][3] +
                mat_A[135][3] * mat_B[248][3];
    mat_C[129][0] <=
                mat_A[128][0] * mat_B[1][0] +
                mat_A[128][1] * mat_B[9][0] +
                mat_A[128][2] * mat_B[17][0] +
                mat_A[128][3] * mat_B[25][0] +
                mat_A[129][0] * mat_B[33][0] +
                mat_A[129][1] * mat_B[41][0] +
                mat_A[129][2] * mat_B[49][0] +
                mat_A[129][3] * mat_B[57][0] +
                mat_A[130][0] * mat_B[65][0] +
                mat_A[130][1] * mat_B[73][0] +
                mat_A[130][2] * mat_B[81][0] +
                mat_A[130][3] * mat_B[89][0] +
                mat_A[131][0] * mat_B[97][0] +
                mat_A[131][1] * mat_B[105][0] +
                mat_A[131][2] * mat_B[113][0] +
                mat_A[131][3] * mat_B[121][0] +
                mat_A[132][0] * mat_B[129][0] +
                mat_A[132][1] * mat_B[137][0] +
                mat_A[132][2] * mat_B[145][0] +
                mat_A[132][3] * mat_B[153][0] +
                mat_A[133][0] * mat_B[161][0] +
                mat_A[133][1] * mat_B[169][0] +
                mat_A[133][2] * mat_B[177][0] +
                mat_A[133][3] * mat_B[185][0] +
                mat_A[134][0] * mat_B[193][0] +
                mat_A[134][1] * mat_B[201][0] +
                mat_A[134][2] * mat_B[209][0] +
                mat_A[134][3] * mat_B[217][0] +
                mat_A[135][0] * mat_B[225][0] +
                mat_A[135][1] * mat_B[233][0] +
                mat_A[135][2] * mat_B[241][0] +
                mat_A[135][3] * mat_B[249][0];
    mat_C[129][1] <=
                mat_A[128][0] * mat_B[1][1] +
                mat_A[128][1] * mat_B[9][1] +
                mat_A[128][2] * mat_B[17][1] +
                mat_A[128][3] * mat_B[25][1] +
                mat_A[129][0] * mat_B[33][1] +
                mat_A[129][1] * mat_B[41][1] +
                mat_A[129][2] * mat_B[49][1] +
                mat_A[129][3] * mat_B[57][1] +
                mat_A[130][0] * mat_B[65][1] +
                mat_A[130][1] * mat_B[73][1] +
                mat_A[130][2] * mat_B[81][1] +
                mat_A[130][3] * mat_B[89][1] +
                mat_A[131][0] * mat_B[97][1] +
                mat_A[131][1] * mat_B[105][1] +
                mat_A[131][2] * mat_B[113][1] +
                mat_A[131][3] * mat_B[121][1] +
                mat_A[132][0] * mat_B[129][1] +
                mat_A[132][1] * mat_B[137][1] +
                mat_A[132][2] * mat_B[145][1] +
                mat_A[132][3] * mat_B[153][1] +
                mat_A[133][0] * mat_B[161][1] +
                mat_A[133][1] * mat_B[169][1] +
                mat_A[133][2] * mat_B[177][1] +
                mat_A[133][3] * mat_B[185][1] +
                mat_A[134][0] * mat_B[193][1] +
                mat_A[134][1] * mat_B[201][1] +
                mat_A[134][2] * mat_B[209][1] +
                mat_A[134][3] * mat_B[217][1] +
                mat_A[135][0] * mat_B[225][1] +
                mat_A[135][1] * mat_B[233][1] +
                mat_A[135][2] * mat_B[241][1] +
                mat_A[135][3] * mat_B[249][1];
    mat_C[129][2] <=
                mat_A[128][0] * mat_B[1][2] +
                mat_A[128][1] * mat_B[9][2] +
                mat_A[128][2] * mat_B[17][2] +
                mat_A[128][3] * mat_B[25][2] +
                mat_A[129][0] * mat_B[33][2] +
                mat_A[129][1] * mat_B[41][2] +
                mat_A[129][2] * mat_B[49][2] +
                mat_A[129][3] * mat_B[57][2] +
                mat_A[130][0] * mat_B[65][2] +
                mat_A[130][1] * mat_B[73][2] +
                mat_A[130][2] * mat_B[81][2] +
                mat_A[130][3] * mat_B[89][2] +
                mat_A[131][0] * mat_B[97][2] +
                mat_A[131][1] * mat_B[105][2] +
                mat_A[131][2] * mat_B[113][2] +
                mat_A[131][3] * mat_B[121][2] +
                mat_A[132][0] * mat_B[129][2] +
                mat_A[132][1] * mat_B[137][2] +
                mat_A[132][2] * mat_B[145][2] +
                mat_A[132][3] * mat_B[153][2] +
                mat_A[133][0] * mat_B[161][2] +
                mat_A[133][1] * mat_B[169][2] +
                mat_A[133][2] * mat_B[177][2] +
                mat_A[133][3] * mat_B[185][2] +
                mat_A[134][0] * mat_B[193][2] +
                mat_A[134][1] * mat_B[201][2] +
                mat_A[134][2] * mat_B[209][2] +
                mat_A[134][3] * mat_B[217][2] +
                mat_A[135][0] * mat_B[225][2] +
                mat_A[135][1] * mat_B[233][2] +
                mat_A[135][2] * mat_B[241][2] +
                mat_A[135][3] * mat_B[249][2];
    mat_C[129][3] <=
                mat_A[128][0] * mat_B[1][3] +
                mat_A[128][1] * mat_B[9][3] +
                mat_A[128][2] * mat_B[17][3] +
                mat_A[128][3] * mat_B[25][3] +
                mat_A[129][0] * mat_B[33][3] +
                mat_A[129][1] * mat_B[41][3] +
                mat_A[129][2] * mat_B[49][3] +
                mat_A[129][3] * mat_B[57][3] +
                mat_A[130][0] * mat_B[65][3] +
                mat_A[130][1] * mat_B[73][3] +
                mat_A[130][2] * mat_B[81][3] +
                mat_A[130][3] * mat_B[89][3] +
                mat_A[131][0] * mat_B[97][3] +
                mat_A[131][1] * mat_B[105][3] +
                mat_A[131][2] * mat_B[113][3] +
                mat_A[131][3] * mat_B[121][3] +
                mat_A[132][0] * mat_B[129][3] +
                mat_A[132][1] * mat_B[137][3] +
                mat_A[132][2] * mat_B[145][3] +
                mat_A[132][3] * mat_B[153][3] +
                mat_A[133][0] * mat_B[161][3] +
                mat_A[133][1] * mat_B[169][3] +
                mat_A[133][2] * mat_B[177][3] +
                mat_A[133][3] * mat_B[185][3] +
                mat_A[134][0] * mat_B[193][3] +
                mat_A[134][1] * mat_B[201][3] +
                mat_A[134][2] * mat_B[209][3] +
                mat_A[134][3] * mat_B[217][3] +
                mat_A[135][0] * mat_B[225][3] +
                mat_A[135][1] * mat_B[233][3] +
                mat_A[135][2] * mat_B[241][3] +
                mat_A[135][3] * mat_B[249][3];
    mat_C[130][0] <=
                mat_A[128][0] * mat_B[2][0] +
                mat_A[128][1] * mat_B[10][0] +
                mat_A[128][2] * mat_B[18][0] +
                mat_A[128][3] * mat_B[26][0] +
                mat_A[129][0] * mat_B[34][0] +
                mat_A[129][1] * mat_B[42][0] +
                mat_A[129][2] * mat_B[50][0] +
                mat_A[129][3] * mat_B[58][0] +
                mat_A[130][0] * mat_B[66][0] +
                mat_A[130][1] * mat_B[74][0] +
                mat_A[130][2] * mat_B[82][0] +
                mat_A[130][3] * mat_B[90][0] +
                mat_A[131][0] * mat_B[98][0] +
                mat_A[131][1] * mat_B[106][0] +
                mat_A[131][2] * mat_B[114][0] +
                mat_A[131][3] * mat_B[122][0] +
                mat_A[132][0] * mat_B[130][0] +
                mat_A[132][1] * mat_B[138][0] +
                mat_A[132][2] * mat_B[146][0] +
                mat_A[132][3] * mat_B[154][0] +
                mat_A[133][0] * mat_B[162][0] +
                mat_A[133][1] * mat_B[170][0] +
                mat_A[133][2] * mat_B[178][0] +
                mat_A[133][3] * mat_B[186][0] +
                mat_A[134][0] * mat_B[194][0] +
                mat_A[134][1] * mat_B[202][0] +
                mat_A[134][2] * mat_B[210][0] +
                mat_A[134][3] * mat_B[218][0] +
                mat_A[135][0] * mat_B[226][0] +
                mat_A[135][1] * mat_B[234][0] +
                mat_A[135][2] * mat_B[242][0] +
                mat_A[135][3] * mat_B[250][0];
    mat_C[130][1] <=
                mat_A[128][0] * mat_B[2][1] +
                mat_A[128][1] * mat_B[10][1] +
                mat_A[128][2] * mat_B[18][1] +
                mat_A[128][3] * mat_B[26][1] +
                mat_A[129][0] * mat_B[34][1] +
                mat_A[129][1] * mat_B[42][1] +
                mat_A[129][2] * mat_B[50][1] +
                mat_A[129][3] * mat_B[58][1] +
                mat_A[130][0] * mat_B[66][1] +
                mat_A[130][1] * mat_B[74][1] +
                mat_A[130][2] * mat_B[82][1] +
                mat_A[130][3] * mat_B[90][1] +
                mat_A[131][0] * mat_B[98][1] +
                mat_A[131][1] * mat_B[106][1] +
                mat_A[131][2] * mat_B[114][1] +
                mat_A[131][3] * mat_B[122][1] +
                mat_A[132][0] * mat_B[130][1] +
                mat_A[132][1] * mat_B[138][1] +
                mat_A[132][2] * mat_B[146][1] +
                mat_A[132][3] * mat_B[154][1] +
                mat_A[133][0] * mat_B[162][1] +
                mat_A[133][1] * mat_B[170][1] +
                mat_A[133][2] * mat_B[178][1] +
                mat_A[133][3] * mat_B[186][1] +
                mat_A[134][0] * mat_B[194][1] +
                mat_A[134][1] * mat_B[202][1] +
                mat_A[134][2] * mat_B[210][1] +
                mat_A[134][3] * mat_B[218][1] +
                mat_A[135][0] * mat_B[226][1] +
                mat_A[135][1] * mat_B[234][1] +
                mat_A[135][2] * mat_B[242][1] +
                mat_A[135][3] * mat_B[250][1];
    mat_C[130][2] <=
                mat_A[128][0] * mat_B[2][2] +
                mat_A[128][1] * mat_B[10][2] +
                mat_A[128][2] * mat_B[18][2] +
                mat_A[128][3] * mat_B[26][2] +
                mat_A[129][0] * mat_B[34][2] +
                mat_A[129][1] * mat_B[42][2] +
                mat_A[129][2] * mat_B[50][2] +
                mat_A[129][3] * mat_B[58][2] +
                mat_A[130][0] * mat_B[66][2] +
                mat_A[130][1] * mat_B[74][2] +
                mat_A[130][2] * mat_B[82][2] +
                mat_A[130][3] * mat_B[90][2] +
                mat_A[131][0] * mat_B[98][2] +
                mat_A[131][1] * mat_B[106][2] +
                mat_A[131][2] * mat_B[114][2] +
                mat_A[131][3] * mat_B[122][2] +
                mat_A[132][0] * mat_B[130][2] +
                mat_A[132][1] * mat_B[138][2] +
                mat_A[132][2] * mat_B[146][2] +
                mat_A[132][3] * mat_B[154][2] +
                mat_A[133][0] * mat_B[162][2] +
                mat_A[133][1] * mat_B[170][2] +
                mat_A[133][2] * mat_B[178][2] +
                mat_A[133][3] * mat_B[186][2] +
                mat_A[134][0] * mat_B[194][2] +
                mat_A[134][1] * mat_B[202][2] +
                mat_A[134][2] * mat_B[210][2] +
                mat_A[134][3] * mat_B[218][2] +
                mat_A[135][0] * mat_B[226][2] +
                mat_A[135][1] * mat_B[234][2] +
                mat_A[135][2] * mat_B[242][2] +
                mat_A[135][3] * mat_B[250][2];
    mat_C[130][3] <=
                mat_A[128][0] * mat_B[2][3] +
                mat_A[128][1] * mat_B[10][3] +
                mat_A[128][2] * mat_B[18][3] +
                mat_A[128][3] * mat_B[26][3] +
                mat_A[129][0] * mat_B[34][3] +
                mat_A[129][1] * mat_B[42][3] +
                mat_A[129][2] * mat_B[50][3] +
                mat_A[129][3] * mat_B[58][3] +
                mat_A[130][0] * mat_B[66][3] +
                mat_A[130][1] * mat_B[74][3] +
                mat_A[130][2] * mat_B[82][3] +
                mat_A[130][3] * mat_B[90][3] +
                mat_A[131][0] * mat_B[98][3] +
                mat_A[131][1] * mat_B[106][3] +
                mat_A[131][2] * mat_B[114][3] +
                mat_A[131][3] * mat_B[122][3] +
                mat_A[132][0] * mat_B[130][3] +
                mat_A[132][1] * mat_B[138][3] +
                mat_A[132][2] * mat_B[146][3] +
                mat_A[132][3] * mat_B[154][3] +
                mat_A[133][0] * mat_B[162][3] +
                mat_A[133][1] * mat_B[170][3] +
                mat_A[133][2] * mat_B[178][3] +
                mat_A[133][3] * mat_B[186][3] +
                mat_A[134][0] * mat_B[194][3] +
                mat_A[134][1] * mat_B[202][3] +
                mat_A[134][2] * mat_B[210][3] +
                mat_A[134][3] * mat_B[218][3] +
                mat_A[135][0] * mat_B[226][3] +
                mat_A[135][1] * mat_B[234][3] +
                mat_A[135][2] * mat_B[242][3] +
                mat_A[135][3] * mat_B[250][3];
    mat_C[131][0] <=
                mat_A[128][0] * mat_B[3][0] +
                mat_A[128][1] * mat_B[11][0] +
                mat_A[128][2] * mat_B[19][0] +
                mat_A[128][3] * mat_B[27][0] +
                mat_A[129][0] * mat_B[35][0] +
                mat_A[129][1] * mat_B[43][0] +
                mat_A[129][2] * mat_B[51][0] +
                mat_A[129][3] * mat_B[59][0] +
                mat_A[130][0] * mat_B[67][0] +
                mat_A[130][1] * mat_B[75][0] +
                mat_A[130][2] * mat_B[83][0] +
                mat_A[130][3] * mat_B[91][0] +
                mat_A[131][0] * mat_B[99][0] +
                mat_A[131][1] * mat_B[107][0] +
                mat_A[131][2] * mat_B[115][0] +
                mat_A[131][3] * mat_B[123][0] +
                mat_A[132][0] * mat_B[131][0] +
                mat_A[132][1] * mat_B[139][0] +
                mat_A[132][2] * mat_B[147][0] +
                mat_A[132][3] * mat_B[155][0] +
                mat_A[133][0] * mat_B[163][0] +
                mat_A[133][1] * mat_B[171][0] +
                mat_A[133][2] * mat_B[179][0] +
                mat_A[133][3] * mat_B[187][0] +
                mat_A[134][0] * mat_B[195][0] +
                mat_A[134][1] * mat_B[203][0] +
                mat_A[134][2] * mat_B[211][0] +
                mat_A[134][3] * mat_B[219][0] +
                mat_A[135][0] * mat_B[227][0] +
                mat_A[135][1] * mat_B[235][0] +
                mat_A[135][2] * mat_B[243][0] +
                mat_A[135][3] * mat_B[251][0];
    mat_C[131][1] <=
                mat_A[128][0] * mat_B[3][1] +
                mat_A[128][1] * mat_B[11][1] +
                mat_A[128][2] * mat_B[19][1] +
                mat_A[128][3] * mat_B[27][1] +
                mat_A[129][0] * mat_B[35][1] +
                mat_A[129][1] * mat_B[43][1] +
                mat_A[129][2] * mat_B[51][1] +
                mat_A[129][3] * mat_B[59][1] +
                mat_A[130][0] * mat_B[67][1] +
                mat_A[130][1] * mat_B[75][1] +
                mat_A[130][2] * mat_B[83][1] +
                mat_A[130][3] * mat_B[91][1] +
                mat_A[131][0] * mat_B[99][1] +
                mat_A[131][1] * mat_B[107][1] +
                mat_A[131][2] * mat_B[115][1] +
                mat_A[131][3] * mat_B[123][1] +
                mat_A[132][0] * mat_B[131][1] +
                mat_A[132][1] * mat_B[139][1] +
                mat_A[132][2] * mat_B[147][1] +
                mat_A[132][3] * mat_B[155][1] +
                mat_A[133][0] * mat_B[163][1] +
                mat_A[133][1] * mat_B[171][1] +
                mat_A[133][2] * mat_B[179][1] +
                mat_A[133][3] * mat_B[187][1] +
                mat_A[134][0] * mat_B[195][1] +
                mat_A[134][1] * mat_B[203][1] +
                mat_A[134][2] * mat_B[211][1] +
                mat_A[134][3] * mat_B[219][1] +
                mat_A[135][0] * mat_B[227][1] +
                mat_A[135][1] * mat_B[235][1] +
                mat_A[135][2] * mat_B[243][1] +
                mat_A[135][3] * mat_B[251][1];
    mat_C[131][2] <=
                mat_A[128][0] * mat_B[3][2] +
                mat_A[128][1] * mat_B[11][2] +
                mat_A[128][2] * mat_B[19][2] +
                mat_A[128][3] * mat_B[27][2] +
                mat_A[129][0] * mat_B[35][2] +
                mat_A[129][1] * mat_B[43][2] +
                mat_A[129][2] * mat_B[51][2] +
                mat_A[129][3] * mat_B[59][2] +
                mat_A[130][0] * mat_B[67][2] +
                mat_A[130][1] * mat_B[75][2] +
                mat_A[130][2] * mat_B[83][2] +
                mat_A[130][3] * mat_B[91][2] +
                mat_A[131][0] * mat_B[99][2] +
                mat_A[131][1] * mat_B[107][2] +
                mat_A[131][2] * mat_B[115][2] +
                mat_A[131][3] * mat_B[123][2] +
                mat_A[132][0] * mat_B[131][2] +
                mat_A[132][1] * mat_B[139][2] +
                mat_A[132][2] * mat_B[147][2] +
                mat_A[132][3] * mat_B[155][2] +
                mat_A[133][0] * mat_B[163][2] +
                mat_A[133][1] * mat_B[171][2] +
                mat_A[133][2] * mat_B[179][2] +
                mat_A[133][3] * mat_B[187][2] +
                mat_A[134][0] * mat_B[195][2] +
                mat_A[134][1] * mat_B[203][2] +
                mat_A[134][2] * mat_B[211][2] +
                mat_A[134][3] * mat_B[219][2] +
                mat_A[135][0] * mat_B[227][2] +
                mat_A[135][1] * mat_B[235][2] +
                mat_A[135][2] * mat_B[243][2] +
                mat_A[135][3] * mat_B[251][2];
    mat_C[131][3] <=
                mat_A[128][0] * mat_B[3][3] +
                mat_A[128][1] * mat_B[11][3] +
                mat_A[128][2] * mat_B[19][3] +
                mat_A[128][3] * mat_B[27][3] +
                mat_A[129][0] * mat_B[35][3] +
                mat_A[129][1] * mat_B[43][3] +
                mat_A[129][2] * mat_B[51][3] +
                mat_A[129][3] * mat_B[59][3] +
                mat_A[130][0] * mat_B[67][3] +
                mat_A[130][1] * mat_B[75][3] +
                mat_A[130][2] * mat_B[83][3] +
                mat_A[130][3] * mat_B[91][3] +
                mat_A[131][0] * mat_B[99][3] +
                mat_A[131][1] * mat_B[107][3] +
                mat_A[131][2] * mat_B[115][3] +
                mat_A[131][3] * mat_B[123][3] +
                mat_A[132][0] * mat_B[131][3] +
                mat_A[132][1] * mat_B[139][3] +
                mat_A[132][2] * mat_B[147][3] +
                mat_A[132][3] * mat_B[155][3] +
                mat_A[133][0] * mat_B[163][3] +
                mat_A[133][1] * mat_B[171][3] +
                mat_A[133][2] * mat_B[179][3] +
                mat_A[133][3] * mat_B[187][3] +
                mat_A[134][0] * mat_B[195][3] +
                mat_A[134][1] * mat_B[203][3] +
                mat_A[134][2] * mat_B[211][3] +
                mat_A[134][3] * mat_B[219][3] +
                mat_A[135][0] * mat_B[227][3] +
                mat_A[135][1] * mat_B[235][3] +
                mat_A[135][2] * mat_B[243][3] +
                mat_A[135][3] * mat_B[251][3];
    mat_C[132][0] <=
                mat_A[128][0] * mat_B[4][0] +
                mat_A[128][1] * mat_B[12][0] +
                mat_A[128][2] * mat_B[20][0] +
                mat_A[128][3] * mat_B[28][0] +
                mat_A[129][0] * mat_B[36][0] +
                mat_A[129][1] * mat_B[44][0] +
                mat_A[129][2] * mat_B[52][0] +
                mat_A[129][3] * mat_B[60][0] +
                mat_A[130][0] * mat_B[68][0] +
                mat_A[130][1] * mat_B[76][0] +
                mat_A[130][2] * mat_B[84][0] +
                mat_A[130][3] * mat_B[92][0] +
                mat_A[131][0] * mat_B[100][0] +
                mat_A[131][1] * mat_B[108][0] +
                mat_A[131][2] * mat_B[116][0] +
                mat_A[131][3] * mat_B[124][0] +
                mat_A[132][0] * mat_B[132][0] +
                mat_A[132][1] * mat_B[140][0] +
                mat_A[132][2] * mat_B[148][0] +
                mat_A[132][3] * mat_B[156][0] +
                mat_A[133][0] * mat_B[164][0] +
                mat_A[133][1] * mat_B[172][0] +
                mat_A[133][2] * mat_B[180][0] +
                mat_A[133][3] * mat_B[188][0] +
                mat_A[134][0] * mat_B[196][0] +
                mat_A[134][1] * mat_B[204][0] +
                mat_A[134][2] * mat_B[212][0] +
                mat_A[134][3] * mat_B[220][0] +
                mat_A[135][0] * mat_B[228][0] +
                mat_A[135][1] * mat_B[236][0] +
                mat_A[135][2] * mat_B[244][0] +
                mat_A[135][3] * mat_B[252][0];
    mat_C[132][1] <=
                mat_A[128][0] * mat_B[4][1] +
                mat_A[128][1] * mat_B[12][1] +
                mat_A[128][2] * mat_B[20][1] +
                mat_A[128][3] * mat_B[28][1] +
                mat_A[129][0] * mat_B[36][1] +
                mat_A[129][1] * mat_B[44][1] +
                mat_A[129][2] * mat_B[52][1] +
                mat_A[129][3] * mat_B[60][1] +
                mat_A[130][0] * mat_B[68][1] +
                mat_A[130][1] * mat_B[76][1] +
                mat_A[130][2] * mat_B[84][1] +
                mat_A[130][3] * mat_B[92][1] +
                mat_A[131][0] * mat_B[100][1] +
                mat_A[131][1] * mat_B[108][1] +
                mat_A[131][2] * mat_B[116][1] +
                mat_A[131][3] * mat_B[124][1] +
                mat_A[132][0] * mat_B[132][1] +
                mat_A[132][1] * mat_B[140][1] +
                mat_A[132][2] * mat_B[148][1] +
                mat_A[132][3] * mat_B[156][1] +
                mat_A[133][0] * mat_B[164][1] +
                mat_A[133][1] * mat_B[172][1] +
                mat_A[133][2] * mat_B[180][1] +
                mat_A[133][3] * mat_B[188][1] +
                mat_A[134][0] * mat_B[196][1] +
                mat_A[134][1] * mat_B[204][1] +
                mat_A[134][2] * mat_B[212][1] +
                mat_A[134][3] * mat_B[220][1] +
                mat_A[135][0] * mat_B[228][1] +
                mat_A[135][1] * mat_B[236][1] +
                mat_A[135][2] * mat_B[244][1] +
                mat_A[135][3] * mat_B[252][1];
    mat_C[132][2] <=
                mat_A[128][0] * mat_B[4][2] +
                mat_A[128][1] * mat_B[12][2] +
                mat_A[128][2] * mat_B[20][2] +
                mat_A[128][3] * mat_B[28][2] +
                mat_A[129][0] * mat_B[36][2] +
                mat_A[129][1] * mat_B[44][2] +
                mat_A[129][2] * mat_B[52][2] +
                mat_A[129][3] * mat_B[60][2] +
                mat_A[130][0] * mat_B[68][2] +
                mat_A[130][1] * mat_B[76][2] +
                mat_A[130][2] * mat_B[84][2] +
                mat_A[130][3] * mat_B[92][2] +
                mat_A[131][0] * mat_B[100][2] +
                mat_A[131][1] * mat_B[108][2] +
                mat_A[131][2] * mat_B[116][2] +
                mat_A[131][3] * mat_B[124][2] +
                mat_A[132][0] * mat_B[132][2] +
                mat_A[132][1] * mat_B[140][2] +
                mat_A[132][2] * mat_B[148][2] +
                mat_A[132][3] * mat_B[156][2] +
                mat_A[133][0] * mat_B[164][2] +
                mat_A[133][1] * mat_B[172][2] +
                mat_A[133][2] * mat_B[180][2] +
                mat_A[133][3] * mat_B[188][2] +
                mat_A[134][0] * mat_B[196][2] +
                mat_A[134][1] * mat_B[204][2] +
                mat_A[134][2] * mat_B[212][2] +
                mat_A[134][3] * mat_B[220][2] +
                mat_A[135][0] * mat_B[228][2] +
                mat_A[135][1] * mat_B[236][2] +
                mat_A[135][2] * mat_B[244][2] +
                mat_A[135][3] * mat_B[252][2];
    mat_C[132][3] <=
                mat_A[128][0] * mat_B[4][3] +
                mat_A[128][1] * mat_B[12][3] +
                mat_A[128][2] * mat_B[20][3] +
                mat_A[128][3] * mat_B[28][3] +
                mat_A[129][0] * mat_B[36][3] +
                mat_A[129][1] * mat_B[44][3] +
                mat_A[129][2] * mat_B[52][3] +
                mat_A[129][3] * mat_B[60][3] +
                mat_A[130][0] * mat_B[68][3] +
                mat_A[130][1] * mat_B[76][3] +
                mat_A[130][2] * mat_B[84][3] +
                mat_A[130][3] * mat_B[92][3] +
                mat_A[131][0] * mat_B[100][3] +
                mat_A[131][1] * mat_B[108][3] +
                mat_A[131][2] * mat_B[116][3] +
                mat_A[131][3] * mat_B[124][3] +
                mat_A[132][0] * mat_B[132][3] +
                mat_A[132][1] * mat_B[140][3] +
                mat_A[132][2] * mat_B[148][3] +
                mat_A[132][3] * mat_B[156][3] +
                mat_A[133][0] * mat_B[164][3] +
                mat_A[133][1] * mat_B[172][3] +
                mat_A[133][2] * mat_B[180][3] +
                mat_A[133][3] * mat_B[188][3] +
                mat_A[134][0] * mat_B[196][3] +
                mat_A[134][1] * mat_B[204][3] +
                mat_A[134][2] * mat_B[212][3] +
                mat_A[134][3] * mat_B[220][3] +
                mat_A[135][0] * mat_B[228][3] +
                mat_A[135][1] * mat_B[236][3] +
                mat_A[135][2] * mat_B[244][3] +
                mat_A[135][3] * mat_B[252][3];
    mat_C[133][0] <=
                mat_A[128][0] * mat_B[5][0] +
                mat_A[128][1] * mat_B[13][0] +
                mat_A[128][2] * mat_B[21][0] +
                mat_A[128][3] * mat_B[29][0] +
                mat_A[129][0] * mat_B[37][0] +
                mat_A[129][1] * mat_B[45][0] +
                mat_A[129][2] * mat_B[53][0] +
                mat_A[129][3] * mat_B[61][0] +
                mat_A[130][0] * mat_B[69][0] +
                mat_A[130][1] * mat_B[77][0] +
                mat_A[130][2] * mat_B[85][0] +
                mat_A[130][3] * mat_B[93][0] +
                mat_A[131][0] * mat_B[101][0] +
                mat_A[131][1] * mat_B[109][0] +
                mat_A[131][2] * mat_B[117][0] +
                mat_A[131][3] * mat_B[125][0] +
                mat_A[132][0] * mat_B[133][0] +
                mat_A[132][1] * mat_B[141][0] +
                mat_A[132][2] * mat_B[149][0] +
                mat_A[132][3] * mat_B[157][0] +
                mat_A[133][0] * mat_B[165][0] +
                mat_A[133][1] * mat_B[173][0] +
                mat_A[133][2] * mat_B[181][0] +
                mat_A[133][3] * mat_B[189][0] +
                mat_A[134][0] * mat_B[197][0] +
                mat_A[134][1] * mat_B[205][0] +
                mat_A[134][2] * mat_B[213][0] +
                mat_A[134][3] * mat_B[221][0] +
                mat_A[135][0] * mat_B[229][0] +
                mat_A[135][1] * mat_B[237][0] +
                mat_A[135][2] * mat_B[245][0] +
                mat_A[135][3] * mat_B[253][0];
    mat_C[133][1] <=
                mat_A[128][0] * mat_B[5][1] +
                mat_A[128][1] * mat_B[13][1] +
                mat_A[128][2] * mat_B[21][1] +
                mat_A[128][3] * mat_B[29][1] +
                mat_A[129][0] * mat_B[37][1] +
                mat_A[129][1] * mat_B[45][1] +
                mat_A[129][2] * mat_B[53][1] +
                mat_A[129][3] * mat_B[61][1] +
                mat_A[130][0] * mat_B[69][1] +
                mat_A[130][1] * mat_B[77][1] +
                mat_A[130][2] * mat_B[85][1] +
                mat_A[130][3] * mat_B[93][1] +
                mat_A[131][0] * mat_B[101][1] +
                mat_A[131][1] * mat_B[109][1] +
                mat_A[131][2] * mat_B[117][1] +
                mat_A[131][3] * mat_B[125][1] +
                mat_A[132][0] * mat_B[133][1] +
                mat_A[132][1] * mat_B[141][1] +
                mat_A[132][2] * mat_B[149][1] +
                mat_A[132][3] * mat_B[157][1] +
                mat_A[133][0] * mat_B[165][1] +
                mat_A[133][1] * mat_B[173][1] +
                mat_A[133][2] * mat_B[181][1] +
                mat_A[133][3] * mat_B[189][1] +
                mat_A[134][0] * mat_B[197][1] +
                mat_A[134][1] * mat_B[205][1] +
                mat_A[134][2] * mat_B[213][1] +
                mat_A[134][3] * mat_B[221][1] +
                mat_A[135][0] * mat_B[229][1] +
                mat_A[135][1] * mat_B[237][1] +
                mat_A[135][2] * mat_B[245][1] +
                mat_A[135][3] * mat_B[253][1];
    mat_C[133][2] <=
                mat_A[128][0] * mat_B[5][2] +
                mat_A[128][1] * mat_B[13][2] +
                mat_A[128][2] * mat_B[21][2] +
                mat_A[128][3] * mat_B[29][2] +
                mat_A[129][0] * mat_B[37][2] +
                mat_A[129][1] * mat_B[45][2] +
                mat_A[129][2] * mat_B[53][2] +
                mat_A[129][3] * mat_B[61][2] +
                mat_A[130][0] * mat_B[69][2] +
                mat_A[130][1] * mat_B[77][2] +
                mat_A[130][2] * mat_B[85][2] +
                mat_A[130][3] * mat_B[93][2] +
                mat_A[131][0] * mat_B[101][2] +
                mat_A[131][1] * mat_B[109][2] +
                mat_A[131][2] * mat_B[117][2] +
                mat_A[131][3] * mat_B[125][2] +
                mat_A[132][0] * mat_B[133][2] +
                mat_A[132][1] * mat_B[141][2] +
                mat_A[132][2] * mat_B[149][2] +
                mat_A[132][3] * mat_B[157][2] +
                mat_A[133][0] * mat_B[165][2] +
                mat_A[133][1] * mat_B[173][2] +
                mat_A[133][2] * mat_B[181][2] +
                mat_A[133][3] * mat_B[189][2] +
                mat_A[134][0] * mat_B[197][2] +
                mat_A[134][1] * mat_B[205][2] +
                mat_A[134][2] * mat_B[213][2] +
                mat_A[134][3] * mat_B[221][2] +
                mat_A[135][0] * mat_B[229][2] +
                mat_A[135][1] * mat_B[237][2] +
                mat_A[135][2] * mat_B[245][2] +
                mat_A[135][3] * mat_B[253][2];
    mat_C[133][3] <=
                mat_A[128][0] * mat_B[5][3] +
                mat_A[128][1] * mat_B[13][3] +
                mat_A[128][2] * mat_B[21][3] +
                mat_A[128][3] * mat_B[29][3] +
                mat_A[129][0] * mat_B[37][3] +
                mat_A[129][1] * mat_B[45][3] +
                mat_A[129][2] * mat_B[53][3] +
                mat_A[129][3] * mat_B[61][3] +
                mat_A[130][0] * mat_B[69][3] +
                mat_A[130][1] * mat_B[77][3] +
                mat_A[130][2] * mat_B[85][3] +
                mat_A[130][3] * mat_B[93][3] +
                mat_A[131][0] * mat_B[101][3] +
                mat_A[131][1] * mat_B[109][3] +
                mat_A[131][2] * mat_B[117][3] +
                mat_A[131][3] * mat_B[125][3] +
                mat_A[132][0] * mat_B[133][3] +
                mat_A[132][1] * mat_B[141][3] +
                mat_A[132][2] * mat_B[149][3] +
                mat_A[132][3] * mat_B[157][3] +
                mat_A[133][0] * mat_B[165][3] +
                mat_A[133][1] * mat_B[173][3] +
                mat_A[133][2] * mat_B[181][3] +
                mat_A[133][3] * mat_B[189][3] +
                mat_A[134][0] * mat_B[197][3] +
                mat_A[134][1] * mat_B[205][3] +
                mat_A[134][2] * mat_B[213][3] +
                mat_A[134][3] * mat_B[221][3] +
                mat_A[135][0] * mat_B[229][3] +
                mat_A[135][1] * mat_B[237][3] +
                mat_A[135][2] * mat_B[245][3] +
                mat_A[135][3] * mat_B[253][3];
    mat_C[134][0] <=
                mat_A[128][0] * mat_B[6][0] +
                mat_A[128][1] * mat_B[14][0] +
                mat_A[128][2] * mat_B[22][0] +
                mat_A[128][3] * mat_B[30][0] +
                mat_A[129][0] * mat_B[38][0] +
                mat_A[129][1] * mat_B[46][0] +
                mat_A[129][2] * mat_B[54][0] +
                mat_A[129][3] * mat_B[62][0] +
                mat_A[130][0] * mat_B[70][0] +
                mat_A[130][1] * mat_B[78][0] +
                mat_A[130][2] * mat_B[86][0] +
                mat_A[130][3] * mat_B[94][0] +
                mat_A[131][0] * mat_B[102][0] +
                mat_A[131][1] * mat_B[110][0] +
                mat_A[131][2] * mat_B[118][0] +
                mat_A[131][3] * mat_B[126][0] +
                mat_A[132][0] * mat_B[134][0] +
                mat_A[132][1] * mat_B[142][0] +
                mat_A[132][2] * mat_B[150][0] +
                mat_A[132][3] * mat_B[158][0] +
                mat_A[133][0] * mat_B[166][0] +
                mat_A[133][1] * mat_B[174][0] +
                mat_A[133][2] * mat_B[182][0] +
                mat_A[133][3] * mat_B[190][0] +
                mat_A[134][0] * mat_B[198][0] +
                mat_A[134][1] * mat_B[206][0] +
                mat_A[134][2] * mat_B[214][0] +
                mat_A[134][3] * mat_B[222][0] +
                mat_A[135][0] * mat_B[230][0] +
                mat_A[135][1] * mat_B[238][0] +
                mat_A[135][2] * mat_B[246][0] +
                mat_A[135][3] * mat_B[254][0];
    mat_C[134][1] <=
                mat_A[128][0] * mat_B[6][1] +
                mat_A[128][1] * mat_B[14][1] +
                mat_A[128][2] * mat_B[22][1] +
                mat_A[128][3] * mat_B[30][1] +
                mat_A[129][0] * mat_B[38][1] +
                mat_A[129][1] * mat_B[46][1] +
                mat_A[129][2] * mat_B[54][1] +
                mat_A[129][3] * mat_B[62][1] +
                mat_A[130][0] * mat_B[70][1] +
                mat_A[130][1] * mat_B[78][1] +
                mat_A[130][2] * mat_B[86][1] +
                mat_A[130][3] * mat_B[94][1] +
                mat_A[131][0] * mat_B[102][1] +
                mat_A[131][1] * mat_B[110][1] +
                mat_A[131][2] * mat_B[118][1] +
                mat_A[131][3] * mat_B[126][1] +
                mat_A[132][0] * mat_B[134][1] +
                mat_A[132][1] * mat_B[142][1] +
                mat_A[132][2] * mat_B[150][1] +
                mat_A[132][3] * mat_B[158][1] +
                mat_A[133][0] * mat_B[166][1] +
                mat_A[133][1] * mat_B[174][1] +
                mat_A[133][2] * mat_B[182][1] +
                mat_A[133][3] * mat_B[190][1] +
                mat_A[134][0] * mat_B[198][1] +
                mat_A[134][1] * mat_B[206][1] +
                mat_A[134][2] * mat_B[214][1] +
                mat_A[134][3] * mat_B[222][1] +
                mat_A[135][0] * mat_B[230][1] +
                mat_A[135][1] * mat_B[238][1] +
                mat_A[135][2] * mat_B[246][1] +
                mat_A[135][3] * mat_B[254][1];
    mat_C[134][2] <=
                mat_A[128][0] * mat_B[6][2] +
                mat_A[128][1] * mat_B[14][2] +
                mat_A[128][2] * mat_B[22][2] +
                mat_A[128][3] * mat_B[30][2] +
                mat_A[129][0] * mat_B[38][2] +
                mat_A[129][1] * mat_B[46][2] +
                mat_A[129][2] * mat_B[54][2] +
                mat_A[129][3] * mat_B[62][2] +
                mat_A[130][0] * mat_B[70][2] +
                mat_A[130][1] * mat_B[78][2] +
                mat_A[130][2] * mat_B[86][2] +
                mat_A[130][3] * mat_B[94][2] +
                mat_A[131][0] * mat_B[102][2] +
                mat_A[131][1] * mat_B[110][2] +
                mat_A[131][2] * mat_B[118][2] +
                mat_A[131][3] * mat_B[126][2] +
                mat_A[132][0] * mat_B[134][2] +
                mat_A[132][1] * mat_B[142][2] +
                mat_A[132][2] * mat_B[150][2] +
                mat_A[132][3] * mat_B[158][2] +
                mat_A[133][0] * mat_B[166][2] +
                mat_A[133][1] * mat_B[174][2] +
                mat_A[133][2] * mat_B[182][2] +
                mat_A[133][3] * mat_B[190][2] +
                mat_A[134][0] * mat_B[198][2] +
                mat_A[134][1] * mat_B[206][2] +
                mat_A[134][2] * mat_B[214][2] +
                mat_A[134][3] * mat_B[222][2] +
                mat_A[135][0] * mat_B[230][2] +
                mat_A[135][1] * mat_B[238][2] +
                mat_A[135][2] * mat_B[246][2] +
                mat_A[135][3] * mat_B[254][2];
    mat_C[134][3] <=
                mat_A[128][0] * mat_B[6][3] +
                mat_A[128][1] * mat_B[14][3] +
                mat_A[128][2] * mat_B[22][3] +
                mat_A[128][3] * mat_B[30][3] +
                mat_A[129][0] * mat_B[38][3] +
                mat_A[129][1] * mat_B[46][3] +
                mat_A[129][2] * mat_B[54][3] +
                mat_A[129][3] * mat_B[62][3] +
                mat_A[130][0] * mat_B[70][3] +
                mat_A[130][1] * mat_B[78][3] +
                mat_A[130][2] * mat_B[86][3] +
                mat_A[130][3] * mat_B[94][3] +
                mat_A[131][0] * mat_B[102][3] +
                mat_A[131][1] * mat_B[110][3] +
                mat_A[131][2] * mat_B[118][3] +
                mat_A[131][3] * mat_B[126][3] +
                mat_A[132][0] * mat_B[134][3] +
                mat_A[132][1] * mat_B[142][3] +
                mat_A[132][2] * mat_B[150][3] +
                mat_A[132][3] * mat_B[158][3] +
                mat_A[133][0] * mat_B[166][3] +
                mat_A[133][1] * mat_B[174][3] +
                mat_A[133][2] * mat_B[182][3] +
                mat_A[133][3] * mat_B[190][3] +
                mat_A[134][0] * mat_B[198][3] +
                mat_A[134][1] * mat_B[206][3] +
                mat_A[134][2] * mat_B[214][3] +
                mat_A[134][3] * mat_B[222][3] +
                mat_A[135][0] * mat_B[230][3] +
                mat_A[135][1] * mat_B[238][3] +
                mat_A[135][2] * mat_B[246][3] +
                mat_A[135][3] * mat_B[254][3];
    mat_C[135][0] <=
                mat_A[128][0] * mat_B[7][0] +
                mat_A[128][1] * mat_B[15][0] +
                mat_A[128][2] * mat_B[23][0] +
                mat_A[128][3] * mat_B[31][0] +
                mat_A[129][0] * mat_B[39][0] +
                mat_A[129][1] * mat_B[47][0] +
                mat_A[129][2] * mat_B[55][0] +
                mat_A[129][3] * mat_B[63][0] +
                mat_A[130][0] * mat_B[71][0] +
                mat_A[130][1] * mat_B[79][0] +
                mat_A[130][2] * mat_B[87][0] +
                mat_A[130][3] * mat_B[95][0] +
                mat_A[131][0] * mat_B[103][0] +
                mat_A[131][1] * mat_B[111][0] +
                mat_A[131][2] * mat_B[119][0] +
                mat_A[131][3] * mat_B[127][0] +
                mat_A[132][0] * mat_B[135][0] +
                mat_A[132][1] * mat_B[143][0] +
                mat_A[132][2] * mat_B[151][0] +
                mat_A[132][3] * mat_B[159][0] +
                mat_A[133][0] * mat_B[167][0] +
                mat_A[133][1] * mat_B[175][0] +
                mat_A[133][2] * mat_B[183][0] +
                mat_A[133][3] * mat_B[191][0] +
                mat_A[134][0] * mat_B[199][0] +
                mat_A[134][1] * mat_B[207][0] +
                mat_A[134][2] * mat_B[215][0] +
                mat_A[134][3] * mat_B[223][0] +
                mat_A[135][0] * mat_B[231][0] +
                mat_A[135][1] * mat_B[239][0] +
                mat_A[135][2] * mat_B[247][0] +
                mat_A[135][3] * mat_B[255][0];
    mat_C[135][1] <=
                mat_A[128][0] * mat_B[7][1] +
                mat_A[128][1] * mat_B[15][1] +
                mat_A[128][2] * mat_B[23][1] +
                mat_A[128][3] * mat_B[31][1] +
                mat_A[129][0] * mat_B[39][1] +
                mat_A[129][1] * mat_B[47][1] +
                mat_A[129][2] * mat_B[55][1] +
                mat_A[129][3] * mat_B[63][1] +
                mat_A[130][0] * mat_B[71][1] +
                mat_A[130][1] * mat_B[79][1] +
                mat_A[130][2] * mat_B[87][1] +
                mat_A[130][3] * mat_B[95][1] +
                mat_A[131][0] * mat_B[103][1] +
                mat_A[131][1] * mat_B[111][1] +
                mat_A[131][2] * mat_B[119][1] +
                mat_A[131][3] * mat_B[127][1] +
                mat_A[132][0] * mat_B[135][1] +
                mat_A[132][1] * mat_B[143][1] +
                mat_A[132][2] * mat_B[151][1] +
                mat_A[132][3] * mat_B[159][1] +
                mat_A[133][0] * mat_B[167][1] +
                mat_A[133][1] * mat_B[175][1] +
                mat_A[133][2] * mat_B[183][1] +
                mat_A[133][3] * mat_B[191][1] +
                mat_A[134][0] * mat_B[199][1] +
                mat_A[134][1] * mat_B[207][1] +
                mat_A[134][2] * mat_B[215][1] +
                mat_A[134][3] * mat_B[223][1] +
                mat_A[135][0] * mat_B[231][1] +
                mat_A[135][1] * mat_B[239][1] +
                mat_A[135][2] * mat_B[247][1] +
                mat_A[135][3] * mat_B[255][1];
    mat_C[135][2] <=
                mat_A[128][0] * mat_B[7][2] +
                mat_A[128][1] * mat_B[15][2] +
                mat_A[128][2] * mat_B[23][2] +
                mat_A[128][3] * mat_B[31][2] +
                mat_A[129][0] * mat_B[39][2] +
                mat_A[129][1] * mat_B[47][2] +
                mat_A[129][2] * mat_B[55][2] +
                mat_A[129][3] * mat_B[63][2] +
                mat_A[130][0] * mat_B[71][2] +
                mat_A[130][1] * mat_B[79][2] +
                mat_A[130][2] * mat_B[87][2] +
                mat_A[130][3] * mat_B[95][2] +
                mat_A[131][0] * mat_B[103][2] +
                mat_A[131][1] * mat_B[111][2] +
                mat_A[131][2] * mat_B[119][2] +
                mat_A[131][3] * mat_B[127][2] +
                mat_A[132][0] * mat_B[135][2] +
                mat_A[132][1] * mat_B[143][2] +
                mat_A[132][2] * mat_B[151][2] +
                mat_A[132][3] * mat_B[159][2] +
                mat_A[133][0] * mat_B[167][2] +
                mat_A[133][1] * mat_B[175][2] +
                mat_A[133][2] * mat_B[183][2] +
                mat_A[133][3] * mat_B[191][2] +
                mat_A[134][0] * mat_B[199][2] +
                mat_A[134][1] * mat_B[207][2] +
                mat_A[134][2] * mat_B[215][2] +
                mat_A[134][3] * mat_B[223][2] +
                mat_A[135][0] * mat_B[231][2] +
                mat_A[135][1] * mat_B[239][2] +
                mat_A[135][2] * mat_B[247][2] +
                mat_A[135][3] * mat_B[255][2];
    mat_C[135][3] <=
                mat_A[128][0] * mat_B[7][3] +
                mat_A[128][1] * mat_B[15][3] +
                mat_A[128][2] * mat_B[23][3] +
                mat_A[128][3] * mat_B[31][3] +
                mat_A[129][0] * mat_B[39][3] +
                mat_A[129][1] * mat_B[47][3] +
                mat_A[129][2] * mat_B[55][3] +
                mat_A[129][3] * mat_B[63][3] +
                mat_A[130][0] * mat_B[71][3] +
                mat_A[130][1] * mat_B[79][3] +
                mat_A[130][2] * mat_B[87][3] +
                mat_A[130][3] * mat_B[95][3] +
                mat_A[131][0] * mat_B[103][3] +
                mat_A[131][1] * mat_B[111][3] +
                mat_A[131][2] * mat_B[119][3] +
                mat_A[131][3] * mat_B[127][3] +
                mat_A[132][0] * mat_B[135][3] +
                mat_A[132][1] * mat_B[143][3] +
                mat_A[132][2] * mat_B[151][3] +
                mat_A[132][3] * mat_B[159][3] +
                mat_A[133][0] * mat_B[167][3] +
                mat_A[133][1] * mat_B[175][3] +
                mat_A[133][2] * mat_B[183][3] +
                mat_A[133][3] * mat_B[191][3] +
                mat_A[134][0] * mat_B[199][3] +
                mat_A[134][1] * mat_B[207][3] +
                mat_A[134][2] * mat_B[215][3] +
                mat_A[134][3] * mat_B[223][3] +
                mat_A[135][0] * mat_B[231][3] +
                mat_A[135][1] * mat_B[239][3] +
                mat_A[135][2] * mat_B[247][3] +
                mat_A[135][3] * mat_B[255][3];
    mat_C[136][0] <=
                mat_A[136][0] * mat_B[0][0] +
                mat_A[136][1] * mat_B[8][0] +
                mat_A[136][2] * mat_B[16][0] +
                mat_A[136][3] * mat_B[24][0] +
                mat_A[137][0] * mat_B[32][0] +
                mat_A[137][1] * mat_B[40][0] +
                mat_A[137][2] * mat_B[48][0] +
                mat_A[137][3] * mat_B[56][0] +
                mat_A[138][0] * mat_B[64][0] +
                mat_A[138][1] * mat_B[72][0] +
                mat_A[138][2] * mat_B[80][0] +
                mat_A[138][3] * mat_B[88][0] +
                mat_A[139][0] * mat_B[96][0] +
                mat_A[139][1] * mat_B[104][0] +
                mat_A[139][2] * mat_B[112][0] +
                mat_A[139][3] * mat_B[120][0] +
                mat_A[140][0] * mat_B[128][0] +
                mat_A[140][1] * mat_B[136][0] +
                mat_A[140][2] * mat_B[144][0] +
                mat_A[140][3] * mat_B[152][0] +
                mat_A[141][0] * mat_B[160][0] +
                mat_A[141][1] * mat_B[168][0] +
                mat_A[141][2] * mat_B[176][0] +
                mat_A[141][3] * mat_B[184][0] +
                mat_A[142][0] * mat_B[192][0] +
                mat_A[142][1] * mat_B[200][0] +
                mat_A[142][2] * mat_B[208][0] +
                mat_A[142][3] * mat_B[216][0] +
                mat_A[143][0] * mat_B[224][0] +
                mat_A[143][1] * mat_B[232][0] +
                mat_A[143][2] * mat_B[240][0] +
                mat_A[143][3] * mat_B[248][0];
    mat_C[136][1] <=
                mat_A[136][0] * mat_B[0][1] +
                mat_A[136][1] * mat_B[8][1] +
                mat_A[136][2] * mat_B[16][1] +
                mat_A[136][3] * mat_B[24][1] +
                mat_A[137][0] * mat_B[32][1] +
                mat_A[137][1] * mat_B[40][1] +
                mat_A[137][2] * mat_B[48][1] +
                mat_A[137][3] * mat_B[56][1] +
                mat_A[138][0] * mat_B[64][1] +
                mat_A[138][1] * mat_B[72][1] +
                mat_A[138][2] * mat_B[80][1] +
                mat_A[138][3] * mat_B[88][1] +
                mat_A[139][0] * mat_B[96][1] +
                mat_A[139][1] * mat_B[104][1] +
                mat_A[139][2] * mat_B[112][1] +
                mat_A[139][3] * mat_B[120][1] +
                mat_A[140][0] * mat_B[128][1] +
                mat_A[140][1] * mat_B[136][1] +
                mat_A[140][2] * mat_B[144][1] +
                mat_A[140][3] * mat_B[152][1] +
                mat_A[141][0] * mat_B[160][1] +
                mat_A[141][1] * mat_B[168][1] +
                mat_A[141][2] * mat_B[176][1] +
                mat_A[141][3] * mat_B[184][1] +
                mat_A[142][0] * mat_B[192][1] +
                mat_A[142][1] * mat_B[200][1] +
                mat_A[142][2] * mat_B[208][1] +
                mat_A[142][3] * mat_B[216][1] +
                mat_A[143][0] * mat_B[224][1] +
                mat_A[143][1] * mat_B[232][1] +
                mat_A[143][2] * mat_B[240][1] +
                mat_A[143][3] * mat_B[248][1];
    mat_C[136][2] <=
                mat_A[136][0] * mat_B[0][2] +
                mat_A[136][1] * mat_B[8][2] +
                mat_A[136][2] * mat_B[16][2] +
                mat_A[136][3] * mat_B[24][2] +
                mat_A[137][0] * mat_B[32][2] +
                mat_A[137][1] * mat_B[40][2] +
                mat_A[137][2] * mat_B[48][2] +
                mat_A[137][3] * mat_B[56][2] +
                mat_A[138][0] * mat_B[64][2] +
                mat_A[138][1] * mat_B[72][2] +
                mat_A[138][2] * mat_B[80][2] +
                mat_A[138][3] * mat_B[88][2] +
                mat_A[139][0] * mat_B[96][2] +
                mat_A[139][1] * mat_B[104][2] +
                mat_A[139][2] * mat_B[112][2] +
                mat_A[139][3] * mat_B[120][2] +
                mat_A[140][0] * mat_B[128][2] +
                mat_A[140][1] * mat_B[136][2] +
                mat_A[140][2] * mat_B[144][2] +
                mat_A[140][3] * mat_B[152][2] +
                mat_A[141][0] * mat_B[160][2] +
                mat_A[141][1] * mat_B[168][2] +
                mat_A[141][2] * mat_B[176][2] +
                mat_A[141][3] * mat_B[184][2] +
                mat_A[142][0] * mat_B[192][2] +
                mat_A[142][1] * mat_B[200][2] +
                mat_A[142][2] * mat_B[208][2] +
                mat_A[142][3] * mat_B[216][2] +
                mat_A[143][0] * mat_B[224][2] +
                mat_A[143][1] * mat_B[232][2] +
                mat_A[143][2] * mat_B[240][2] +
                mat_A[143][3] * mat_B[248][2];
    mat_C[136][3] <=
                mat_A[136][0] * mat_B[0][3] +
                mat_A[136][1] * mat_B[8][3] +
                mat_A[136][2] * mat_B[16][3] +
                mat_A[136][3] * mat_B[24][3] +
                mat_A[137][0] * mat_B[32][3] +
                mat_A[137][1] * mat_B[40][3] +
                mat_A[137][2] * mat_B[48][3] +
                mat_A[137][3] * mat_B[56][3] +
                mat_A[138][0] * mat_B[64][3] +
                mat_A[138][1] * mat_B[72][3] +
                mat_A[138][2] * mat_B[80][3] +
                mat_A[138][3] * mat_B[88][3] +
                mat_A[139][0] * mat_B[96][3] +
                mat_A[139][1] * mat_B[104][3] +
                mat_A[139][2] * mat_B[112][3] +
                mat_A[139][3] * mat_B[120][3] +
                mat_A[140][0] * mat_B[128][3] +
                mat_A[140][1] * mat_B[136][3] +
                mat_A[140][2] * mat_B[144][3] +
                mat_A[140][3] * mat_B[152][3] +
                mat_A[141][0] * mat_B[160][3] +
                mat_A[141][1] * mat_B[168][3] +
                mat_A[141][2] * mat_B[176][3] +
                mat_A[141][3] * mat_B[184][3] +
                mat_A[142][0] * mat_B[192][3] +
                mat_A[142][1] * mat_B[200][3] +
                mat_A[142][2] * mat_B[208][3] +
                mat_A[142][3] * mat_B[216][3] +
                mat_A[143][0] * mat_B[224][3] +
                mat_A[143][1] * mat_B[232][3] +
                mat_A[143][2] * mat_B[240][3] +
                mat_A[143][3] * mat_B[248][3];
    mat_C[137][0] <=
                mat_A[136][0] * mat_B[1][0] +
                mat_A[136][1] * mat_B[9][0] +
                mat_A[136][2] * mat_B[17][0] +
                mat_A[136][3] * mat_B[25][0] +
                mat_A[137][0] * mat_B[33][0] +
                mat_A[137][1] * mat_B[41][0] +
                mat_A[137][2] * mat_B[49][0] +
                mat_A[137][3] * mat_B[57][0] +
                mat_A[138][0] * mat_B[65][0] +
                mat_A[138][1] * mat_B[73][0] +
                mat_A[138][2] * mat_B[81][0] +
                mat_A[138][3] * mat_B[89][0] +
                mat_A[139][0] * mat_B[97][0] +
                mat_A[139][1] * mat_B[105][0] +
                mat_A[139][2] * mat_B[113][0] +
                mat_A[139][3] * mat_B[121][0] +
                mat_A[140][0] * mat_B[129][0] +
                mat_A[140][1] * mat_B[137][0] +
                mat_A[140][2] * mat_B[145][0] +
                mat_A[140][3] * mat_B[153][0] +
                mat_A[141][0] * mat_B[161][0] +
                mat_A[141][1] * mat_B[169][0] +
                mat_A[141][2] * mat_B[177][0] +
                mat_A[141][3] * mat_B[185][0] +
                mat_A[142][0] * mat_B[193][0] +
                mat_A[142][1] * mat_B[201][0] +
                mat_A[142][2] * mat_B[209][0] +
                mat_A[142][3] * mat_B[217][0] +
                mat_A[143][0] * mat_B[225][0] +
                mat_A[143][1] * mat_B[233][0] +
                mat_A[143][2] * mat_B[241][0] +
                mat_A[143][3] * mat_B[249][0];
    mat_C[137][1] <=
                mat_A[136][0] * mat_B[1][1] +
                mat_A[136][1] * mat_B[9][1] +
                mat_A[136][2] * mat_B[17][1] +
                mat_A[136][3] * mat_B[25][1] +
                mat_A[137][0] * mat_B[33][1] +
                mat_A[137][1] * mat_B[41][1] +
                mat_A[137][2] * mat_B[49][1] +
                mat_A[137][3] * mat_B[57][1] +
                mat_A[138][0] * mat_B[65][1] +
                mat_A[138][1] * mat_B[73][1] +
                mat_A[138][2] * mat_B[81][1] +
                mat_A[138][3] * mat_B[89][1] +
                mat_A[139][0] * mat_B[97][1] +
                mat_A[139][1] * mat_B[105][1] +
                mat_A[139][2] * mat_B[113][1] +
                mat_A[139][3] * mat_B[121][1] +
                mat_A[140][0] * mat_B[129][1] +
                mat_A[140][1] * mat_B[137][1] +
                mat_A[140][2] * mat_B[145][1] +
                mat_A[140][3] * mat_B[153][1] +
                mat_A[141][0] * mat_B[161][1] +
                mat_A[141][1] * mat_B[169][1] +
                mat_A[141][2] * mat_B[177][1] +
                mat_A[141][3] * mat_B[185][1] +
                mat_A[142][0] * mat_B[193][1] +
                mat_A[142][1] * mat_B[201][1] +
                mat_A[142][2] * mat_B[209][1] +
                mat_A[142][3] * mat_B[217][1] +
                mat_A[143][0] * mat_B[225][1] +
                mat_A[143][1] * mat_B[233][1] +
                mat_A[143][2] * mat_B[241][1] +
                mat_A[143][3] * mat_B[249][1];
    mat_C[137][2] <=
                mat_A[136][0] * mat_B[1][2] +
                mat_A[136][1] * mat_B[9][2] +
                mat_A[136][2] * mat_B[17][2] +
                mat_A[136][3] * mat_B[25][2] +
                mat_A[137][0] * mat_B[33][2] +
                mat_A[137][1] * mat_B[41][2] +
                mat_A[137][2] * mat_B[49][2] +
                mat_A[137][3] * mat_B[57][2] +
                mat_A[138][0] * mat_B[65][2] +
                mat_A[138][1] * mat_B[73][2] +
                mat_A[138][2] * mat_B[81][2] +
                mat_A[138][3] * mat_B[89][2] +
                mat_A[139][0] * mat_B[97][2] +
                mat_A[139][1] * mat_B[105][2] +
                mat_A[139][2] * mat_B[113][2] +
                mat_A[139][3] * mat_B[121][2] +
                mat_A[140][0] * mat_B[129][2] +
                mat_A[140][1] * mat_B[137][2] +
                mat_A[140][2] * mat_B[145][2] +
                mat_A[140][3] * mat_B[153][2] +
                mat_A[141][0] * mat_B[161][2] +
                mat_A[141][1] * mat_B[169][2] +
                mat_A[141][2] * mat_B[177][2] +
                mat_A[141][3] * mat_B[185][2] +
                mat_A[142][0] * mat_B[193][2] +
                mat_A[142][1] * mat_B[201][2] +
                mat_A[142][2] * mat_B[209][2] +
                mat_A[142][3] * mat_B[217][2] +
                mat_A[143][0] * mat_B[225][2] +
                mat_A[143][1] * mat_B[233][2] +
                mat_A[143][2] * mat_B[241][2] +
                mat_A[143][3] * mat_B[249][2];
    mat_C[137][3] <=
                mat_A[136][0] * mat_B[1][3] +
                mat_A[136][1] * mat_B[9][3] +
                mat_A[136][2] * mat_B[17][3] +
                mat_A[136][3] * mat_B[25][3] +
                mat_A[137][0] * mat_B[33][3] +
                mat_A[137][1] * mat_B[41][3] +
                mat_A[137][2] * mat_B[49][3] +
                mat_A[137][3] * mat_B[57][3] +
                mat_A[138][0] * mat_B[65][3] +
                mat_A[138][1] * mat_B[73][3] +
                mat_A[138][2] * mat_B[81][3] +
                mat_A[138][3] * mat_B[89][3] +
                mat_A[139][0] * mat_B[97][3] +
                mat_A[139][1] * mat_B[105][3] +
                mat_A[139][2] * mat_B[113][3] +
                mat_A[139][3] * mat_B[121][3] +
                mat_A[140][0] * mat_B[129][3] +
                mat_A[140][1] * mat_B[137][3] +
                mat_A[140][2] * mat_B[145][3] +
                mat_A[140][3] * mat_B[153][3] +
                mat_A[141][0] * mat_B[161][3] +
                mat_A[141][1] * mat_B[169][3] +
                mat_A[141][2] * mat_B[177][3] +
                mat_A[141][3] * mat_B[185][3] +
                mat_A[142][0] * mat_B[193][3] +
                mat_A[142][1] * mat_B[201][3] +
                mat_A[142][2] * mat_B[209][3] +
                mat_A[142][3] * mat_B[217][3] +
                mat_A[143][0] * mat_B[225][3] +
                mat_A[143][1] * mat_B[233][3] +
                mat_A[143][2] * mat_B[241][3] +
                mat_A[143][3] * mat_B[249][3];
    mat_C[138][0] <=
                mat_A[136][0] * mat_B[2][0] +
                mat_A[136][1] * mat_B[10][0] +
                mat_A[136][2] * mat_B[18][0] +
                mat_A[136][3] * mat_B[26][0] +
                mat_A[137][0] * mat_B[34][0] +
                mat_A[137][1] * mat_B[42][0] +
                mat_A[137][2] * mat_B[50][0] +
                mat_A[137][3] * mat_B[58][0] +
                mat_A[138][0] * mat_B[66][0] +
                mat_A[138][1] * mat_B[74][0] +
                mat_A[138][2] * mat_B[82][0] +
                mat_A[138][3] * mat_B[90][0] +
                mat_A[139][0] * mat_B[98][0] +
                mat_A[139][1] * mat_B[106][0] +
                mat_A[139][2] * mat_B[114][0] +
                mat_A[139][3] * mat_B[122][0] +
                mat_A[140][0] * mat_B[130][0] +
                mat_A[140][1] * mat_B[138][0] +
                mat_A[140][2] * mat_B[146][0] +
                mat_A[140][3] * mat_B[154][0] +
                mat_A[141][0] * mat_B[162][0] +
                mat_A[141][1] * mat_B[170][0] +
                mat_A[141][2] * mat_B[178][0] +
                mat_A[141][3] * mat_B[186][0] +
                mat_A[142][0] * mat_B[194][0] +
                mat_A[142][1] * mat_B[202][0] +
                mat_A[142][2] * mat_B[210][0] +
                mat_A[142][3] * mat_B[218][0] +
                mat_A[143][0] * mat_B[226][0] +
                mat_A[143][1] * mat_B[234][0] +
                mat_A[143][2] * mat_B[242][0] +
                mat_A[143][3] * mat_B[250][0];
    mat_C[138][1] <=
                mat_A[136][0] * mat_B[2][1] +
                mat_A[136][1] * mat_B[10][1] +
                mat_A[136][2] * mat_B[18][1] +
                mat_A[136][3] * mat_B[26][1] +
                mat_A[137][0] * mat_B[34][1] +
                mat_A[137][1] * mat_B[42][1] +
                mat_A[137][2] * mat_B[50][1] +
                mat_A[137][3] * mat_B[58][1] +
                mat_A[138][0] * mat_B[66][1] +
                mat_A[138][1] * mat_B[74][1] +
                mat_A[138][2] * mat_B[82][1] +
                mat_A[138][3] * mat_B[90][1] +
                mat_A[139][0] * mat_B[98][1] +
                mat_A[139][1] * mat_B[106][1] +
                mat_A[139][2] * mat_B[114][1] +
                mat_A[139][3] * mat_B[122][1] +
                mat_A[140][0] * mat_B[130][1] +
                mat_A[140][1] * mat_B[138][1] +
                mat_A[140][2] * mat_B[146][1] +
                mat_A[140][3] * mat_B[154][1] +
                mat_A[141][0] * mat_B[162][1] +
                mat_A[141][1] * mat_B[170][1] +
                mat_A[141][2] * mat_B[178][1] +
                mat_A[141][3] * mat_B[186][1] +
                mat_A[142][0] * mat_B[194][1] +
                mat_A[142][1] * mat_B[202][1] +
                mat_A[142][2] * mat_B[210][1] +
                mat_A[142][3] * mat_B[218][1] +
                mat_A[143][0] * mat_B[226][1] +
                mat_A[143][1] * mat_B[234][1] +
                mat_A[143][2] * mat_B[242][1] +
                mat_A[143][3] * mat_B[250][1];
    mat_C[138][2] <=
                mat_A[136][0] * mat_B[2][2] +
                mat_A[136][1] * mat_B[10][2] +
                mat_A[136][2] * mat_B[18][2] +
                mat_A[136][3] * mat_B[26][2] +
                mat_A[137][0] * mat_B[34][2] +
                mat_A[137][1] * mat_B[42][2] +
                mat_A[137][2] * mat_B[50][2] +
                mat_A[137][3] * mat_B[58][2] +
                mat_A[138][0] * mat_B[66][2] +
                mat_A[138][1] * mat_B[74][2] +
                mat_A[138][2] * mat_B[82][2] +
                mat_A[138][3] * mat_B[90][2] +
                mat_A[139][0] * mat_B[98][2] +
                mat_A[139][1] * mat_B[106][2] +
                mat_A[139][2] * mat_B[114][2] +
                mat_A[139][3] * mat_B[122][2] +
                mat_A[140][0] * mat_B[130][2] +
                mat_A[140][1] * mat_B[138][2] +
                mat_A[140][2] * mat_B[146][2] +
                mat_A[140][3] * mat_B[154][2] +
                mat_A[141][0] * mat_B[162][2] +
                mat_A[141][1] * mat_B[170][2] +
                mat_A[141][2] * mat_B[178][2] +
                mat_A[141][3] * mat_B[186][2] +
                mat_A[142][0] * mat_B[194][2] +
                mat_A[142][1] * mat_B[202][2] +
                mat_A[142][2] * mat_B[210][2] +
                mat_A[142][3] * mat_B[218][2] +
                mat_A[143][0] * mat_B[226][2] +
                mat_A[143][1] * mat_B[234][2] +
                mat_A[143][2] * mat_B[242][2] +
                mat_A[143][3] * mat_B[250][2];
    mat_C[138][3] <=
                mat_A[136][0] * mat_B[2][3] +
                mat_A[136][1] * mat_B[10][3] +
                mat_A[136][2] * mat_B[18][3] +
                mat_A[136][3] * mat_B[26][3] +
                mat_A[137][0] * mat_B[34][3] +
                mat_A[137][1] * mat_B[42][3] +
                mat_A[137][2] * mat_B[50][3] +
                mat_A[137][3] * mat_B[58][3] +
                mat_A[138][0] * mat_B[66][3] +
                mat_A[138][1] * mat_B[74][3] +
                mat_A[138][2] * mat_B[82][3] +
                mat_A[138][3] * mat_B[90][3] +
                mat_A[139][0] * mat_B[98][3] +
                mat_A[139][1] * mat_B[106][3] +
                mat_A[139][2] * mat_B[114][3] +
                mat_A[139][3] * mat_B[122][3] +
                mat_A[140][0] * mat_B[130][3] +
                mat_A[140][1] * mat_B[138][3] +
                mat_A[140][2] * mat_B[146][3] +
                mat_A[140][3] * mat_B[154][3] +
                mat_A[141][0] * mat_B[162][3] +
                mat_A[141][1] * mat_B[170][3] +
                mat_A[141][2] * mat_B[178][3] +
                mat_A[141][3] * mat_B[186][3] +
                mat_A[142][0] * mat_B[194][3] +
                mat_A[142][1] * mat_B[202][3] +
                mat_A[142][2] * mat_B[210][3] +
                mat_A[142][3] * mat_B[218][3] +
                mat_A[143][0] * mat_B[226][3] +
                mat_A[143][1] * mat_B[234][3] +
                mat_A[143][2] * mat_B[242][3] +
                mat_A[143][3] * mat_B[250][3];
    mat_C[139][0] <=
                mat_A[136][0] * mat_B[3][0] +
                mat_A[136][1] * mat_B[11][0] +
                mat_A[136][2] * mat_B[19][0] +
                mat_A[136][3] * mat_B[27][0] +
                mat_A[137][0] * mat_B[35][0] +
                mat_A[137][1] * mat_B[43][0] +
                mat_A[137][2] * mat_B[51][0] +
                mat_A[137][3] * mat_B[59][0] +
                mat_A[138][0] * mat_B[67][0] +
                mat_A[138][1] * mat_B[75][0] +
                mat_A[138][2] * mat_B[83][0] +
                mat_A[138][3] * mat_B[91][0] +
                mat_A[139][0] * mat_B[99][0] +
                mat_A[139][1] * mat_B[107][0] +
                mat_A[139][2] * mat_B[115][0] +
                mat_A[139][3] * mat_B[123][0] +
                mat_A[140][0] * mat_B[131][0] +
                mat_A[140][1] * mat_B[139][0] +
                mat_A[140][2] * mat_B[147][0] +
                mat_A[140][3] * mat_B[155][0] +
                mat_A[141][0] * mat_B[163][0] +
                mat_A[141][1] * mat_B[171][0] +
                mat_A[141][2] * mat_B[179][0] +
                mat_A[141][3] * mat_B[187][0] +
                mat_A[142][0] * mat_B[195][0] +
                mat_A[142][1] * mat_B[203][0] +
                mat_A[142][2] * mat_B[211][0] +
                mat_A[142][3] * mat_B[219][0] +
                mat_A[143][0] * mat_B[227][0] +
                mat_A[143][1] * mat_B[235][0] +
                mat_A[143][2] * mat_B[243][0] +
                mat_A[143][3] * mat_B[251][0];
    mat_C[139][1] <=
                mat_A[136][0] * mat_B[3][1] +
                mat_A[136][1] * mat_B[11][1] +
                mat_A[136][2] * mat_B[19][1] +
                mat_A[136][3] * mat_B[27][1] +
                mat_A[137][0] * mat_B[35][1] +
                mat_A[137][1] * mat_B[43][1] +
                mat_A[137][2] * mat_B[51][1] +
                mat_A[137][3] * mat_B[59][1] +
                mat_A[138][0] * mat_B[67][1] +
                mat_A[138][1] * mat_B[75][1] +
                mat_A[138][2] * mat_B[83][1] +
                mat_A[138][3] * mat_B[91][1] +
                mat_A[139][0] * mat_B[99][1] +
                mat_A[139][1] * mat_B[107][1] +
                mat_A[139][2] * mat_B[115][1] +
                mat_A[139][3] * mat_B[123][1] +
                mat_A[140][0] * mat_B[131][1] +
                mat_A[140][1] * mat_B[139][1] +
                mat_A[140][2] * mat_B[147][1] +
                mat_A[140][3] * mat_B[155][1] +
                mat_A[141][0] * mat_B[163][1] +
                mat_A[141][1] * mat_B[171][1] +
                mat_A[141][2] * mat_B[179][1] +
                mat_A[141][3] * mat_B[187][1] +
                mat_A[142][0] * mat_B[195][1] +
                mat_A[142][1] * mat_B[203][1] +
                mat_A[142][2] * mat_B[211][1] +
                mat_A[142][3] * mat_B[219][1] +
                mat_A[143][0] * mat_B[227][1] +
                mat_A[143][1] * mat_B[235][1] +
                mat_A[143][2] * mat_B[243][1] +
                mat_A[143][3] * mat_B[251][1];
    mat_C[139][2] <=
                mat_A[136][0] * mat_B[3][2] +
                mat_A[136][1] * mat_B[11][2] +
                mat_A[136][2] * mat_B[19][2] +
                mat_A[136][3] * mat_B[27][2] +
                mat_A[137][0] * mat_B[35][2] +
                mat_A[137][1] * mat_B[43][2] +
                mat_A[137][2] * mat_B[51][2] +
                mat_A[137][3] * mat_B[59][2] +
                mat_A[138][0] * mat_B[67][2] +
                mat_A[138][1] * mat_B[75][2] +
                mat_A[138][2] * mat_B[83][2] +
                mat_A[138][3] * mat_B[91][2] +
                mat_A[139][0] * mat_B[99][2] +
                mat_A[139][1] * mat_B[107][2] +
                mat_A[139][2] * mat_B[115][2] +
                mat_A[139][3] * mat_B[123][2] +
                mat_A[140][0] * mat_B[131][2] +
                mat_A[140][1] * mat_B[139][2] +
                mat_A[140][2] * mat_B[147][2] +
                mat_A[140][3] * mat_B[155][2] +
                mat_A[141][0] * mat_B[163][2] +
                mat_A[141][1] * mat_B[171][2] +
                mat_A[141][2] * mat_B[179][2] +
                mat_A[141][3] * mat_B[187][2] +
                mat_A[142][0] * mat_B[195][2] +
                mat_A[142][1] * mat_B[203][2] +
                mat_A[142][2] * mat_B[211][2] +
                mat_A[142][3] * mat_B[219][2] +
                mat_A[143][0] * mat_B[227][2] +
                mat_A[143][1] * mat_B[235][2] +
                mat_A[143][2] * mat_B[243][2] +
                mat_A[143][3] * mat_B[251][2];
    mat_C[139][3] <=
                mat_A[136][0] * mat_B[3][3] +
                mat_A[136][1] * mat_B[11][3] +
                mat_A[136][2] * mat_B[19][3] +
                mat_A[136][3] * mat_B[27][3] +
                mat_A[137][0] * mat_B[35][3] +
                mat_A[137][1] * mat_B[43][3] +
                mat_A[137][2] * mat_B[51][3] +
                mat_A[137][3] * mat_B[59][3] +
                mat_A[138][0] * mat_B[67][3] +
                mat_A[138][1] * mat_B[75][3] +
                mat_A[138][2] * mat_B[83][3] +
                mat_A[138][3] * mat_B[91][3] +
                mat_A[139][0] * mat_B[99][3] +
                mat_A[139][1] * mat_B[107][3] +
                mat_A[139][2] * mat_B[115][3] +
                mat_A[139][3] * mat_B[123][3] +
                mat_A[140][0] * mat_B[131][3] +
                mat_A[140][1] * mat_B[139][3] +
                mat_A[140][2] * mat_B[147][3] +
                mat_A[140][3] * mat_B[155][3] +
                mat_A[141][0] * mat_B[163][3] +
                mat_A[141][1] * mat_B[171][3] +
                mat_A[141][2] * mat_B[179][3] +
                mat_A[141][3] * mat_B[187][3] +
                mat_A[142][0] * mat_B[195][3] +
                mat_A[142][1] * mat_B[203][3] +
                mat_A[142][2] * mat_B[211][3] +
                mat_A[142][3] * mat_B[219][3] +
                mat_A[143][0] * mat_B[227][3] +
                mat_A[143][1] * mat_B[235][3] +
                mat_A[143][2] * mat_B[243][3] +
                mat_A[143][3] * mat_B[251][3];
    mat_C[140][0] <=
                mat_A[136][0] * mat_B[4][0] +
                mat_A[136][1] * mat_B[12][0] +
                mat_A[136][2] * mat_B[20][0] +
                mat_A[136][3] * mat_B[28][0] +
                mat_A[137][0] * mat_B[36][0] +
                mat_A[137][1] * mat_B[44][0] +
                mat_A[137][2] * mat_B[52][0] +
                mat_A[137][3] * mat_B[60][0] +
                mat_A[138][0] * mat_B[68][0] +
                mat_A[138][1] * mat_B[76][0] +
                mat_A[138][2] * mat_B[84][0] +
                mat_A[138][3] * mat_B[92][0] +
                mat_A[139][0] * mat_B[100][0] +
                mat_A[139][1] * mat_B[108][0] +
                mat_A[139][2] * mat_B[116][0] +
                mat_A[139][3] * mat_B[124][0] +
                mat_A[140][0] * mat_B[132][0] +
                mat_A[140][1] * mat_B[140][0] +
                mat_A[140][2] * mat_B[148][0] +
                mat_A[140][3] * mat_B[156][0] +
                mat_A[141][0] * mat_B[164][0] +
                mat_A[141][1] * mat_B[172][0] +
                mat_A[141][2] * mat_B[180][0] +
                mat_A[141][3] * mat_B[188][0] +
                mat_A[142][0] * mat_B[196][0] +
                mat_A[142][1] * mat_B[204][0] +
                mat_A[142][2] * mat_B[212][0] +
                mat_A[142][3] * mat_B[220][0] +
                mat_A[143][0] * mat_B[228][0] +
                mat_A[143][1] * mat_B[236][0] +
                mat_A[143][2] * mat_B[244][0] +
                mat_A[143][3] * mat_B[252][0];
    mat_C[140][1] <=
                mat_A[136][0] * mat_B[4][1] +
                mat_A[136][1] * mat_B[12][1] +
                mat_A[136][2] * mat_B[20][1] +
                mat_A[136][3] * mat_B[28][1] +
                mat_A[137][0] * mat_B[36][1] +
                mat_A[137][1] * mat_B[44][1] +
                mat_A[137][2] * mat_B[52][1] +
                mat_A[137][3] * mat_B[60][1] +
                mat_A[138][0] * mat_B[68][1] +
                mat_A[138][1] * mat_B[76][1] +
                mat_A[138][2] * mat_B[84][1] +
                mat_A[138][3] * mat_B[92][1] +
                mat_A[139][0] * mat_B[100][1] +
                mat_A[139][1] * mat_B[108][1] +
                mat_A[139][2] * mat_B[116][1] +
                mat_A[139][3] * mat_B[124][1] +
                mat_A[140][0] * mat_B[132][1] +
                mat_A[140][1] * mat_B[140][1] +
                mat_A[140][2] * mat_B[148][1] +
                mat_A[140][3] * mat_B[156][1] +
                mat_A[141][0] * mat_B[164][1] +
                mat_A[141][1] * mat_B[172][1] +
                mat_A[141][2] * mat_B[180][1] +
                mat_A[141][3] * mat_B[188][1] +
                mat_A[142][0] * mat_B[196][1] +
                mat_A[142][1] * mat_B[204][1] +
                mat_A[142][2] * mat_B[212][1] +
                mat_A[142][3] * mat_B[220][1] +
                mat_A[143][0] * mat_B[228][1] +
                mat_A[143][1] * mat_B[236][1] +
                mat_A[143][2] * mat_B[244][1] +
                mat_A[143][3] * mat_B[252][1];
    mat_C[140][2] <=
                mat_A[136][0] * mat_B[4][2] +
                mat_A[136][1] * mat_B[12][2] +
                mat_A[136][2] * mat_B[20][2] +
                mat_A[136][3] * mat_B[28][2] +
                mat_A[137][0] * mat_B[36][2] +
                mat_A[137][1] * mat_B[44][2] +
                mat_A[137][2] * mat_B[52][2] +
                mat_A[137][3] * mat_B[60][2] +
                mat_A[138][0] * mat_B[68][2] +
                mat_A[138][1] * mat_B[76][2] +
                mat_A[138][2] * mat_B[84][2] +
                mat_A[138][3] * mat_B[92][2] +
                mat_A[139][0] * mat_B[100][2] +
                mat_A[139][1] * mat_B[108][2] +
                mat_A[139][2] * mat_B[116][2] +
                mat_A[139][3] * mat_B[124][2] +
                mat_A[140][0] * mat_B[132][2] +
                mat_A[140][1] * mat_B[140][2] +
                mat_A[140][2] * mat_B[148][2] +
                mat_A[140][3] * mat_B[156][2] +
                mat_A[141][0] * mat_B[164][2] +
                mat_A[141][1] * mat_B[172][2] +
                mat_A[141][2] * mat_B[180][2] +
                mat_A[141][3] * mat_B[188][2] +
                mat_A[142][0] * mat_B[196][2] +
                mat_A[142][1] * mat_B[204][2] +
                mat_A[142][2] * mat_B[212][2] +
                mat_A[142][3] * mat_B[220][2] +
                mat_A[143][0] * mat_B[228][2] +
                mat_A[143][1] * mat_B[236][2] +
                mat_A[143][2] * mat_B[244][2] +
                mat_A[143][3] * mat_B[252][2];
    mat_C[140][3] <=
                mat_A[136][0] * mat_B[4][3] +
                mat_A[136][1] * mat_B[12][3] +
                mat_A[136][2] * mat_B[20][3] +
                mat_A[136][3] * mat_B[28][3] +
                mat_A[137][0] * mat_B[36][3] +
                mat_A[137][1] * mat_B[44][3] +
                mat_A[137][2] * mat_B[52][3] +
                mat_A[137][3] * mat_B[60][3] +
                mat_A[138][0] * mat_B[68][3] +
                mat_A[138][1] * mat_B[76][3] +
                mat_A[138][2] * mat_B[84][3] +
                mat_A[138][3] * mat_B[92][3] +
                mat_A[139][0] * mat_B[100][3] +
                mat_A[139][1] * mat_B[108][3] +
                mat_A[139][2] * mat_B[116][3] +
                mat_A[139][3] * mat_B[124][3] +
                mat_A[140][0] * mat_B[132][3] +
                mat_A[140][1] * mat_B[140][3] +
                mat_A[140][2] * mat_B[148][3] +
                mat_A[140][3] * mat_B[156][3] +
                mat_A[141][0] * mat_B[164][3] +
                mat_A[141][1] * mat_B[172][3] +
                mat_A[141][2] * mat_B[180][3] +
                mat_A[141][3] * mat_B[188][3] +
                mat_A[142][0] * mat_B[196][3] +
                mat_A[142][1] * mat_B[204][3] +
                mat_A[142][2] * mat_B[212][3] +
                mat_A[142][3] * mat_B[220][3] +
                mat_A[143][0] * mat_B[228][3] +
                mat_A[143][1] * mat_B[236][3] +
                mat_A[143][2] * mat_B[244][3] +
                mat_A[143][3] * mat_B[252][3];
    mat_C[141][0] <=
                mat_A[136][0] * mat_B[5][0] +
                mat_A[136][1] * mat_B[13][0] +
                mat_A[136][2] * mat_B[21][0] +
                mat_A[136][3] * mat_B[29][0] +
                mat_A[137][0] * mat_B[37][0] +
                mat_A[137][1] * mat_B[45][0] +
                mat_A[137][2] * mat_B[53][0] +
                mat_A[137][3] * mat_B[61][0] +
                mat_A[138][0] * mat_B[69][0] +
                mat_A[138][1] * mat_B[77][0] +
                mat_A[138][2] * mat_B[85][0] +
                mat_A[138][3] * mat_B[93][0] +
                mat_A[139][0] * mat_B[101][0] +
                mat_A[139][1] * mat_B[109][0] +
                mat_A[139][2] * mat_B[117][0] +
                mat_A[139][3] * mat_B[125][0] +
                mat_A[140][0] * mat_B[133][0] +
                mat_A[140][1] * mat_B[141][0] +
                mat_A[140][2] * mat_B[149][0] +
                mat_A[140][3] * mat_B[157][0] +
                mat_A[141][0] * mat_B[165][0] +
                mat_A[141][1] * mat_B[173][0] +
                mat_A[141][2] * mat_B[181][0] +
                mat_A[141][3] * mat_B[189][0] +
                mat_A[142][0] * mat_B[197][0] +
                mat_A[142][1] * mat_B[205][0] +
                mat_A[142][2] * mat_B[213][0] +
                mat_A[142][3] * mat_B[221][0] +
                mat_A[143][0] * mat_B[229][0] +
                mat_A[143][1] * mat_B[237][0] +
                mat_A[143][2] * mat_B[245][0] +
                mat_A[143][3] * mat_B[253][0];
    mat_C[141][1] <=
                mat_A[136][0] * mat_B[5][1] +
                mat_A[136][1] * mat_B[13][1] +
                mat_A[136][2] * mat_B[21][1] +
                mat_A[136][3] * mat_B[29][1] +
                mat_A[137][0] * mat_B[37][1] +
                mat_A[137][1] * mat_B[45][1] +
                mat_A[137][2] * mat_B[53][1] +
                mat_A[137][3] * mat_B[61][1] +
                mat_A[138][0] * mat_B[69][1] +
                mat_A[138][1] * mat_B[77][1] +
                mat_A[138][2] * mat_B[85][1] +
                mat_A[138][3] * mat_B[93][1] +
                mat_A[139][0] * mat_B[101][1] +
                mat_A[139][1] * mat_B[109][1] +
                mat_A[139][2] * mat_B[117][1] +
                mat_A[139][3] * mat_B[125][1] +
                mat_A[140][0] * mat_B[133][1] +
                mat_A[140][1] * mat_B[141][1] +
                mat_A[140][2] * mat_B[149][1] +
                mat_A[140][3] * mat_B[157][1] +
                mat_A[141][0] * mat_B[165][1] +
                mat_A[141][1] * mat_B[173][1] +
                mat_A[141][2] * mat_B[181][1] +
                mat_A[141][3] * mat_B[189][1] +
                mat_A[142][0] * mat_B[197][1] +
                mat_A[142][1] * mat_B[205][1] +
                mat_A[142][2] * mat_B[213][1] +
                mat_A[142][3] * mat_B[221][1] +
                mat_A[143][0] * mat_B[229][1] +
                mat_A[143][1] * mat_B[237][1] +
                mat_A[143][2] * mat_B[245][1] +
                mat_A[143][3] * mat_B[253][1];
    mat_C[141][2] <=
                mat_A[136][0] * mat_B[5][2] +
                mat_A[136][1] * mat_B[13][2] +
                mat_A[136][2] * mat_B[21][2] +
                mat_A[136][3] * mat_B[29][2] +
                mat_A[137][0] * mat_B[37][2] +
                mat_A[137][1] * mat_B[45][2] +
                mat_A[137][2] * mat_B[53][2] +
                mat_A[137][3] * mat_B[61][2] +
                mat_A[138][0] * mat_B[69][2] +
                mat_A[138][1] * mat_B[77][2] +
                mat_A[138][2] * mat_B[85][2] +
                mat_A[138][3] * mat_B[93][2] +
                mat_A[139][0] * mat_B[101][2] +
                mat_A[139][1] * mat_B[109][2] +
                mat_A[139][2] * mat_B[117][2] +
                mat_A[139][3] * mat_B[125][2] +
                mat_A[140][0] * mat_B[133][2] +
                mat_A[140][1] * mat_B[141][2] +
                mat_A[140][2] * mat_B[149][2] +
                mat_A[140][3] * mat_B[157][2] +
                mat_A[141][0] * mat_B[165][2] +
                mat_A[141][1] * mat_B[173][2] +
                mat_A[141][2] * mat_B[181][2] +
                mat_A[141][3] * mat_B[189][2] +
                mat_A[142][0] * mat_B[197][2] +
                mat_A[142][1] * mat_B[205][2] +
                mat_A[142][2] * mat_B[213][2] +
                mat_A[142][3] * mat_B[221][2] +
                mat_A[143][0] * mat_B[229][2] +
                mat_A[143][1] * mat_B[237][2] +
                mat_A[143][2] * mat_B[245][2] +
                mat_A[143][3] * mat_B[253][2];
    mat_C[141][3] <=
                mat_A[136][0] * mat_B[5][3] +
                mat_A[136][1] * mat_B[13][3] +
                mat_A[136][2] * mat_B[21][3] +
                mat_A[136][3] * mat_B[29][3] +
                mat_A[137][0] * mat_B[37][3] +
                mat_A[137][1] * mat_B[45][3] +
                mat_A[137][2] * mat_B[53][3] +
                mat_A[137][3] * mat_B[61][3] +
                mat_A[138][0] * mat_B[69][3] +
                mat_A[138][1] * mat_B[77][3] +
                mat_A[138][2] * mat_B[85][3] +
                mat_A[138][3] * mat_B[93][3] +
                mat_A[139][0] * mat_B[101][3] +
                mat_A[139][1] * mat_B[109][3] +
                mat_A[139][2] * mat_B[117][3] +
                mat_A[139][3] * mat_B[125][3] +
                mat_A[140][0] * mat_B[133][3] +
                mat_A[140][1] * mat_B[141][3] +
                mat_A[140][2] * mat_B[149][3] +
                mat_A[140][3] * mat_B[157][3] +
                mat_A[141][0] * mat_B[165][3] +
                mat_A[141][1] * mat_B[173][3] +
                mat_A[141][2] * mat_B[181][3] +
                mat_A[141][3] * mat_B[189][3] +
                mat_A[142][0] * mat_B[197][3] +
                mat_A[142][1] * mat_B[205][3] +
                mat_A[142][2] * mat_B[213][3] +
                mat_A[142][3] * mat_B[221][3] +
                mat_A[143][0] * mat_B[229][3] +
                mat_A[143][1] * mat_B[237][3] +
                mat_A[143][2] * mat_B[245][3] +
                mat_A[143][3] * mat_B[253][3];
    mat_C[142][0] <=
                mat_A[136][0] * mat_B[6][0] +
                mat_A[136][1] * mat_B[14][0] +
                mat_A[136][2] * mat_B[22][0] +
                mat_A[136][3] * mat_B[30][0] +
                mat_A[137][0] * mat_B[38][0] +
                mat_A[137][1] * mat_B[46][0] +
                mat_A[137][2] * mat_B[54][0] +
                mat_A[137][3] * mat_B[62][0] +
                mat_A[138][0] * mat_B[70][0] +
                mat_A[138][1] * mat_B[78][0] +
                mat_A[138][2] * mat_B[86][0] +
                mat_A[138][3] * mat_B[94][0] +
                mat_A[139][0] * mat_B[102][0] +
                mat_A[139][1] * mat_B[110][0] +
                mat_A[139][2] * mat_B[118][0] +
                mat_A[139][3] * mat_B[126][0] +
                mat_A[140][0] * mat_B[134][0] +
                mat_A[140][1] * mat_B[142][0] +
                mat_A[140][2] * mat_B[150][0] +
                mat_A[140][3] * mat_B[158][0] +
                mat_A[141][0] * mat_B[166][0] +
                mat_A[141][1] * mat_B[174][0] +
                mat_A[141][2] * mat_B[182][0] +
                mat_A[141][3] * mat_B[190][0] +
                mat_A[142][0] * mat_B[198][0] +
                mat_A[142][1] * mat_B[206][0] +
                mat_A[142][2] * mat_B[214][0] +
                mat_A[142][3] * mat_B[222][0] +
                mat_A[143][0] * mat_B[230][0] +
                mat_A[143][1] * mat_B[238][0] +
                mat_A[143][2] * mat_B[246][0] +
                mat_A[143][3] * mat_B[254][0];
    mat_C[142][1] <=
                mat_A[136][0] * mat_B[6][1] +
                mat_A[136][1] * mat_B[14][1] +
                mat_A[136][2] * mat_B[22][1] +
                mat_A[136][3] * mat_B[30][1] +
                mat_A[137][0] * mat_B[38][1] +
                mat_A[137][1] * mat_B[46][1] +
                mat_A[137][2] * mat_B[54][1] +
                mat_A[137][3] * mat_B[62][1] +
                mat_A[138][0] * mat_B[70][1] +
                mat_A[138][1] * mat_B[78][1] +
                mat_A[138][2] * mat_B[86][1] +
                mat_A[138][3] * mat_B[94][1] +
                mat_A[139][0] * mat_B[102][1] +
                mat_A[139][1] * mat_B[110][1] +
                mat_A[139][2] * mat_B[118][1] +
                mat_A[139][3] * mat_B[126][1] +
                mat_A[140][0] * mat_B[134][1] +
                mat_A[140][1] * mat_B[142][1] +
                mat_A[140][2] * mat_B[150][1] +
                mat_A[140][3] * mat_B[158][1] +
                mat_A[141][0] * mat_B[166][1] +
                mat_A[141][1] * mat_B[174][1] +
                mat_A[141][2] * mat_B[182][1] +
                mat_A[141][3] * mat_B[190][1] +
                mat_A[142][0] * mat_B[198][1] +
                mat_A[142][1] * mat_B[206][1] +
                mat_A[142][2] * mat_B[214][1] +
                mat_A[142][3] * mat_B[222][1] +
                mat_A[143][0] * mat_B[230][1] +
                mat_A[143][1] * mat_B[238][1] +
                mat_A[143][2] * mat_B[246][1] +
                mat_A[143][3] * mat_B[254][1];
    mat_C[142][2] <=
                mat_A[136][0] * mat_B[6][2] +
                mat_A[136][1] * mat_B[14][2] +
                mat_A[136][2] * mat_B[22][2] +
                mat_A[136][3] * mat_B[30][2] +
                mat_A[137][0] * mat_B[38][2] +
                mat_A[137][1] * mat_B[46][2] +
                mat_A[137][2] * mat_B[54][2] +
                mat_A[137][3] * mat_B[62][2] +
                mat_A[138][0] * mat_B[70][2] +
                mat_A[138][1] * mat_B[78][2] +
                mat_A[138][2] * mat_B[86][2] +
                mat_A[138][3] * mat_B[94][2] +
                mat_A[139][0] * mat_B[102][2] +
                mat_A[139][1] * mat_B[110][2] +
                mat_A[139][2] * mat_B[118][2] +
                mat_A[139][3] * mat_B[126][2] +
                mat_A[140][0] * mat_B[134][2] +
                mat_A[140][1] * mat_B[142][2] +
                mat_A[140][2] * mat_B[150][2] +
                mat_A[140][3] * mat_B[158][2] +
                mat_A[141][0] * mat_B[166][2] +
                mat_A[141][1] * mat_B[174][2] +
                mat_A[141][2] * mat_B[182][2] +
                mat_A[141][3] * mat_B[190][2] +
                mat_A[142][0] * mat_B[198][2] +
                mat_A[142][1] * mat_B[206][2] +
                mat_A[142][2] * mat_B[214][2] +
                mat_A[142][3] * mat_B[222][2] +
                mat_A[143][0] * mat_B[230][2] +
                mat_A[143][1] * mat_B[238][2] +
                mat_A[143][2] * mat_B[246][2] +
                mat_A[143][3] * mat_B[254][2];
    mat_C[142][3] <=
                mat_A[136][0] * mat_B[6][3] +
                mat_A[136][1] * mat_B[14][3] +
                mat_A[136][2] * mat_B[22][3] +
                mat_A[136][3] * mat_B[30][3] +
                mat_A[137][0] * mat_B[38][3] +
                mat_A[137][1] * mat_B[46][3] +
                mat_A[137][2] * mat_B[54][3] +
                mat_A[137][3] * mat_B[62][3] +
                mat_A[138][0] * mat_B[70][3] +
                mat_A[138][1] * mat_B[78][3] +
                mat_A[138][2] * mat_B[86][3] +
                mat_A[138][3] * mat_B[94][3] +
                mat_A[139][0] * mat_B[102][3] +
                mat_A[139][1] * mat_B[110][3] +
                mat_A[139][2] * mat_B[118][3] +
                mat_A[139][3] * mat_B[126][3] +
                mat_A[140][0] * mat_B[134][3] +
                mat_A[140][1] * mat_B[142][3] +
                mat_A[140][2] * mat_B[150][3] +
                mat_A[140][3] * mat_B[158][3] +
                mat_A[141][0] * mat_B[166][3] +
                mat_A[141][1] * mat_B[174][3] +
                mat_A[141][2] * mat_B[182][3] +
                mat_A[141][3] * mat_B[190][3] +
                mat_A[142][0] * mat_B[198][3] +
                mat_A[142][1] * mat_B[206][3] +
                mat_A[142][2] * mat_B[214][3] +
                mat_A[142][3] * mat_B[222][3] +
                mat_A[143][0] * mat_B[230][3] +
                mat_A[143][1] * mat_B[238][3] +
                mat_A[143][2] * mat_B[246][3] +
                mat_A[143][3] * mat_B[254][3];
    mat_C[143][0] <=
                mat_A[136][0] * mat_B[7][0] +
                mat_A[136][1] * mat_B[15][0] +
                mat_A[136][2] * mat_B[23][0] +
                mat_A[136][3] * mat_B[31][0] +
                mat_A[137][0] * mat_B[39][0] +
                mat_A[137][1] * mat_B[47][0] +
                mat_A[137][2] * mat_B[55][0] +
                mat_A[137][3] * mat_B[63][0] +
                mat_A[138][0] * mat_B[71][0] +
                mat_A[138][1] * mat_B[79][0] +
                mat_A[138][2] * mat_B[87][0] +
                mat_A[138][3] * mat_B[95][0] +
                mat_A[139][0] * mat_B[103][0] +
                mat_A[139][1] * mat_B[111][0] +
                mat_A[139][2] * mat_B[119][0] +
                mat_A[139][3] * mat_B[127][0] +
                mat_A[140][0] * mat_B[135][0] +
                mat_A[140][1] * mat_B[143][0] +
                mat_A[140][2] * mat_B[151][0] +
                mat_A[140][3] * mat_B[159][0] +
                mat_A[141][0] * mat_B[167][0] +
                mat_A[141][1] * mat_B[175][0] +
                mat_A[141][2] * mat_B[183][0] +
                mat_A[141][3] * mat_B[191][0] +
                mat_A[142][0] * mat_B[199][0] +
                mat_A[142][1] * mat_B[207][0] +
                mat_A[142][2] * mat_B[215][0] +
                mat_A[142][3] * mat_B[223][0] +
                mat_A[143][0] * mat_B[231][0] +
                mat_A[143][1] * mat_B[239][0] +
                mat_A[143][2] * mat_B[247][0] +
                mat_A[143][3] * mat_B[255][0];
    mat_C[143][1] <=
                mat_A[136][0] * mat_B[7][1] +
                mat_A[136][1] * mat_B[15][1] +
                mat_A[136][2] * mat_B[23][1] +
                mat_A[136][3] * mat_B[31][1] +
                mat_A[137][0] * mat_B[39][1] +
                mat_A[137][1] * mat_B[47][1] +
                mat_A[137][2] * mat_B[55][1] +
                mat_A[137][3] * mat_B[63][1] +
                mat_A[138][0] * mat_B[71][1] +
                mat_A[138][1] * mat_B[79][1] +
                mat_A[138][2] * mat_B[87][1] +
                mat_A[138][3] * mat_B[95][1] +
                mat_A[139][0] * mat_B[103][1] +
                mat_A[139][1] * mat_B[111][1] +
                mat_A[139][2] * mat_B[119][1] +
                mat_A[139][3] * mat_B[127][1] +
                mat_A[140][0] * mat_B[135][1] +
                mat_A[140][1] * mat_B[143][1] +
                mat_A[140][2] * mat_B[151][1] +
                mat_A[140][3] * mat_B[159][1] +
                mat_A[141][0] * mat_B[167][1] +
                mat_A[141][1] * mat_B[175][1] +
                mat_A[141][2] * mat_B[183][1] +
                mat_A[141][3] * mat_B[191][1] +
                mat_A[142][0] * mat_B[199][1] +
                mat_A[142][1] * mat_B[207][1] +
                mat_A[142][2] * mat_B[215][1] +
                mat_A[142][3] * mat_B[223][1] +
                mat_A[143][0] * mat_B[231][1] +
                mat_A[143][1] * mat_B[239][1] +
                mat_A[143][2] * mat_B[247][1] +
                mat_A[143][3] * mat_B[255][1];
    mat_C[143][2] <=
                mat_A[136][0] * mat_B[7][2] +
                mat_A[136][1] * mat_B[15][2] +
                mat_A[136][2] * mat_B[23][2] +
                mat_A[136][3] * mat_B[31][2] +
                mat_A[137][0] * mat_B[39][2] +
                mat_A[137][1] * mat_B[47][2] +
                mat_A[137][2] * mat_B[55][2] +
                mat_A[137][3] * mat_B[63][2] +
                mat_A[138][0] * mat_B[71][2] +
                mat_A[138][1] * mat_B[79][2] +
                mat_A[138][2] * mat_B[87][2] +
                mat_A[138][3] * mat_B[95][2] +
                mat_A[139][0] * mat_B[103][2] +
                mat_A[139][1] * mat_B[111][2] +
                mat_A[139][2] * mat_B[119][2] +
                mat_A[139][3] * mat_B[127][2] +
                mat_A[140][0] * mat_B[135][2] +
                mat_A[140][1] * mat_B[143][2] +
                mat_A[140][2] * mat_B[151][2] +
                mat_A[140][3] * mat_B[159][2] +
                mat_A[141][0] * mat_B[167][2] +
                mat_A[141][1] * mat_B[175][2] +
                mat_A[141][2] * mat_B[183][2] +
                mat_A[141][3] * mat_B[191][2] +
                mat_A[142][0] * mat_B[199][2] +
                mat_A[142][1] * mat_B[207][2] +
                mat_A[142][2] * mat_B[215][2] +
                mat_A[142][3] * mat_B[223][2] +
                mat_A[143][0] * mat_B[231][2] +
                mat_A[143][1] * mat_B[239][2] +
                mat_A[143][2] * mat_B[247][2] +
                mat_A[143][3] * mat_B[255][2];
    mat_C[143][3] <=
                mat_A[136][0] * mat_B[7][3] +
                mat_A[136][1] * mat_B[15][3] +
                mat_A[136][2] * mat_B[23][3] +
                mat_A[136][3] * mat_B[31][3] +
                mat_A[137][0] * mat_B[39][3] +
                mat_A[137][1] * mat_B[47][3] +
                mat_A[137][2] * mat_B[55][3] +
                mat_A[137][3] * mat_B[63][3] +
                mat_A[138][0] * mat_B[71][3] +
                mat_A[138][1] * mat_B[79][3] +
                mat_A[138][2] * mat_B[87][3] +
                mat_A[138][3] * mat_B[95][3] +
                mat_A[139][0] * mat_B[103][3] +
                mat_A[139][1] * mat_B[111][3] +
                mat_A[139][2] * mat_B[119][3] +
                mat_A[139][3] * mat_B[127][3] +
                mat_A[140][0] * mat_B[135][3] +
                mat_A[140][1] * mat_B[143][3] +
                mat_A[140][2] * mat_B[151][3] +
                mat_A[140][3] * mat_B[159][3] +
                mat_A[141][0] * mat_B[167][3] +
                mat_A[141][1] * mat_B[175][3] +
                mat_A[141][2] * mat_B[183][3] +
                mat_A[141][3] * mat_B[191][3] +
                mat_A[142][0] * mat_B[199][3] +
                mat_A[142][1] * mat_B[207][3] +
                mat_A[142][2] * mat_B[215][3] +
                mat_A[142][3] * mat_B[223][3] +
                mat_A[143][0] * mat_B[231][3] +
                mat_A[143][1] * mat_B[239][3] +
                mat_A[143][2] * mat_B[247][3] +
                mat_A[143][3] * mat_B[255][3];
    mat_C[144][0] <=
                mat_A[144][0] * mat_B[0][0] +
                mat_A[144][1] * mat_B[8][0] +
                mat_A[144][2] * mat_B[16][0] +
                mat_A[144][3] * mat_B[24][0] +
                mat_A[145][0] * mat_B[32][0] +
                mat_A[145][1] * mat_B[40][0] +
                mat_A[145][2] * mat_B[48][0] +
                mat_A[145][3] * mat_B[56][0] +
                mat_A[146][0] * mat_B[64][0] +
                mat_A[146][1] * mat_B[72][0] +
                mat_A[146][2] * mat_B[80][0] +
                mat_A[146][3] * mat_B[88][0] +
                mat_A[147][0] * mat_B[96][0] +
                mat_A[147][1] * mat_B[104][0] +
                mat_A[147][2] * mat_B[112][0] +
                mat_A[147][3] * mat_B[120][0] +
                mat_A[148][0] * mat_B[128][0] +
                mat_A[148][1] * mat_B[136][0] +
                mat_A[148][2] * mat_B[144][0] +
                mat_A[148][3] * mat_B[152][0] +
                mat_A[149][0] * mat_B[160][0] +
                mat_A[149][1] * mat_B[168][0] +
                mat_A[149][2] * mat_B[176][0] +
                mat_A[149][3] * mat_B[184][0] +
                mat_A[150][0] * mat_B[192][0] +
                mat_A[150][1] * mat_B[200][0] +
                mat_A[150][2] * mat_B[208][0] +
                mat_A[150][3] * mat_B[216][0] +
                mat_A[151][0] * mat_B[224][0] +
                mat_A[151][1] * mat_B[232][0] +
                mat_A[151][2] * mat_B[240][0] +
                mat_A[151][3] * mat_B[248][0];
    mat_C[144][1] <=
                mat_A[144][0] * mat_B[0][1] +
                mat_A[144][1] * mat_B[8][1] +
                mat_A[144][2] * mat_B[16][1] +
                mat_A[144][3] * mat_B[24][1] +
                mat_A[145][0] * mat_B[32][1] +
                mat_A[145][1] * mat_B[40][1] +
                mat_A[145][2] * mat_B[48][1] +
                mat_A[145][3] * mat_B[56][1] +
                mat_A[146][0] * mat_B[64][1] +
                mat_A[146][1] * mat_B[72][1] +
                mat_A[146][2] * mat_B[80][1] +
                mat_A[146][3] * mat_B[88][1] +
                mat_A[147][0] * mat_B[96][1] +
                mat_A[147][1] * mat_B[104][1] +
                mat_A[147][2] * mat_B[112][1] +
                mat_A[147][3] * mat_B[120][1] +
                mat_A[148][0] * mat_B[128][1] +
                mat_A[148][1] * mat_B[136][1] +
                mat_A[148][2] * mat_B[144][1] +
                mat_A[148][3] * mat_B[152][1] +
                mat_A[149][0] * mat_B[160][1] +
                mat_A[149][1] * mat_B[168][1] +
                mat_A[149][2] * mat_B[176][1] +
                mat_A[149][3] * mat_B[184][1] +
                mat_A[150][0] * mat_B[192][1] +
                mat_A[150][1] * mat_B[200][1] +
                mat_A[150][2] * mat_B[208][1] +
                mat_A[150][3] * mat_B[216][1] +
                mat_A[151][0] * mat_B[224][1] +
                mat_A[151][1] * mat_B[232][1] +
                mat_A[151][2] * mat_B[240][1] +
                mat_A[151][3] * mat_B[248][1];
    mat_C[144][2] <=
                mat_A[144][0] * mat_B[0][2] +
                mat_A[144][1] * mat_B[8][2] +
                mat_A[144][2] * mat_B[16][2] +
                mat_A[144][3] * mat_B[24][2] +
                mat_A[145][0] * mat_B[32][2] +
                mat_A[145][1] * mat_B[40][2] +
                mat_A[145][2] * mat_B[48][2] +
                mat_A[145][3] * mat_B[56][2] +
                mat_A[146][0] * mat_B[64][2] +
                mat_A[146][1] * mat_B[72][2] +
                mat_A[146][2] * mat_B[80][2] +
                mat_A[146][3] * mat_B[88][2] +
                mat_A[147][0] * mat_B[96][2] +
                mat_A[147][1] * mat_B[104][2] +
                mat_A[147][2] * mat_B[112][2] +
                mat_A[147][3] * mat_B[120][2] +
                mat_A[148][0] * mat_B[128][2] +
                mat_A[148][1] * mat_B[136][2] +
                mat_A[148][2] * mat_B[144][2] +
                mat_A[148][3] * mat_B[152][2] +
                mat_A[149][0] * mat_B[160][2] +
                mat_A[149][1] * mat_B[168][2] +
                mat_A[149][2] * mat_B[176][2] +
                mat_A[149][3] * mat_B[184][2] +
                mat_A[150][0] * mat_B[192][2] +
                mat_A[150][1] * mat_B[200][2] +
                mat_A[150][2] * mat_B[208][2] +
                mat_A[150][3] * mat_B[216][2] +
                mat_A[151][0] * mat_B[224][2] +
                mat_A[151][1] * mat_B[232][2] +
                mat_A[151][2] * mat_B[240][2] +
                mat_A[151][3] * mat_B[248][2];
    mat_C[144][3] <=
                mat_A[144][0] * mat_B[0][3] +
                mat_A[144][1] * mat_B[8][3] +
                mat_A[144][2] * mat_B[16][3] +
                mat_A[144][3] * mat_B[24][3] +
                mat_A[145][0] * mat_B[32][3] +
                mat_A[145][1] * mat_B[40][3] +
                mat_A[145][2] * mat_B[48][3] +
                mat_A[145][3] * mat_B[56][3] +
                mat_A[146][0] * mat_B[64][3] +
                mat_A[146][1] * mat_B[72][3] +
                mat_A[146][2] * mat_B[80][3] +
                mat_A[146][3] * mat_B[88][3] +
                mat_A[147][0] * mat_B[96][3] +
                mat_A[147][1] * mat_B[104][3] +
                mat_A[147][2] * mat_B[112][3] +
                mat_A[147][3] * mat_B[120][3] +
                mat_A[148][0] * mat_B[128][3] +
                mat_A[148][1] * mat_B[136][3] +
                mat_A[148][2] * mat_B[144][3] +
                mat_A[148][3] * mat_B[152][3] +
                mat_A[149][0] * mat_B[160][3] +
                mat_A[149][1] * mat_B[168][3] +
                mat_A[149][2] * mat_B[176][3] +
                mat_A[149][3] * mat_B[184][3] +
                mat_A[150][0] * mat_B[192][3] +
                mat_A[150][1] * mat_B[200][3] +
                mat_A[150][2] * mat_B[208][3] +
                mat_A[150][3] * mat_B[216][3] +
                mat_A[151][0] * mat_B[224][3] +
                mat_A[151][1] * mat_B[232][3] +
                mat_A[151][2] * mat_B[240][3] +
                mat_A[151][3] * mat_B[248][3];
    mat_C[145][0] <=
                mat_A[144][0] * mat_B[1][0] +
                mat_A[144][1] * mat_B[9][0] +
                mat_A[144][2] * mat_B[17][0] +
                mat_A[144][3] * mat_B[25][0] +
                mat_A[145][0] * mat_B[33][0] +
                mat_A[145][1] * mat_B[41][0] +
                mat_A[145][2] * mat_B[49][0] +
                mat_A[145][3] * mat_B[57][0] +
                mat_A[146][0] * mat_B[65][0] +
                mat_A[146][1] * mat_B[73][0] +
                mat_A[146][2] * mat_B[81][0] +
                mat_A[146][3] * mat_B[89][0] +
                mat_A[147][0] * mat_B[97][0] +
                mat_A[147][1] * mat_B[105][0] +
                mat_A[147][2] * mat_B[113][0] +
                mat_A[147][3] * mat_B[121][0] +
                mat_A[148][0] * mat_B[129][0] +
                mat_A[148][1] * mat_B[137][0] +
                mat_A[148][2] * mat_B[145][0] +
                mat_A[148][3] * mat_B[153][0] +
                mat_A[149][0] * mat_B[161][0] +
                mat_A[149][1] * mat_B[169][0] +
                mat_A[149][2] * mat_B[177][0] +
                mat_A[149][3] * mat_B[185][0] +
                mat_A[150][0] * mat_B[193][0] +
                mat_A[150][1] * mat_B[201][0] +
                mat_A[150][2] * mat_B[209][0] +
                mat_A[150][3] * mat_B[217][0] +
                mat_A[151][0] * mat_B[225][0] +
                mat_A[151][1] * mat_B[233][0] +
                mat_A[151][2] * mat_B[241][0] +
                mat_A[151][3] * mat_B[249][0];
    mat_C[145][1] <=
                mat_A[144][0] * mat_B[1][1] +
                mat_A[144][1] * mat_B[9][1] +
                mat_A[144][2] * mat_B[17][1] +
                mat_A[144][3] * mat_B[25][1] +
                mat_A[145][0] * mat_B[33][1] +
                mat_A[145][1] * mat_B[41][1] +
                mat_A[145][2] * mat_B[49][1] +
                mat_A[145][3] * mat_B[57][1] +
                mat_A[146][0] * mat_B[65][1] +
                mat_A[146][1] * mat_B[73][1] +
                mat_A[146][2] * mat_B[81][1] +
                mat_A[146][3] * mat_B[89][1] +
                mat_A[147][0] * mat_B[97][1] +
                mat_A[147][1] * mat_B[105][1] +
                mat_A[147][2] * mat_B[113][1] +
                mat_A[147][3] * mat_B[121][1] +
                mat_A[148][0] * mat_B[129][1] +
                mat_A[148][1] * mat_B[137][1] +
                mat_A[148][2] * mat_B[145][1] +
                mat_A[148][3] * mat_B[153][1] +
                mat_A[149][0] * mat_B[161][1] +
                mat_A[149][1] * mat_B[169][1] +
                mat_A[149][2] * mat_B[177][1] +
                mat_A[149][3] * mat_B[185][1] +
                mat_A[150][0] * mat_B[193][1] +
                mat_A[150][1] * mat_B[201][1] +
                mat_A[150][2] * mat_B[209][1] +
                mat_A[150][3] * mat_B[217][1] +
                mat_A[151][0] * mat_B[225][1] +
                mat_A[151][1] * mat_B[233][1] +
                mat_A[151][2] * mat_B[241][1] +
                mat_A[151][3] * mat_B[249][1];
    mat_C[145][2] <=
                mat_A[144][0] * mat_B[1][2] +
                mat_A[144][1] * mat_B[9][2] +
                mat_A[144][2] * mat_B[17][2] +
                mat_A[144][3] * mat_B[25][2] +
                mat_A[145][0] * mat_B[33][2] +
                mat_A[145][1] * mat_B[41][2] +
                mat_A[145][2] * mat_B[49][2] +
                mat_A[145][3] * mat_B[57][2] +
                mat_A[146][0] * mat_B[65][2] +
                mat_A[146][1] * mat_B[73][2] +
                mat_A[146][2] * mat_B[81][2] +
                mat_A[146][3] * mat_B[89][2] +
                mat_A[147][0] * mat_B[97][2] +
                mat_A[147][1] * mat_B[105][2] +
                mat_A[147][2] * mat_B[113][2] +
                mat_A[147][3] * mat_B[121][2] +
                mat_A[148][0] * mat_B[129][2] +
                mat_A[148][1] * mat_B[137][2] +
                mat_A[148][2] * mat_B[145][2] +
                mat_A[148][3] * mat_B[153][2] +
                mat_A[149][0] * mat_B[161][2] +
                mat_A[149][1] * mat_B[169][2] +
                mat_A[149][2] * mat_B[177][2] +
                mat_A[149][3] * mat_B[185][2] +
                mat_A[150][0] * mat_B[193][2] +
                mat_A[150][1] * mat_B[201][2] +
                mat_A[150][2] * mat_B[209][2] +
                mat_A[150][3] * mat_B[217][2] +
                mat_A[151][0] * mat_B[225][2] +
                mat_A[151][1] * mat_B[233][2] +
                mat_A[151][2] * mat_B[241][2] +
                mat_A[151][3] * mat_B[249][2];
    mat_C[145][3] <=
                mat_A[144][0] * mat_B[1][3] +
                mat_A[144][1] * mat_B[9][3] +
                mat_A[144][2] * mat_B[17][3] +
                mat_A[144][3] * mat_B[25][3] +
                mat_A[145][0] * mat_B[33][3] +
                mat_A[145][1] * mat_B[41][3] +
                mat_A[145][2] * mat_B[49][3] +
                mat_A[145][3] * mat_B[57][3] +
                mat_A[146][0] * mat_B[65][3] +
                mat_A[146][1] * mat_B[73][3] +
                mat_A[146][2] * mat_B[81][3] +
                mat_A[146][3] * mat_B[89][3] +
                mat_A[147][0] * mat_B[97][3] +
                mat_A[147][1] * mat_B[105][3] +
                mat_A[147][2] * mat_B[113][3] +
                mat_A[147][3] * mat_B[121][3] +
                mat_A[148][0] * mat_B[129][3] +
                mat_A[148][1] * mat_B[137][3] +
                mat_A[148][2] * mat_B[145][3] +
                mat_A[148][3] * mat_B[153][3] +
                mat_A[149][0] * mat_B[161][3] +
                mat_A[149][1] * mat_B[169][3] +
                mat_A[149][2] * mat_B[177][3] +
                mat_A[149][3] * mat_B[185][3] +
                mat_A[150][0] * mat_B[193][3] +
                mat_A[150][1] * mat_B[201][3] +
                mat_A[150][2] * mat_B[209][3] +
                mat_A[150][3] * mat_B[217][3] +
                mat_A[151][0] * mat_B[225][3] +
                mat_A[151][1] * mat_B[233][3] +
                mat_A[151][2] * mat_B[241][3] +
                mat_A[151][3] * mat_B[249][3];
    mat_C[146][0] <=
                mat_A[144][0] * mat_B[2][0] +
                mat_A[144][1] * mat_B[10][0] +
                mat_A[144][2] * mat_B[18][0] +
                mat_A[144][3] * mat_B[26][0] +
                mat_A[145][0] * mat_B[34][0] +
                mat_A[145][1] * mat_B[42][0] +
                mat_A[145][2] * mat_B[50][0] +
                mat_A[145][3] * mat_B[58][0] +
                mat_A[146][0] * mat_B[66][0] +
                mat_A[146][1] * mat_B[74][0] +
                mat_A[146][2] * mat_B[82][0] +
                mat_A[146][3] * mat_B[90][0] +
                mat_A[147][0] * mat_B[98][0] +
                mat_A[147][1] * mat_B[106][0] +
                mat_A[147][2] * mat_B[114][0] +
                mat_A[147][3] * mat_B[122][0] +
                mat_A[148][0] * mat_B[130][0] +
                mat_A[148][1] * mat_B[138][0] +
                mat_A[148][2] * mat_B[146][0] +
                mat_A[148][3] * mat_B[154][0] +
                mat_A[149][0] * mat_B[162][0] +
                mat_A[149][1] * mat_B[170][0] +
                mat_A[149][2] * mat_B[178][0] +
                mat_A[149][3] * mat_B[186][0] +
                mat_A[150][0] * mat_B[194][0] +
                mat_A[150][1] * mat_B[202][0] +
                mat_A[150][2] * mat_B[210][0] +
                mat_A[150][3] * mat_B[218][0] +
                mat_A[151][0] * mat_B[226][0] +
                mat_A[151][1] * mat_B[234][0] +
                mat_A[151][2] * mat_B[242][0] +
                mat_A[151][3] * mat_B[250][0];
    mat_C[146][1] <=
                mat_A[144][0] * mat_B[2][1] +
                mat_A[144][1] * mat_B[10][1] +
                mat_A[144][2] * mat_B[18][1] +
                mat_A[144][3] * mat_B[26][1] +
                mat_A[145][0] * mat_B[34][1] +
                mat_A[145][1] * mat_B[42][1] +
                mat_A[145][2] * mat_B[50][1] +
                mat_A[145][3] * mat_B[58][1] +
                mat_A[146][0] * mat_B[66][1] +
                mat_A[146][1] * mat_B[74][1] +
                mat_A[146][2] * mat_B[82][1] +
                mat_A[146][3] * mat_B[90][1] +
                mat_A[147][0] * mat_B[98][1] +
                mat_A[147][1] * mat_B[106][1] +
                mat_A[147][2] * mat_B[114][1] +
                mat_A[147][3] * mat_B[122][1] +
                mat_A[148][0] * mat_B[130][1] +
                mat_A[148][1] * mat_B[138][1] +
                mat_A[148][2] * mat_B[146][1] +
                mat_A[148][3] * mat_B[154][1] +
                mat_A[149][0] * mat_B[162][1] +
                mat_A[149][1] * mat_B[170][1] +
                mat_A[149][2] * mat_B[178][1] +
                mat_A[149][3] * mat_B[186][1] +
                mat_A[150][0] * mat_B[194][1] +
                mat_A[150][1] * mat_B[202][1] +
                mat_A[150][2] * mat_B[210][1] +
                mat_A[150][3] * mat_B[218][1] +
                mat_A[151][0] * mat_B[226][1] +
                mat_A[151][1] * mat_B[234][1] +
                mat_A[151][2] * mat_B[242][1] +
                mat_A[151][3] * mat_B[250][1];
    mat_C[146][2] <=
                mat_A[144][0] * mat_B[2][2] +
                mat_A[144][1] * mat_B[10][2] +
                mat_A[144][2] * mat_B[18][2] +
                mat_A[144][3] * mat_B[26][2] +
                mat_A[145][0] * mat_B[34][2] +
                mat_A[145][1] * mat_B[42][2] +
                mat_A[145][2] * mat_B[50][2] +
                mat_A[145][3] * mat_B[58][2] +
                mat_A[146][0] * mat_B[66][2] +
                mat_A[146][1] * mat_B[74][2] +
                mat_A[146][2] * mat_B[82][2] +
                mat_A[146][3] * mat_B[90][2] +
                mat_A[147][0] * mat_B[98][2] +
                mat_A[147][1] * mat_B[106][2] +
                mat_A[147][2] * mat_B[114][2] +
                mat_A[147][3] * mat_B[122][2] +
                mat_A[148][0] * mat_B[130][2] +
                mat_A[148][1] * mat_B[138][2] +
                mat_A[148][2] * mat_B[146][2] +
                mat_A[148][3] * mat_B[154][2] +
                mat_A[149][0] * mat_B[162][2] +
                mat_A[149][1] * mat_B[170][2] +
                mat_A[149][2] * mat_B[178][2] +
                mat_A[149][3] * mat_B[186][2] +
                mat_A[150][0] * mat_B[194][2] +
                mat_A[150][1] * mat_B[202][2] +
                mat_A[150][2] * mat_B[210][2] +
                mat_A[150][3] * mat_B[218][2] +
                mat_A[151][0] * mat_B[226][2] +
                mat_A[151][1] * mat_B[234][2] +
                mat_A[151][2] * mat_B[242][2] +
                mat_A[151][3] * mat_B[250][2];
    mat_C[146][3] <=
                mat_A[144][0] * mat_B[2][3] +
                mat_A[144][1] * mat_B[10][3] +
                mat_A[144][2] * mat_B[18][3] +
                mat_A[144][3] * mat_B[26][3] +
                mat_A[145][0] * mat_B[34][3] +
                mat_A[145][1] * mat_B[42][3] +
                mat_A[145][2] * mat_B[50][3] +
                mat_A[145][3] * mat_B[58][3] +
                mat_A[146][0] * mat_B[66][3] +
                mat_A[146][1] * mat_B[74][3] +
                mat_A[146][2] * mat_B[82][3] +
                mat_A[146][3] * mat_B[90][3] +
                mat_A[147][0] * mat_B[98][3] +
                mat_A[147][1] * mat_B[106][3] +
                mat_A[147][2] * mat_B[114][3] +
                mat_A[147][3] * mat_B[122][3] +
                mat_A[148][0] * mat_B[130][3] +
                mat_A[148][1] * mat_B[138][3] +
                mat_A[148][2] * mat_B[146][3] +
                mat_A[148][3] * mat_B[154][3] +
                mat_A[149][0] * mat_B[162][3] +
                mat_A[149][1] * mat_B[170][3] +
                mat_A[149][2] * mat_B[178][3] +
                mat_A[149][3] * mat_B[186][3] +
                mat_A[150][0] * mat_B[194][3] +
                mat_A[150][1] * mat_B[202][3] +
                mat_A[150][2] * mat_B[210][3] +
                mat_A[150][3] * mat_B[218][3] +
                mat_A[151][0] * mat_B[226][3] +
                mat_A[151][1] * mat_B[234][3] +
                mat_A[151][2] * mat_B[242][3] +
                mat_A[151][3] * mat_B[250][3];
    mat_C[147][0] <=
                mat_A[144][0] * mat_B[3][0] +
                mat_A[144][1] * mat_B[11][0] +
                mat_A[144][2] * mat_B[19][0] +
                mat_A[144][3] * mat_B[27][0] +
                mat_A[145][0] * mat_B[35][0] +
                mat_A[145][1] * mat_B[43][0] +
                mat_A[145][2] * mat_B[51][0] +
                mat_A[145][3] * mat_B[59][0] +
                mat_A[146][0] * mat_B[67][0] +
                mat_A[146][1] * mat_B[75][0] +
                mat_A[146][2] * mat_B[83][0] +
                mat_A[146][3] * mat_B[91][0] +
                mat_A[147][0] * mat_B[99][0] +
                mat_A[147][1] * mat_B[107][0] +
                mat_A[147][2] * mat_B[115][0] +
                mat_A[147][3] * mat_B[123][0] +
                mat_A[148][0] * mat_B[131][0] +
                mat_A[148][1] * mat_B[139][0] +
                mat_A[148][2] * mat_B[147][0] +
                mat_A[148][3] * mat_B[155][0] +
                mat_A[149][0] * mat_B[163][0] +
                mat_A[149][1] * mat_B[171][0] +
                mat_A[149][2] * mat_B[179][0] +
                mat_A[149][3] * mat_B[187][0] +
                mat_A[150][0] * mat_B[195][0] +
                mat_A[150][1] * mat_B[203][0] +
                mat_A[150][2] * mat_B[211][0] +
                mat_A[150][3] * mat_B[219][0] +
                mat_A[151][0] * mat_B[227][0] +
                mat_A[151][1] * mat_B[235][0] +
                mat_A[151][2] * mat_B[243][0] +
                mat_A[151][3] * mat_B[251][0];
    mat_C[147][1] <=
                mat_A[144][0] * mat_B[3][1] +
                mat_A[144][1] * mat_B[11][1] +
                mat_A[144][2] * mat_B[19][1] +
                mat_A[144][3] * mat_B[27][1] +
                mat_A[145][0] * mat_B[35][1] +
                mat_A[145][1] * mat_B[43][1] +
                mat_A[145][2] * mat_B[51][1] +
                mat_A[145][3] * mat_B[59][1] +
                mat_A[146][0] * mat_B[67][1] +
                mat_A[146][1] * mat_B[75][1] +
                mat_A[146][2] * mat_B[83][1] +
                mat_A[146][3] * mat_B[91][1] +
                mat_A[147][0] * mat_B[99][1] +
                mat_A[147][1] * mat_B[107][1] +
                mat_A[147][2] * mat_B[115][1] +
                mat_A[147][3] * mat_B[123][1] +
                mat_A[148][0] * mat_B[131][1] +
                mat_A[148][1] * mat_B[139][1] +
                mat_A[148][2] * mat_B[147][1] +
                mat_A[148][3] * mat_B[155][1] +
                mat_A[149][0] * mat_B[163][1] +
                mat_A[149][1] * mat_B[171][1] +
                mat_A[149][2] * mat_B[179][1] +
                mat_A[149][3] * mat_B[187][1] +
                mat_A[150][0] * mat_B[195][1] +
                mat_A[150][1] * mat_B[203][1] +
                mat_A[150][2] * mat_B[211][1] +
                mat_A[150][3] * mat_B[219][1] +
                mat_A[151][0] * mat_B[227][1] +
                mat_A[151][1] * mat_B[235][1] +
                mat_A[151][2] * mat_B[243][1] +
                mat_A[151][3] * mat_B[251][1];
    mat_C[147][2] <=
                mat_A[144][0] * mat_B[3][2] +
                mat_A[144][1] * mat_B[11][2] +
                mat_A[144][2] * mat_B[19][2] +
                mat_A[144][3] * mat_B[27][2] +
                mat_A[145][0] * mat_B[35][2] +
                mat_A[145][1] * mat_B[43][2] +
                mat_A[145][2] * mat_B[51][2] +
                mat_A[145][3] * mat_B[59][2] +
                mat_A[146][0] * mat_B[67][2] +
                mat_A[146][1] * mat_B[75][2] +
                mat_A[146][2] * mat_B[83][2] +
                mat_A[146][3] * mat_B[91][2] +
                mat_A[147][0] * mat_B[99][2] +
                mat_A[147][1] * mat_B[107][2] +
                mat_A[147][2] * mat_B[115][2] +
                mat_A[147][3] * mat_B[123][2] +
                mat_A[148][0] * mat_B[131][2] +
                mat_A[148][1] * mat_B[139][2] +
                mat_A[148][2] * mat_B[147][2] +
                mat_A[148][3] * mat_B[155][2] +
                mat_A[149][0] * mat_B[163][2] +
                mat_A[149][1] * mat_B[171][2] +
                mat_A[149][2] * mat_B[179][2] +
                mat_A[149][3] * mat_B[187][2] +
                mat_A[150][0] * mat_B[195][2] +
                mat_A[150][1] * mat_B[203][2] +
                mat_A[150][2] * mat_B[211][2] +
                mat_A[150][3] * mat_B[219][2] +
                mat_A[151][0] * mat_B[227][2] +
                mat_A[151][1] * mat_B[235][2] +
                mat_A[151][2] * mat_B[243][2] +
                mat_A[151][3] * mat_B[251][2];
    mat_C[147][3] <=
                mat_A[144][0] * mat_B[3][3] +
                mat_A[144][1] * mat_B[11][3] +
                mat_A[144][2] * mat_B[19][3] +
                mat_A[144][3] * mat_B[27][3] +
                mat_A[145][0] * mat_B[35][3] +
                mat_A[145][1] * mat_B[43][3] +
                mat_A[145][2] * mat_B[51][3] +
                mat_A[145][3] * mat_B[59][3] +
                mat_A[146][0] * mat_B[67][3] +
                mat_A[146][1] * mat_B[75][3] +
                mat_A[146][2] * mat_B[83][3] +
                mat_A[146][3] * mat_B[91][3] +
                mat_A[147][0] * mat_B[99][3] +
                mat_A[147][1] * mat_B[107][3] +
                mat_A[147][2] * mat_B[115][3] +
                mat_A[147][3] * mat_B[123][3] +
                mat_A[148][0] * mat_B[131][3] +
                mat_A[148][1] * mat_B[139][3] +
                mat_A[148][2] * mat_B[147][3] +
                mat_A[148][3] * mat_B[155][3] +
                mat_A[149][0] * mat_B[163][3] +
                mat_A[149][1] * mat_B[171][3] +
                mat_A[149][2] * mat_B[179][3] +
                mat_A[149][3] * mat_B[187][3] +
                mat_A[150][0] * mat_B[195][3] +
                mat_A[150][1] * mat_B[203][3] +
                mat_A[150][2] * mat_B[211][3] +
                mat_A[150][3] * mat_B[219][3] +
                mat_A[151][0] * mat_B[227][3] +
                mat_A[151][1] * mat_B[235][3] +
                mat_A[151][2] * mat_B[243][3] +
                mat_A[151][3] * mat_B[251][3];
    mat_C[148][0] <=
                mat_A[144][0] * mat_B[4][0] +
                mat_A[144][1] * mat_B[12][0] +
                mat_A[144][2] * mat_B[20][0] +
                mat_A[144][3] * mat_B[28][0] +
                mat_A[145][0] * mat_B[36][0] +
                mat_A[145][1] * mat_B[44][0] +
                mat_A[145][2] * mat_B[52][0] +
                mat_A[145][3] * mat_B[60][0] +
                mat_A[146][0] * mat_B[68][0] +
                mat_A[146][1] * mat_B[76][0] +
                mat_A[146][2] * mat_B[84][0] +
                mat_A[146][3] * mat_B[92][0] +
                mat_A[147][0] * mat_B[100][0] +
                mat_A[147][1] * mat_B[108][0] +
                mat_A[147][2] * mat_B[116][0] +
                mat_A[147][3] * mat_B[124][0] +
                mat_A[148][0] * mat_B[132][0] +
                mat_A[148][1] * mat_B[140][0] +
                mat_A[148][2] * mat_B[148][0] +
                mat_A[148][3] * mat_B[156][0] +
                mat_A[149][0] * mat_B[164][0] +
                mat_A[149][1] * mat_B[172][0] +
                mat_A[149][2] * mat_B[180][0] +
                mat_A[149][3] * mat_B[188][0] +
                mat_A[150][0] * mat_B[196][0] +
                mat_A[150][1] * mat_B[204][0] +
                mat_A[150][2] * mat_B[212][0] +
                mat_A[150][3] * mat_B[220][0] +
                mat_A[151][0] * mat_B[228][0] +
                mat_A[151][1] * mat_B[236][0] +
                mat_A[151][2] * mat_B[244][0] +
                mat_A[151][3] * mat_B[252][0];
    mat_C[148][1] <=
                mat_A[144][0] * mat_B[4][1] +
                mat_A[144][1] * mat_B[12][1] +
                mat_A[144][2] * mat_B[20][1] +
                mat_A[144][3] * mat_B[28][1] +
                mat_A[145][0] * mat_B[36][1] +
                mat_A[145][1] * mat_B[44][1] +
                mat_A[145][2] * mat_B[52][1] +
                mat_A[145][3] * mat_B[60][1] +
                mat_A[146][0] * mat_B[68][1] +
                mat_A[146][1] * mat_B[76][1] +
                mat_A[146][2] * mat_B[84][1] +
                mat_A[146][3] * mat_B[92][1] +
                mat_A[147][0] * mat_B[100][1] +
                mat_A[147][1] * mat_B[108][1] +
                mat_A[147][2] * mat_B[116][1] +
                mat_A[147][3] * mat_B[124][1] +
                mat_A[148][0] * mat_B[132][1] +
                mat_A[148][1] * mat_B[140][1] +
                mat_A[148][2] * mat_B[148][1] +
                mat_A[148][3] * mat_B[156][1] +
                mat_A[149][0] * mat_B[164][1] +
                mat_A[149][1] * mat_B[172][1] +
                mat_A[149][2] * mat_B[180][1] +
                mat_A[149][3] * mat_B[188][1] +
                mat_A[150][0] * mat_B[196][1] +
                mat_A[150][1] * mat_B[204][1] +
                mat_A[150][2] * mat_B[212][1] +
                mat_A[150][3] * mat_B[220][1] +
                mat_A[151][0] * mat_B[228][1] +
                mat_A[151][1] * mat_B[236][1] +
                mat_A[151][2] * mat_B[244][1] +
                mat_A[151][3] * mat_B[252][1];
    mat_C[148][2] <=
                mat_A[144][0] * mat_B[4][2] +
                mat_A[144][1] * mat_B[12][2] +
                mat_A[144][2] * mat_B[20][2] +
                mat_A[144][3] * mat_B[28][2] +
                mat_A[145][0] * mat_B[36][2] +
                mat_A[145][1] * mat_B[44][2] +
                mat_A[145][2] * mat_B[52][2] +
                mat_A[145][3] * mat_B[60][2] +
                mat_A[146][0] * mat_B[68][2] +
                mat_A[146][1] * mat_B[76][2] +
                mat_A[146][2] * mat_B[84][2] +
                mat_A[146][3] * mat_B[92][2] +
                mat_A[147][0] * mat_B[100][2] +
                mat_A[147][1] * mat_B[108][2] +
                mat_A[147][2] * mat_B[116][2] +
                mat_A[147][3] * mat_B[124][2] +
                mat_A[148][0] * mat_B[132][2] +
                mat_A[148][1] * mat_B[140][2] +
                mat_A[148][2] * mat_B[148][2] +
                mat_A[148][3] * mat_B[156][2] +
                mat_A[149][0] * mat_B[164][2] +
                mat_A[149][1] * mat_B[172][2] +
                mat_A[149][2] * mat_B[180][2] +
                mat_A[149][3] * mat_B[188][2] +
                mat_A[150][0] * mat_B[196][2] +
                mat_A[150][1] * mat_B[204][2] +
                mat_A[150][2] * mat_B[212][2] +
                mat_A[150][3] * mat_B[220][2] +
                mat_A[151][0] * mat_B[228][2] +
                mat_A[151][1] * mat_B[236][2] +
                mat_A[151][2] * mat_B[244][2] +
                mat_A[151][3] * mat_B[252][2];
    mat_C[148][3] <=
                mat_A[144][0] * mat_B[4][3] +
                mat_A[144][1] * mat_B[12][3] +
                mat_A[144][2] * mat_B[20][3] +
                mat_A[144][3] * mat_B[28][3] +
                mat_A[145][0] * mat_B[36][3] +
                mat_A[145][1] * mat_B[44][3] +
                mat_A[145][2] * mat_B[52][3] +
                mat_A[145][3] * mat_B[60][3] +
                mat_A[146][0] * mat_B[68][3] +
                mat_A[146][1] * mat_B[76][3] +
                mat_A[146][2] * mat_B[84][3] +
                mat_A[146][3] * mat_B[92][3] +
                mat_A[147][0] * mat_B[100][3] +
                mat_A[147][1] * mat_B[108][3] +
                mat_A[147][2] * mat_B[116][3] +
                mat_A[147][3] * mat_B[124][3] +
                mat_A[148][0] * mat_B[132][3] +
                mat_A[148][1] * mat_B[140][3] +
                mat_A[148][2] * mat_B[148][3] +
                mat_A[148][3] * mat_B[156][3] +
                mat_A[149][0] * mat_B[164][3] +
                mat_A[149][1] * mat_B[172][3] +
                mat_A[149][2] * mat_B[180][3] +
                mat_A[149][3] * mat_B[188][3] +
                mat_A[150][0] * mat_B[196][3] +
                mat_A[150][1] * mat_B[204][3] +
                mat_A[150][2] * mat_B[212][3] +
                mat_A[150][3] * mat_B[220][3] +
                mat_A[151][0] * mat_B[228][3] +
                mat_A[151][1] * mat_B[236][3] +
                mat_A[151][2] * mat_B[244][3] +
                mat_A[151][3] * mat_B[252][3];
    mat_C[149][0] <=
                mat_A[144][0] * mat_B[5][0] +
                mat_A[144][1] * mat_B[13][0] +
                mat_A[144][2] * mat_B[21][0] +
                mat_A[144][3] * mat_B[29][0] +
                mat_A[145][0] * mat_B[37][0] +
                mat_A[145][1] * mat_B[45][0] +
                mat_A[145][2] * mat_B[53][0] +
                mat_A[145][3] * mat_B[61][0] +
                mat_A[146][0] * mat_B[69][0] +
                mat_A[146][1] * mat_B[77][0] +
                mat_A[146][2] * mat_B[85][0] +
                mat_A[146][3] * mat_B[93][0] +
                mat_A[147][0] * mat_B[101][0] +
                mat_A[147][1] * mat_B[109][0] +
                mat_A[147][2] * mat_B[117][0] +
                mat_A[147][3] * mat_B[125][0] +
                mat_A[148][0] * mat_B[133][0] +
                mat_A[148][1] * mat_B[141][0] +
                mat_A[148][2] * mat_B[149][0] +
                mat_A[148][3] * mat_B[157][0] +
                mat_A[149][0] * mat_B[165][0] +
                mat_A[149][1] * mat_B[173][0] +
                mat_A[149][2] * mat_B[181][0] +
                mat_A[149][3] * mat_B[189][0] +
                mat_A[150][0] * mat_B[197][0] +
                mat_A[150][1] * mat_B[205][0] +
                mat_A[150][2] * mat_B[213][0] +
                mat_A[150][3] * mat_B[221][0] +
                mat_A[151][0] * mat_B[229][0] +
                mat_A[151][1] * mat_B[237][0] +
                mat_A[151][2] * mat_B[245][0] +
                mat_A[151][3] * mat_B[253][0];
    mat_C[149][1] <=
                mat_A[144][0] * mat_B[5][1] +
                mat_A[144][1] * mat_B[13][1] +
                mat_A[144][2] * mat_B[21][1] +
                mat_A[144][3] * mat_B[29][1] +
                mat_A[145][0] * mat_B[37][1] +
                mat_A[145][1] * mat_B[45][1] +
                mat_A[145][2] * mat_B[53][1] +
                mat_A[145][3] * mat_B[61][1] +
                mat_A[146][0] * mat_B[69][1] +
                mat_A[146][1] * mat_B[77][1] +
                mat_A[146][2] * mat_B[85][1] +
                mat_A[146][3] * mat_B[93][1] +
                mat_A[147][0] * mat_B[101][1] +
                mat_A[147][1] * mat_B[109][1] +
                mat_A[147][2] * mat_B[117][1] +
                mat_A[147][3] * mat_B[125][1] +
                mat_A[148][0] * mat_B[133][1] +
                mat_A[148][1] * mat_B[141][1] +
                mat_A[148][2] * mat_B[149][1] +
                mat_A[148][3] * mat_B[157][1] +
                mat_A[149][0] * mat_B[165][1] +
                mat_A[149][1] * mat_B[173][1] +
                mat_A[149][2] * mat_B[181][1] +
                mat_A[149][3] * mat_B[189][1] +
                mat_A[150][0] * mat_B[197][1] +
                mat_A[150][1] * mat_B[205][1] +
                mat_A[150][2] * mat_B[213][1] +
                mat_A[150][3] * mat_B[221][1] +
                mat_A[151][0] * mat_B[229][1] +
                mat_A[151][1] * mat_B[237][1] +
                mat_A[151][2] * mat_B[245][1] +
                mat_A[151][3] * mat_B[253][1];
    mat_C[149][2] <=
                mat_A[144][0] * mat_B[5][2] +
                mat_A[144][1] * mat_B[13][2] +
                mat_A[144][2] * mat_B[21][2] +
                mat_A[144][3] * mat_B[29][2] +
                mat_A[145][0] * mat_B[37][2] +
                mat_A[145][1] * mat_B[45][2] +
                mat_A[145][2] * mat_B[53][2] +
                mat_A[145][3] * mat_B[61][2] +
                mat_A[146][0] * mat_B[69][2] +
                mat_A[146][1] * mat_B[77][2] +
                mat_A[146][2] * mat_B[85][2] +
                mat_A[146][3] * mat_B[93][2] +
                mat_A[147][0] * mat_B[101][2] +
                mat_A[147][1] * mat_B[109][2] +
                mat_A[147][2] * mat_B[117][2] +
                mat_A[147][3] * mat_B[125][2] +
                mat_A[148][0] * mat_B[133][2] +
                mat_A[148][1] * mat_B[141][2] +
                mat_A[148][2] * mat_B[149][2] +
                mat_A[148][3] * mat_B[157][2] +
                mat_A[149][0] * mat_B[165][2] +
                mat_A[149][1] * mat_B[173][2] +
                mat_A[149][2] * mat_B[181][2] +
                mat_A[149][3] * mat_B[189][2] +
                mat_A[150][0] * mat_B[197][2] +
                mat_A[150][1] * mat_B[205][2] +
                mat_A[150][2] * mat_B[213][2] +
                mat_A[150][3] * mat_B[221][2] +
                mat_A[151][0] * mat_B[229][2] +
                mat_A[151][1] * mat_B[237][2] +
                mat_A[151][2] * mat_B[245][2] +
                mat_A[151][3] * mat_B[253][2];
    mat_C[149][3] <=
                mat_A[144][0] * mat_B[5][3] +
                mat_A[144][1] * mat_B[13][3] +
                mat_A[144][2] * mat_B[21][3] +
                mat_A[144][3] * mat_B[29][3] +
                mat_A[145][0] * mat_B[37][3] +
                mat_A[145][1] * mat_B[45][3] +
                mat_A[145][2] * mat_B[53][3] +
                mat_A[145][3] * mat_B[61][3] +
                mat_A[146][0] * mat_B[69][3] +
                mat_A[146][1] * mat_B[77][3] +
                mat_A[146][2] * mat_B[85][3] +
                mat_A[146][3] * mat_B[93][3] +
                mat_A[147][0] * mat_B[101][3] +
                mat_A[147][1] * mat_B[109][3] +
                mat_A[147][2] * mat_B[117][3] +
                mat_A[147][3] * mat_B[125][3] +
                mat_A[148][0] * mat_B[133][3] +
                mat_A[148][1] * mat_B[141][3] +
                mat_A[148][2] * mat_B[149][3] +
                mat_A[148][3] * mat_B[157][3] +
                mat_A[149][0] * mat_B[165][3] +
                mat_A[149][1] * mat_B[173][3] +
                mat_A[149][2] * mat_B[181][3] +
                mat_A[149][3] * mat_B[189][3] +
                mat_A[150][0] * mat_B[197][3] +
                mat_A[150][1] * mat_B[205][3] +
                mat_A[150][2] * mat_B[213][3] +
                mat_A[150][3] * mat_B[221][3] +
                mat_A[151][0] * mat_B[229][3] +
                mat_A[151][1] * mat_B[237][3] +
                mat_A[151][2] * mat_B[245][3] +
                mat_A[151][3] * mat_B[253][3];
    mat_C[150][0] <=
                mat_A[144][0] * mat_B[6][0] +
                mat_A[144][1] * mat_B[14][0] +
                mat_A[144][2] * mat_B[22][0] +
                mat_A[144][3] * mat_B[30][0] +
                mat_A[145][0] * mat_B[38][0] +
                mat_A[145][1] * mat_B[46][0] +
                mat_A[145][2] * mat_B[54][0] +
                mat_A[145][3] * mat_B[62][0] +
                mat_A[146][0] * mat_B[70][0] +
                mat_A[146][1] * mat_B[78][0] +
                mat_A[146][2] * mat_B[86][0] +
                mat_A[146][3] * mat_B[94][0] +
                mat_A[147][0] * mat_B[102][0] +
                mat_A[147][1] * mat_B[110][0] +
                mat_A[147][2] * mat_B[118][0] +
                mat_A[147][3] * mat_B[126][0] +
                mat_A[148][0] * mat_B[134][0] +
                mat_A[148][1] * mat_B[142][0] +
                mat_A[148][2] * mat_B[150][0] +
                mat_A[148][3] * mat_B[158][0] +
                mat_A[149][0] * mat_B[166][0] +
                mat_A[149][1] * mat_B[174][0] +
                mat_A[149][2] * mat_B[182][0] +
                mat_A[149][3] * mat_B[190][0] +
                mat_A[150][0] * mat_B[198][0] +
                mat_A[150][1] * mat_B[206][0] +
                mat_A[150][2] * mat_B[214][0] +
                mat_A[150][3] * mat_B[222][0] +
                mat_A[151][0] * mat_B[230][0] +
                mat_A[151][1] * mat_B[238][0] +
                mat_A[151][2] * mat_B[246][0] +
                mat_A[151][3] * mat_B[254][0];
    mat_C[150][1] <=
                mat_A[144][0] * mat_B[6][1] +
                mat_A[144][1] * mat_B[14][1] +
                mat_A[144][2] * mat_B[22][1] +
                mat_A[144][3] * mat_B[30][1] +
                mat_A[145][0] * mat_B[38][1] +
                mat_A[145][1] * mat_B[46][1] +
                mat_A[145][2] * mat_B[54][1] +
                mat_A[145][3] * mat_B[62][1] +
                mat_A[146][0] * mat_B[70][1] +
                mat_A[146][1] * mat_B[78][1] +
                mat_A[146][2] * mat_B[86][1] +
                mat_A[146][3] * mat_B[94][1] +
                mat_A[147][0] * mat_B[102][1] +
                mat_A[147][1] * mat_B[110][1] +
                mat_A[147][2] * mat_B[118][1] +
                mat_A[147][3] * mat_B[126][1] +
                mat_A[148][0] * mat_B[134][1] +
                mat_A[148][1] * mat_B[142][1] +
                mat_A[148][2] * mat_B[150][1] +
                mat_A[148][3] * mat_B[158][1] +
                mat_A[149][0] * mat_B[166][1] +
                mat_A[149][1] * mat_B[174][1] +
                mat_A[149][2] * mat_B[182][1] +
                mat_A[149][3] * mat_B[190][1] +
                mat_A[150][0] * mat_B[198][1] +
                mat_A[150][1] * mat_B[206][1] +
                mat_A[150][2] * mat_B[214][1] +
                mat_A[150][3] * mat_B[222][1] +
                mat_A[151][0] * mat_B[230][1] +
                mat_A[151][1] * mat_B[238][1] +
                mat_A[151][2] * mat_B[246][1] +
                mat_A[151][3] * mat_B[254][1];
    mat_C[150][2] <=
                mat_A[144][0] * mat_B[6][2] +
                mat_A[144][1] * mat_B[14][2] +
                mat_A[144][2] * mat_B[22][2] +
                mat_A[144][3] * mat_B[30][2] +
                mat_A[145][0] * mat_B[38][2] +
                mat_A[145][1] * mat_B[46][2] +
                mat_A[145][2] * mat_B[54][2] +
                mat_A[145][3] * mat_B[62][2] +
                mat_A[146][0] * mat_B[70][2] +
                mat_A[146][1] * mat_B[78][2] +
                mat_A[146][2] * mat_B[86][2] +
                mat_A[146][3] * mat_B[94][2] +
                mat_A[147][0] * mat_B[102][2] +
                mat_A[147][1] * mat_B[110][2] +
                mat_A[147][2] * mat_B[118][2] +
                mat_A[147][3] * mat_B[126][2] +
                mat_A[148][0] * mat_B[134][2] +
                mat_A[148][1] * mat_B[142][2] +
                mat_A[148][2] * mat_B[150][2] +
                mat_A[148][3] * mat_B[158][2] +
                mat_A[149][0] * mat_B[166][2] +
                mat_A[149][1] * mat_B[174][2] +
                mat_A[149][2] * mat_B[182][2] +
                mat_A[149][3] * mat_B[190][2] +
                mat_A[150][0] * mat_B[198][2] +
                mat_A[150][1] * mat_B[206][2] +
                mat_A[150][2] * mat_B[214][2] +
                mat_A[150][3] * mat_B[222][2] +
                mat_A[151][0] * mat_B[230][2] +
                mat_A[151][1] * mat_B[238][2] +
                mat_A[151][2] * mat_B[246][2] +
                mat_A[151][3] * mat_B[254][2];
    mat_C[150][3] <=
                mat_A[144][0] * mat_B[6][3] +
                mat_A[144][1] * mat_B[14][3] +
                mat_A[144][2] * mat_B[22][3] +
                mat_A[144][3] * mat_B[30][3] +
                mat_A[145][0] * mat_B[38][3] +
                mat_A[145][1] * mat_B[46][3] +
                mat_A[145][2] * mat_B[54][3] +
                mat_A[145][3] * mat_B[62][3] +
                mat_A[146][0] * mat_B[70][3] +
                mat_A[146][1] * mat_B[78][3] +
                mat_A[146][2] * mat_B[86][3] +
                mat_A[146][3] * mat_B[94][3] +
                mat_A[147][0] * mat_B[102][3] +
                mat_A[147][1] * mat_B[110][3] +
                mat_A[147][2] * mat_B[118][3] +
                mat_A[147][3] * mat_B[126][3] +
                mat_A[148][0] * mat_B[134][3] +
                mat_A[148][1] * mat_B[142][3] +
                mat_A[148][2] * mat_B[150][3] +
                mat_A[148][3] * mat_B[158][3] +
                mat_A[149][0] * mat_B[166][3] +
                mat_A[149][1] * mat_B[174][3] +
                mat_A[149][2] * mat_B[182][3] +
                mat_A[149][3] * mat_B[190][3] +
                mat_A[150][0] * mat_B[198][3] +
                mat_A[150][1] * mat_B[206][3] +
                mat_A[150][2] * mat_B[214][3] +
                mat_A[150][3] * mat_B[222][3] +
                mat_A[151][0] * mat_B[230][3] +
                mat_A[151][1] * mat_B[238][3] +
                mat_A[151][2] * mat_B[246][3] +
                mat_A[151][3] * mat_B[254][3];
    mat_C[151][0] <=
                mat_A[144][0] * mat_B[7][0] +
                mat_A[144][1] * mat_B[15][0] +
                mat_A[144][2] * mat_B[23][0] +
                mat_A[144][3] * mat_B[31][0] +
                mat_A[145][0] * mat_B[39][0] +
                mat_A[145][1] * mat_B[47][0] +
                mat_A[145][2] * mat_B[55][0] +
                mat_A[145][3] * mat_B[63][0] +
                mat_A[146][0] * mat_B[71][0] +
                mat_A[146][1] * mat_B[79][0] +
                mat_A[146][2] * mat_B[87][0] +
                mat_A[146][3] * mat_B[95][0] +
                mat_A[147][0] * mat_B[103][0] +
                mat_A[147][1] * mat_B[111][0] +
                mat_A[147][2] * mat_B[119][0] +
                mat_A[147][3] * mat_B[127][0] +
                mat_A[148][0] * mat_B[135][0] +
                mat_A[148][1] * mat_B[143][0] +
                mat_A[148][2] * mat_B[151][0] +
                mat_A[148][3] * mat_B[159][0] +
                mat_A[149][0] * mat_B[167][0] +
                mat_A[149][1] * mat_B[175][0] +
                mat_A[149][2] * mat_B[183][0] +
                mat_A[149][3] * mat_B[191][0] +
                mat_A[150][0] * mat_B[199][0] +
                mat_A[150][1] * mat_B[207][0] +
                mat_A[150][2] * mat_B[215][0] +
                mat_A[150][3] * mat_B[223][0] +
                mat_A[151][0] * mat_B[231][0] +
                mat_A[151][1] * mat_B[239][0] +
                mat_A[151][2] * mat_B[247][0] +
                mat_A[151][3] * mat_B[255][0];
    mat_C[151][1] <=
                mat_A[144][0] * mat_B[7][1] +
                mat_A[144][1] * mat_B[15][1] +
                mat_A[144][2] * mat_B[23][1] +
                mat_A[144][3] * mat_B[31][1] +
                mat_A[145][0] * mat_B[39][1] +
                mat_A[145][1] * mat_B[47][1] +
                mat_A[145][2] * mat_B[55][1] +
                mat_A[145][3] * mat_B[63][1] +
                mat_A[146][0] * mat_B[71][1] +
                mat_A[146][1] * mat_B[79][1] +
                mat_A[146][2] * mat_B[87][1] +
                mat_A[146][3] * mat_B[95][1] +
                mat_A[147][0] * mat_B[103][1] +
                mat_A[147][1] * mat_B[111][1] +
                mat_A[147][2] * mat_B[119][1] +
                mat_A[147][3] * mat_B[127][1] +
                mat_A[148][0] * mat_B[135][1] +
                mat_A[148][1] * mat_B[143][1] +
                mat_A[148][2] * mat_B[151][1] +
                mat_A[148][3] * mat_B[159][1] +
                mat_A[149][0] * mat_B[167][1] +
                mat_A[149][1] * mat_B[175][1] +
                mat_A[149][2] * mat_B[183][1] +
                mat_A[149][3] * mat_B[191][1] +
                mat_A[150][0] * mat_B[199][1] +
                mat_A[150][1] * mat_B[207][1] +
                mat_A[150][2] * mat_B[215][1] +
                mat_A[150][3] * mat_B[223][1] +
                mat_A[151][0] * mat_B[231][1] +
                mat_A[151][1] * mat_B[239][1] +
                mat_A[151][2] * mat_B[247][1] +
                mat_A[151][3] * mat_B[255][1];
    mat_C[151][2] <=
                mat_A[144][0] * mat_B[7][2] +
                mat_A[144][1] * mat_B[15][2] +
                mat_A[144][2] * mat_B[23][2] +
                mat_A[144][3] * mat_B[31][2] +
                mat_A[145][0] * mat_B[39][2] +
                mat_A[145][1] * mat_B[47][2] +
                mat_A[145][2] * mat_B[55][2] +
                mat_A[145][3] * mat_B[63][2] +
                mat_A[146][0] * mat_B[71][2] +
                mat_A[146][1] * mat_B[79][2] +
                mat_A[146][2] * mat_B[87][2] +
                mat_A[146][3] * mat_B[95][2] +
                mat_A[147][0] * mat_B[103][2] +
                mat_A[147][1] * mat_B[111][2] +
                mat_A[147][2] * mat_B[119][2] +
                mat_A[147][3] * mat_B[127][2] +
                mat_A[148][0] * mat_B[135][2] +
                mat_A[148][1] * mat_B[143][2] +
                mat_A[148][2] * mat_B[151][2] +
                mat_A[148][3] * mat_B[159][2] +
                mat_A[149][0] * mat_B[167][2] +
                mat_A[149][1] * mat_B[175][2] +
                mat_A[149][2] * mat_B[183][2] +
                mat_A[149][3] * mat_B[191][2] +
                mat_A[150][0] * mat_B[199][2] +
                mat_A[150][1] * mat_B[207][2] +
                mat_A[150][2] * mat_B[215][2] +
                mat_A[150][3] * mat_B[223][2] +
                mat_A[151][0] * mat_B[231][2] +
                mat_A[151][1] * mat_B[239][2] +
                mat_A[151][2] * mat_B[247][2] +
                mat_A[151][3] * mat_B[255][2];
    mat_C[151][3] <=
                mat_A[144][0] * mat_B[7][3] +
                mat_A[144][1] * mat_B[15][3] +
                mat_A[144][2] * mat_B[23][3] +
                mat_A[144][3] * mat_B[31][3] +
                mat_A[145][0] * mat_B[39][3] +
                mat_A[145][1] * mat_B[47][3] +
                mat_A[145][2] * mat_B[55][3] +
                mat_A[145][3] * mat_B[63][3] +
                mat_A[146][0] * mat_B[71][3] +
                mat_A[146][1] * mat_B[79][3] +
                mat_A[146][2] * mat_B[87][3] +
                mat_A[146][3] * mat_B[95][3] +
                mat_A[147][0] * mat_B[103][3] +
                mat_A[147][1] * mat_B[111][3] +
                mat_A[147][2] * mat_B[119][3] +
                mat_A[147][3] * mat_B[127][3] +
                mat_A[148][0] * mat_B[135][3] +
                mat_A[148][1] * mat_B[143][3] +
                mat_A[148][2] * mat_B[151][3] +
                mat_A[148][3] * mat_B[159][3] +
                mat_A[149][0] * mat_B[167][3] +
                mat_A[149][1] * mat_B[175][3] +
                mat_A[149][2] * mat_B[183][3] +
                mat_A[149][3] * mat_B[191][3] +
                mat_A[150][0] * mat_B[199][3] +
                mat_A[150][1] * mat_B[207][3] +
                mat_A[150][2] * mat_B[215][3] +
                mat_A[150][3] * mat_B[223][3] +
                mat_A[151][0] * mat_B[231][3] +
                mat_A[151][1] * mat_B[239][3] +
                mat_A[151][2] * mat_B[247][3] +
                mat_A[151][3] * mat_B[255][3];
    mat_C[152][0] <=
                mat_A[152][0] * mat_B[0][0] +
                mat_A[152][1] * mat_B[8][0] +
                mat_A[152][2] * mat_B[16][0] +
                mat_A[152][3] * mat_B[24][0] +
                mat_A[153][0] * mat_B[32][0] +
                mat_A[153][1] * mat_B[40][0] +
                mat_A[153][2] * mat_B[48][0] +
                mat_A[153][3] * mat_B[56][0] +
                mat_A[154][0] * mat_B[64][0] +
                mat_A[154][1] * mat_B[72][0] +
                mat_A[154][2] * mat_B[80][0] +
                mat_A[154][3] * mat_B[88][0] +
                mat_A[155][0] * mat_B[96][0] +
                mat_A[155][1] * mat_B[104][0] +
                mat_A[155][2] * mat_B[112][0] +
                mat_A[155][3] * mat_B[120][0] +
                mat_A[156][0] * mat_B[128][0] +
                mat_A[156][1] * mat_B[136][0] +
                mat_A[156][2] * mat_B[144][0] +
                mat_A[156][3] * mat_B[152][0] +
                mat_A[157][0] * mat_B[160][0] +
                mat_A[157][1] * mat_B[168][0] +
                mat_A[157][2] * mat_B[176][0] +
                mat_A[157][3] * mat_B[184][0] +
                mat_A[158][0] * mat_B[192][0] +
                mat_A[158][1] * mat_B[200][0] +
                mat_A[158][2] * mat_B[208][0] +
                mat_A[158][3] * mat_B[216][0] +
                mat_A[159][0] * mat_B[224][0] +
                mat_A[159][1] * mat_B[232][0] +
                mat_A[159][2] * mat_B[240][0] +
                mat_A[159][3] * mat_B[248][0];
    mat_C[152][1] <=
                mat_A[152][0] * mat_B[0][1] +
                mat_A[152][1] * mat_B[8][1] +
                mat_A[152][2] * mat_B[16][1] +
                mat_A[152][3] * mat_B[24][1] +
                mat_A[153][0] * mat_B[32][1] +
                mat_A[153][1] * mat_B[40][1] +
                mat_A[153][2] * mat_B[48][1] +
                mat_A[153][3] * mat_B[56][1] +
                mat_A[154][0] * mat_B[64][1] +
                mat_A[154][1] * mat_B[72][1] +
                mat_A[154][2] * mat_B[80][1] +
                mat_A[154][3] * mat_B[88][1] +
                mat_A[155][0] * mat_B[96][1] +
                mat_A[155][1] * mat_B[104][1] +
                mat_A[155][2] * mat_B[112][1] +
                mat_A[155][3] * mat_B[120][1] +
                mat_A[156][0] * mat_B[128][1] +
                mat_A[156][1] * mat_B[136][1] +
                mat_A[156][2] * mat_B[144][1] +
                mat_A[156][3] * mat_B[152][1] +
                mat_A[157][0] * mat_B[160][1] +
                mat_A[157][1] * mat_B[168][1] +
                mat_A[157][2] * mat_B[176][1] +
                mat_A[157][3] * mat_B[184][1] +
                mat_A[158][0] * mat_B[192][1] +
                mat_A[158][1] * mat_B[200][1] +
                mat_A[158][2] * mat_B[208][1] +
                mat_A[158][3] * mat_B[216][1] +
                mat_A[159][0] * mat_B[224][1] +
                mat_A[159][1] * mat_B[232][1] +
                mat_A[159][2] * mat_B[240][1] +
                mat_A[159][3] * mat_B[248][1];
    mat_C[152][2] <=
                mat_A[152][0] * mat_B[0][2] +
                mat_A[152][1] * mat_B[8][2] +
                mat_A[152][2] * mat_B[16][2] +
                mat_A[152][3] * mat_B[24][2] +
                mat_A[153][0] * mat_B[32][2] +
                mat_A[153][1] * mat_B[40][2] +
                mat_A[153][2] * mat_B[48][2] +
                mat_A[153][3] * mat_B[56][2] +
                mat_A[154][0] * mat_B[64][2] +
                mat_A[154][1] * mat_B[72][2] +
                mat_A[154][2] * mat_B[80][2] +
                mat_A[154][3] * mat_B[88][2] +
                mat_A[155][0] * mat_B[96][2] +
                mat_A[155][1] * mat_B[104][2] +
                mat_A[155][2] * mat_B[112][2] +
                mat_A[155][3] * mat_B[120][2] +
                mat_A[156][0] * mat_B[128][2] +
                mat_A[156][1] * mat_B[136][2] +
                mat_A[156][2] * mat_B[144][2] +
                mat_A[156][3] * mat_B[152][2] +
                mat_A[157][0] * mat_B[160][2] +
                mat_A[157][1] * mat_B[168][2] +
                mat_A[157][2] * mat_B[176][2] +
                mat_A[157][3] * mat_B[184][2] +
                mat_A[158][0] * mat_B[192][2] +
                mat_A[158][1] * mat_B[200][2] +
                mat_A[158][2] * mat_B[208][2] +
                mat_A[158][3] * mat_B[216][2] +
                mat_A[159][0] * mat_B[224][2] +
                mat_A[159][1] * mat_B[232][2] +
                mat_A[159][2] * mat_B[240][2] +
                mat_A[159][3] * mat_B[248][2];
    mat_C[152][3] <=
                mat_A[152][0] * mat_B[0][3] +
                mat_A[152][1] * mat_B[8][3] +
                mat_A[152][2] * mat_B[16][3] +
                mat_A[152][3] * mat_B[24][3] +
                mat_A[153][0] * mat_B[32][3] +
                mat_A[153][1] * mat_B[40][3] +
                mat_A[153][2] * mat_B[48][3] +
                mat_A[153][3] * mat_B[56][3] +
                mat_A[154][0] * mat_B[64][3] +
                mat_A[154][1] * mat_B[72][3] +
                mat_A[154][2] * mat_B[80][3] +
                mat_A[154][3] * mat_B[88][3] +
                mat_A[155][0] * mat_B[96][3] +
                mat_A[155][1] * mat_B[104][3] +
                mat_A[155][2] * mat_B[112][3] +
                mat_A[155][3] * mat_B[120][3] +
                mat_A[156][0] * mat_B[128][3] +
                mat_A[156][1] * mat_B[136][3] +
                mat_A[156][2] * mat_B[144][3] +
                mat_A[156][3] * mat_B[152][3] +
                mat_A[157][0] * mat_B[160][3] +
                mat_A[157][1] * mat_B[168][3] +
                mat_A[157][2] * mat_B[176][3] +
                mat_A[157][3] * mat_B[184][3] +
                mat_A[158][0] * mat_B[192][3] +
                mat_A[158][1] * mat_B[200][3] +
                mat_A[158][2] * mat_B[208][3] +
                mat_A[158][3] * mat_B[216][3] +
                mat_A[159][0] * mat_B[224][3] +
                mat_A[159][1] * mat_B[232][3] +
                mat_A[159][2] * mat_B[240][3] +
                mat_A[159][3] * mat_B[248][3];
    mat_C[153][0] <=
                mat_A[152][0] * mat_B[1][0] +
                mat_A[152][1] * mat_B[9][0] +
                mat_A[152][2] * mat_B[17][0] +
                mat_A[152][3] * mat_B[25][0] +
                mat_A[153][0] * mat_B[33][0] +
                mat_A[153][1] * mat_B[41][0] +
                mat_A[153][2] * mat_B[49][0] +
                mat_A[153][3] * mat_B[57][0] +
                mat_A[154][0] * mat_B[65][0] +
                mat_A[154][1] * mat_B[73][0] +
                mat_A[154][2] * mat_B[81][0] +
                mat_A[154][3] * mat_B[89][0] +
                mat_A[155][0] * mat_B[97][0] +
                mat_A[155][1] * mat_B[105][0] +
                mat_A[155][2] * mat_B[113][0] +
                mat_A[155][3] * mat_B[121][0] +
                mat_A[156][0] * mat_B[129][0] +
                mat_A[156][1] * mat_B[137][0] +
                mat_A[156][2] * mat_B[145][0] +
                mat_A[156][3] * mat_B[153][0] +
                mat_A[157][0] * mat_B[161][0] +
                mat_A[157][1] * mat_B[169][0] +
                mat_A[157][2] * mat_B[177][0] +
                mat_A[157][3] * mat_B[185][0] +
                mat_A[158][0] * mat_B[193][0] +
                mat_A[158][1] * mat_B[201][0] +
                mat_A[158][2] * mat_B[209][0] +
                mat_A[158][3] * mat_B[217][0] +
                mat_A[159][0] * mat_B[225][0] +
                mat_A[159][1] * mat_B[233][0] +
                mat_A[159][2] * mat_B[241][0] +
                mat_A[159][3] * mat_B[249][0];
    mat_C[153][1] <=
                mat_A[152][0] * mat_B[1][1] +
                mat_A[152][1] * mat_B[9][1] +
                mat_A[152][2] * mat_B[17][1] +
                mat_A[152][3] * mat_B[25][1] +
                mat_A[153][0] * mat_B[33][1] +
                mat_A[153][1] * mat_B[41][1] +
                mat_A[153][2] * mat_B[49][1] +
                mat_A[153][3] * mat_B[57][1] +
                mat_A[154][0] * mat_B[65][1] +
                mat_A[154][1] * mat_B[73][1] +
                mat_A[154][2] * mat_B[81][1] +
                mat_A[154][3] * mat_B[89][1] +
                mat_A[155][0] * mat_B[97][1] +
                mat_A[155][1] * mat_B[105][1] +
                mat_A[155][2] * mat_B[113][1] +
                mat_A[155][3] * mat_B[121][1] +
                mat_A[156][0] * mat_B[129][1] +
                mat_A[156][1] * mat_B[137][1] +
                mat_A[156][2] * mat_B[145][1] +
                mat_A[156][3] * mat_B[153][1] +
                mat_A[157][0] * mat_B[161][1] +
                mat_A[157][1] * mat_B[169][1] +
                mat_A[157][2] * mat_B[177][1] +
                mat_A[157][3] * mat_B[185][1] +
                mat_A[158][0] * mat_B[193][1] +
                mat_A[158][1] * mat_B[201][1] +
                mat_A[158][2] * mat_B[209][1] +
                mat_A[158][3] * mat_B[217][1] +
                mat_A[159][0] * mat_B[225][1] +
                mat_A[159][1] * mat_B[233][1] +
                mat_A[159][2] * mat_B[241][1] +
                mat_A[159][3] * mat_B[249][1];
    mat_C[153][2] <=
                mat_A[152][0] * mat_B[1][2] +
                mat_A[152][1] * mat_B[9][2] +
                mat_A[152][2] * mat_B[17][2] +
                mat_A[152][3] * mat_B[25][2] +
                mat_A[153][0] * mat_B[33][2] +
                mat_A[153][1] * mat_B[41][2] +
                mat_A[153][2] * mat_B[49][2] +
                mat_A[153][3] * mat_B[57][2] +
                mat_A[154][0] * mat_B[65][2] +
                mat_A[154][1] * mat_B[73][2] +
                mat_A[154][2] * mat_B[81][2] +
                mat_A[154][3] * mat_B[89][2] +
                mat_A[155][0] * mat_B[97][2] +
                mat_A[155][1] * mat_B[105][2] +
                mat_A[155][2] * mat_B[113][2] +
                mat_A[155][3] * mat_B[121][2] +
                mat_A[156][0] * mat_B[129][2] +
                mat_A[156][1] * mat_B[137][2] +
                mat_A[156][2] * mat_B[145][2] +
                mat_A[156][3] * mat_B[153][2] +
                mat_A[157][0] * mat_B[161][2] +
                mat_A[157][1] * mat_B[169][2] +
                mat_A[157][2] * mat_B[177][2] +
                mat_A[157][3] * mat_B[185][2] +
                mat_A[158][0] * mat_B[193][2] +
                mat_A[158][1] * mat_B[201][2] +
                mat_A[158][2] * mat_B[209][2] +
                mat_A[158][3] * mat_B[217][2] +
                mat_A[159][0] * mat_B[225][2] +
                mat_A[159][1] * mat_B[233][2] +
                mat_A[159][2] * mat_B[241][2] +
                mat_A[159][3] * mat_B[249][2];
    mat_C[153][3] <=
                mat_A[152][0] * mat_B[1][3] +
                mat_A[152][1] * mat_B[9][3] +
                mat_A[152][2] * mat_B[17][3] +
                mat_A[152][3] * mat_B[25][3] +
                mat_A[153][0] * mat_B[33][3] +
                mat_A[153][1] * mat_B[41][3] +
                mat_A[153][2] * mat_B[49][3] +
                mat_A[153][3] * mat_B[57][3] +
                mat_A[154][0] * mat_B[65][3] +
                mat_A[154][1] * mat_B[73][3] +
                mat_A[154][2] * mat_B[81][3] +
                mat_A[154][3] * mat_B[89][3] +
                mat_A[155][0] * mat_B[97][3] +
                mat_A[155][1] * mat_B[105][3] +
                mat_A[155][2] * mat_B[113][3] +
                mat_A[155][3] * mat_B[121][3] +
                mat_A[156][0] * mat_B[129][3] +
                mat_A[156][1] * mat_B[137][3] +
                mat_A[156][2] * mat_B[145][3] +
                mat_A[156][3] * mat_B[153][3] +
                mat_A[157][0] * mat_B[161][3] +
                mat_A[157][1] * mat_B[169][3] +
                mat_A[157][2] * mat_B[177][3] +
                mat_A[157][3] * mat_B[185][3] +
                mat_A[158][0] * mat_B[193][3] +
                mat_A[158][1] * mat_B[201][3] +
                mat_A[158][2] * mat_B[209][3] +
                mat_A[158][3] * mat_B[217][3] +
                mat_A[159][0] * mat_B[225][3] +
                mat_A[159][1] * mat_B[233][3] +
                mat_A[159][2] * mat_B[241][3] +
                mat_A[159][3] * mat_B[249][3];
    mat_C[154][0] <=
                mat_A[152][0] * mat_B[2][0] +
                mat_A[152][1] * mat_B[10][0] +
                mat_A[152][2] * mat_B[18][0] +
                mat_A[152][3] * mat_B[26][0] +
                mat_A[153][0] * mat_B[34][0] +
                mat_A[153][1] * mat_B[42][0] +
                mat_A[153][2] * mat_B[50][0] +
                mat_A[153][3] * mat_B[58][0] +
                mat_A[154][0] * mat_B[66][0] +
                mat_A[154][1] * mat_B[74][0] +
                mat_A[154][2] * mat_B[82][0] +
                mat_A[154][3] * mat_B[90][0] +
                mat_A[155][0] * mat_B[98][0] +
                mat_A[155][1] * mat_B[106][0] +
                mat_A[155][2] * mat_B[114][0] +
                mat_A[155][3] * mat_B[122][0] +
                mat_A[156][0] * mat_B[130][0] +
                mat_A[156][1] * mat_B[138][0] +
                mat_A[156][2] * mat_B[146][0] +
                mat_A[156][3] * mat_B[154][0] +
                mat_A[157][0] * mat_B[162][0] +
                mat_A[157][1] * mat_B[170][0] +
                mat_A[157][2] * mat_B[178][0] +
                mat_A[157][3] * mat_B[186][0] +
                mat_A[158][0] * mat_B[194][0] +
                mat_A[158][1] * mat_B[202][0] +
                mat_A[158][2] * mat_B[210][0] +
                mat_A[158][3] * mat_B[218][0] +
                mat_A[159][0] * mat_B[226][0] +
                mat_A[159][1] * mat_B[234][0] +
                mat_A[159][2] * mat_B[242][0] +
                mat_A[159][3] * mat_B[250][0];
    mat_C[154][1] <=
                mat_A[152][0] * mat_B[2][1] +
                mat_A[152][1] * mat_B[10][1] +
                mat_A[152][2] * mat_B[18][1] +
                mat_A[152][3] * mat_B[26][1] +
                mat_A[153][0] * mat_B[34][1] +
                mat_A[153][1] * mat_B[42][1] +
                mat_A[153][2] * mat_B[50][1] +
                mat_A[153][3] * mat_B[58][1] +
                mat_A[154][0] * mat_B[66][1] +
                mat_A[154][1] * mat_B[74][1] +
                mat_A[154][2] * mat_B[82][1] +
                mat_A[154][3] * mat_B[90][1] +
                mat_A[155][0] * mat_B[98][1] +
                mat_A[155][1] * mat_B[106][1] +
                mat_A[155][2] * mat_B[114][1] +
                mat_A[155][3] * mat_B[122][1] +
                mat_A[156][0] * mat_B[130][1] +
                mat_A[156][1] * mat_B[138][1] +
                mat_A[156][2] * mat_B[146][1] +
                mat_A[156][3] * mat_B[154][1] +
                mat_A[157][0] * mat_B[162][1] +
                mat_A[157][1] * mat_B[170][1] +
                mat_A[157][2] * mat_B[178][1] +
                mat_A[157][3] * mat_B[186][1] +
                mat_A[158][0] * mat_B[194][1] +
                mat_A[158][1] * mat_B[202][1] +
                mat_A[158][2] * mat_B[210][1] +
                mat_A[158][3] * mat_B[218][1] +
                mat_A[159][0] * mat_B[226][1] +
                mat_A[159][1] * mat_B[234][1] +
                mat_A[159][2] * mat_B[242][1] +
                mat_A[159][3] * mat_B[250][1];
    mat_C[154][2] <=
                mat_A[152][0] * mat_B[2][2] +
                mat_A[152][1] * mat_B[10][2] +
                mat_A[152][2] * mat_B[18][2] +
                mat_A[152][3] * mat_B[26][2] +
                mat_A[153][0] * mat_B[34][2] +
                mat_A[153][1] * mat_B[42][2] +
                mat_A[153][2] * mat_B[50][2] +
                mat_A[153][3] * mat_B[58][2] +
                mat_A[154][0] * mat_B[66][2] +
                mat_A[154][1] * mat_B[74][2] +
                mat_A[154][2] * mat_B[82][2] +
                mat_A[154][3] * mat_B[90][2] +
                mat_A[155][0] * mat_B[98][2] +
                mat_A[155][1] * mat_B[106][2] +
                mat_A[155][2] * mat_B[114][2] +
                mat_A[155][3] * mat_B[122][2] +
                mat_A[156][0] * mat_B[130][2] +
                mat_A[156][1] * mat_B[138][2] +
                mat_A[156][2] * mat_B[146][2] +
                mat_A[156][3] * mat_B[154][2] +
                mat_A[157][0] * mat_B[162][2] +
                mat_A[157][1] * mat_B[170][2] +
                mat_A[157][2] * mat_B[178][2] +
                mat_A[157][3] * mat_B[186][2] +
                mat_A[158][0] * mat_B[194][2] +
                mat_A[158][1] * mat_B[202][2] +
                mat_A[158][2] * mat_B[210][2] +
                mat_A[158][3] * mat_B[218][2] +
                mat_A[159][0] * mat_B[226][2] +
                mat_A[159][1] * mat_B[234][2] +
                mat_A[159][2] * mat_B[242][2] +
                mat_A[159][3] * mat_B[250][2];
    mat_C[154][3] <=
                mat_A[152][0] * mat_B[2][3] +
                mat_A[152][1] * mat_B[10][3] +
                mat_A[152][2] * mat_B[18][3] +
                mat_A[152][3] * mat_B[26][3] +
                mat_A[153][0] * mat_B[34][3] +
                mat_A[153][1] * mat_B[42][3] +
                mat_A[153][2] * mat_B[50][3] +
                mat_A[153][3] * mat_B[58][3] +
                mat_A[154][0] * mat_B[66][3] +
                mat_A[154][1] * mat_B[74][3] +
                mat_A[154][2] * mat_B[82][3] +
                mat_A[154][3] * mat_B[90][3] +
                mat_A[155][0] * mat_B[98][3] +
                mat_A[155][1] * mat_B[106][3] +
                mat_A[155][2] * mat_B[114][3] +
                mat_A[155][3] * mat_B[122][3] +
                mat_A[156][0] * mat_B[130][3] +
                mat_A[156][1] * mat_B[138][3] +
                mat_A[156][2] * mat_B[146][3] +
                mat_A[156][3] * mat_B[154][3] +
                mat_A[157][0] * mat_B[162][3] +
                mat_A[157][1] * mat_B[170][3] +
                mat_A[157][2] * mat_B[178][3] +
                mat_A[157][3] * mat_B[186][3] +
                mat_A[158][0] * mat_B[194][3] +
                mat_A[158][1] * mat_B[202][3] +
                mat_A[158][2] * mat_B[210][3] +
                mat_A[158][3] * mat_B[218][3] +
                mat_A[159][0] * mat_B[226][3] +
                mat_A[159][1] * mat_B[234][3] +
                mat_A[159][2] * mat_B[242][3] +
                mat_A[159][3] * mat_B[250][3];
    mat_C[155][0] <=
                mat_A[152][0] * mat_B[3][0] +
                mat_A[152][1] * mat_B[11][0] +
                mat_A[152][2] * mat_B[19][0] +
                mat_A[152][3] * mat_B[27][0] +
                mat_A[153][0] * mat_B[35][0] +
                mat_A[153][1] * mat_B[43][0] +
                mat_A[153][2] * mat_B[51][0] +
                mat_A[153][3] * mat_B[59][0] +
                mat_A[154][0] * mat_B[67][0] +
                mat_A[154][1] * mat_B[75][0] +
                mat_A[154][2] * mat_B[83][0] +
                mat_A[154][3] * mat_B[91][0] +
                mat_A[155][0] * mat_B[99][0] +
                mat_A[155][1] * mat_B[107][0] +
                mat_A[155][2] * mat_B[115][0] +
                mat_A[155][3] * mat_B[123][0] +
                mat_A[156][0] * mat_B[131][0] +
                mat_A[156][1] * mat_B[139][0] +
                mat_A[156][2] * mat_B[147][0] +
                mat_A[156][3] * mat_B[155][0] +
                mat_A[157][0] * mat_B[163][0] +
                mat_A[157][1] * mat_B[171][0] +
                mat_A[157][2] * mat_B[179][0] +
                mat_A[157][3] * mat_B[187][0] +
                mat_A[158][0] * mat_B[195][0] +
                mat_A[158][1] * mat_B[203][0] +
                mat_A[158][2] * mat_B[211][0] +
                mat_A[158][3] * mat_B[219][0] +
                mat_A[159][0] * mat_B[227][0] +
                mat_A[159][1] * mat_B[235][0] +
                mat_A[159][2] * mat_B[243][0] +
                mat_A[159][3] * mat_B[251][0];
    mat_C[155][1] <=
                mat_A[152][0] * mat_B[3][1] +
                mat_A[152][1] * mat_B[11][1] +
                mat_A[152][2] * mat_B[19][1] +
                mat_A[152][3] * mat_B[27][1] +
                mat_A[153][0] * mat_B[35][1] +
                mat_A[153][1] * mat_B[43][1] +
                mat_A[153][2] * mat_B[51][1] +
                mat_A[153][3] * mat_B[59][1] +
                mat_A[154][0] * mat_B[67][1] +
                mat_A[154][1] * mat_B[75][1] +
                mat_A[154][2] * mat_B[83][1] +
                mat_A[154][3] * mat_B[91][1] +
                mat_A[155][0] * mat_B[99][1] +
                mat_A[155][1] * mat_B[107][1] +
                mat_A[155][2] * mat_B[115][1] +
                mat_A[155][3] * mat_B[123][1] +
                mat_A[156][0] * mat_B[131][1] +
                mat_A[156][1] * mat_B[139][1] +
                mat_A[156][2] * mat_B[147][1] +
                mat_A[156][3] * mat_B[155][1] +
                mat_A[157][0] * mat_B[163][1] +
                mat_A[157][1] * mat_B[171][1] +
                mat_A[157][2] * mat_B[179][1] +
                mat_A[157][3] * mat_B[187][1] +
                mat_A[158][0] * mat_B[195][1] +
                mat_A[158][1] * mat_B[203][1] +
                mat_A[158][2] * mat_B[211][1] +
                mat_A[158][3] * mat_B[219][1] +
                mat_A[159][0] * mat_B[227][1] +
                mat_A[159][1] * mat_B[235][1] +
                mat_A[159][2] * mat_B[243][1] +
                mat_A[159][3] * mat_B[251][1];
    mat_C[155][2] <=
                mat_A[152][0] * mat_B[3][2] +
                mat_A[152][1] * mat_B[11][2] +
                mat_A[152][2] * mat_B[19][2] +
                mat_A[152][3] * mat_B[27][2] +
                mat_A[153][0] * mat_B[35][2] +
                mat_A[153][1] * mat_B[43][2] +
                mat_A[153][2] * mat_B[51][2] +
                mat_A[153][3] * mat_B[59][2] +
                mat_A[154][0] * mat_B[67][2] +
                mat_A[154][1] * mat_B[75][2] +
                mat_A[154][2] * mat_B[83][2] +
                mat_A[154][3] * mat_B[91][2] +
                mat_A[155][0] * mat_B[99][2] +
                mat_A[155][1] * mat_B[107][2] +
                mat_A[155][2] * mat_B[115][2] +
                mat_A[155][3] * mat_B[123][2] +
                mat_A[156][0] * mat_B[131][2] +
                mat_A[156][1] * mat_B[139][2] +
                mat_A[156][2] * mat_B[147][2] +
                mat_A[156][3] * mat_B[155][2] +
                mat_A[157][0] * mat_B[163][2] +
                mat_A[157][1] * mat_B[171][2] +
                mat_A[157][2] * mat_B[179][2] +
                mat_A[157][3] * mat_B[187][2] +
                mat_A[158][0] * mat_B[195][2] +
                mat_A[158][1] * mat_B[203][2] +
                mat_A[158][2] * mat_B[211][2] +
                mat_A[158][3] * mat_B[219][2] +
                mat_A[159][0] * mat_B[227][2] +
                mat_A[159][1] * mat_B[235][2] +
                mat_A[159][2] * mat_B[243][2] +
                mat_A[159][3] * mat_B[251][2];
    mat_C[155][3] <=
                mat_A[152][0] * mat_B[3][3] +
                mat_A[152][1] * mat_B[11][3] +
                mat_A[152][2] * mat_B[19][3] +
                mat_A[152][3] * mat_B[27][3] +
                mat_A[153][0] * mat_B[35][3] +
                mat_A[153][1] * mat_B[43][3] +
                mat_A[153][2] * mat_B[51][3] +
                mat_A[153][3] * mat_B[59][3] +
                mat_A[154][0] * mat_B[67][3] +
                mat_A[154][1] * mat_B[75][3] +
                mat_A[154][2] * mat_B[83][3] +
                mat_A[154][3] * mat_B[91][3] +
                mat_A[155][0] * mat_B[99][3] +
                mat_A[155][1] * mat_B[107][3] +
                mat_A[155][2] * mat_B[115][3] +
                mat_A[155][3] * mat_B[123][3] +
                mat_A[156][0] * mat_B[131][3] +
                mat_A[156][1] * mat_B[139][3] +
                mat_A[156][2] * mat_B[147][3] +
                mat_A[156][3] * mat_B[155][3] +
                mat_A[157][0] * mat_B[163][3] +
                mat_A[157][1] * mat_B[171][3] +
                mat_A[157][2] * mat_B[179][3] +
                mat_A[157][3] * mat_B[187][3] +
                mat_A[158][0] * mat_B[195][3] +
                mat_A[158][1] * mat_B[203][3] +
                mat_A[158][2] * mat_B[211][3] +
                mat_A[158][3] * mat_B[219][3] +
                mat_A[159][0] * mat_B[227][3] +
                mat_A[159][1] * mat_B[235][3] +
                mat_A[159][2] * mat_B[243][3] +
                mat_A[159][3] * mat_B[251][3];
    mat_C[156][0] <=
                mat_A[152][0] * mat_B[4][0] +
                mat_A[152][1] * mat_B[12][0] +
                mat_A[152][2] * mat_B[20][0] +
                mat_A[152][3] * mat_B[28][0] +
                mat_A[153][0] * mat_B[36][0] +
                mat_A[153][1] * mat_B[44][0] +
                mat_A[153][2] * mat_B[52][0] +
                mat_A[153][3] * mat_B[60][0] +
                mat_A[154][0] * mat_B[68][0] +
                mat_A[154][1] * mat_B[76][0] +
                mat_A[154][2] * mat_B[84][0] +
                mat_A[154][3] * mat_B[92][0] +
                mat_A[155][0] * mat_B[100][0] +
                mat_A[155][1] * mat_B[108][0] +
                mat_A[155][2] * mat_B[116][0] +
                mat_A[155][3] * mat_B[124][0] +
                mat_A[156][0] * mat_B[132][0] +
                mat_A[156][1] * mat_B[140][0] +
                mat_A[156][2] * mat_B[148][0] +
                mat_A[156][3] * mat_B[156][0] +
                mat_A[157][0] * mat_B[164][0] +
                mat_A[157][1] * mat_B[172][0] +
                mat_A[157][2] * mat_B[180][0] +
                mat_A[157][3] * mat_B[188][0] +
                mat_A[158][0] * mat_B[196][0] +
                mat_A[158][1] * mat_B[204][0] +
                mat_A[158][2] * mat_B[212][0] +
                mat_A[158][3] * mat_B[220][0] +
                mat_A[159][0] * mat_B[228][0] +
                mat_A[159][1] * mat_B[236][0] +
                mat_A[159][2] * mat_B[244][0] +
                mat_A[159][3] * mat_B[252][0];
    mat_C[156][1] <=
                mat_A[152][0] * mat_B[4][1] +
                mat_A[152][1] * mat_B[12][1] +
                mat_A[152][2] * mat_B[20][1] +
                mat_A[152][3] * mat_B[28][1] +
                mat_A[153][0] * mat_B[36][1] +
                mat_A[153][1] * mat_B[44][1] +
                mat_A[153][2] * mat_B[52][1] +
                mat_A[153][3] * mat_B[60][1] +
                mat_A[154][0] * mat_B[68][1] +
                mat_A[154][1] * mat_B[76][1] +
                mat_A[154][2] * mat_B[84][1] +
                mat_A[154][3] * mat_B[92][1] +
                mat_A[155][0] * mat_B[100][1] +
                mat_A[155][1] * mat_B[108][1] +
                mat_A[155][2] * mat_B[116][1] +
                mat_A[155][3] * mat_B[124][1] +
                mat_A[156][0] * mat_B[132][1] +
                mat_A[156][1] * mat_B[140][1] +
                mat_A[156][2] * mat_B[148][1] +
                mat_A[156][3] * mat_B[156][1] +
                mat_A[157][0] * mat_B[164][1] +
                mat_A[157][1] * mat_B[172][1] +
                mat_A[157][2] * mat_B[180][1] +
                mat_A[157][3] * mat_B[188][1] +
                mat_A[158][0] * mat_B[196][1] +
                mat_A[158][1] * mat_B[204][1] +
                mat_A[158][2] * mat_B[212][1] +
                mat_A[158][3] * mat_B[220][1] +
                mat_A[159][0] * mat_B[228][1] +
                mat_A[159][1] * mat_B[236][1] +
                mat_A[159][2] * mat_B[244][1] +
                mat_A[159][3] * mat_B[252][1];
    mat_C[156][2] <=
                mat_A[152][0] * mat_B[4][2] +
                mat_A[152][1] * mat_B[12][2] +
                mat_A[152][2] * mat_B[20][2] +
                mat_A[152][3] * mat_B[28][2] +
                mat_A[153][0] * mat_B[36][2] +
                mat_A[153][1] * mat_B[44][2] +
                mat_A[153][2] * mat_B[52][2] +
                mat_A[153][3] * mat_B[60][2] +
                mat_A[154][0] * mat_B[68][2] +
                mat_A[154][1] * mat_B[76][2] +
                mat_A[154][2] * mat_B[84][2] +
                mat_A[154][3] * mat_B[92][2] +
                mat_A[155][0] * mat_B[100][2] +
                mat_A[155][1] * mat_B[108][2] +
                mat_A[155][2] * mat_B[116][2] +
                mat_A[155][3] * mat_B[124][2] +
                mat_A[156][0] * mat_B[132][2] +
                mat_A[156][1] * mat_B[140][2] +
                mat_A[156][2] * mat_B[148][2] +
                mat_A[156][3] * mat_B[156][2] +
                mat_A[157][0] * mat_B[164][2] +
                mat_A[157][1] * mat_B[172][2] +
                mat_A[157][2] * mat_B[180][2] +
                mat_A[157][3] * mat_B[188][2] +
                mat_A[158][0] * mat_B[196][2] +
                mat_A[158][1] * mat_B[204][2] +
                mat_A[158][2] * mat_B[212][2] +
                mat_A[158][3] * mat_B[220][2] +
                mat_A[159][0] * mat_B[228][2] +
                mat_A[159][1] * mat_B[236][2] +
                mat_A[159][2] * mat_B[244][2] +
                mat_A[159][3] * mat_B[252][2];
    mat_C[156][3] <=
                mat_A[152][0] * mat_B[4][3] +
                mat_A[152][1] * mat_B[12][3] +
                mat_A[152][2] * mat_B[20][3] +
                mat_A[152][3] * mat_B[28][3] +
                mat_A[153][0] * mat_B[36][3] +
                mat_A[153][1] * mat_B[44][3] +
                mat_A[153][2] * mat_B[52][3] +
                mat_A[153][3] * mat_B[60][3] +
                mat_A[154][0] * mat_B[68][3] +
                mat_A[154][1] * mat_B[76][3] +
                mat_A[154][2] * mat_B[84][3] +
                mat_A[154][3] * mat_B[92][3] +
                mat_A[155][0] * mat_B[100][3] +
                mat_A[155][1] * mat_B[108][3] +
                mat_A[155][2] * mat_B[116][3] +
                mat_A[155][3] * mat_B[124][3] +
                mat_A[156][0] * mat_B[132][3] +
                mat_A[156][1] * mat_B[140][3] +
                mat_A[156][2] * mat_B[148][3] +
                mat_A[156][3] * mat_B[156][3] +
                mat_A[157][0] * mat_B[164][3] +
                mat_A[157][1] * mat_B[172][3] +
                mat_A[157][2] * mat_B[180][3] +
                mat_A[157][3] * mat_B[188][3] +
                mat_A[158][0] * mat_B[196][3] +
                mat_A[158][1] * mat_B[204][3] +
                mat_A[158][2] * mat_B[212][3] +
                mat_A[158][3] * mat_B[220][3] +
                mat_A[159][0] * mat_B[228][3] +
                mat_A[159][1] * mat_B[236][3] +
                mat_A[159][2] * mat_B[244][3] +
                mat_A[159][3] * mat_B[252][3];
    mat_C[157][0] <=
                mat_A[152][0] * mat_B[5][0] +
                mat_A[152][1] * mat_B[13][0] +
                mat_A[152][2] * mat_B[21][0] +
                mat_A[152][3] * mat_B[29][0] +
                mat_A[153][0] * mat_B[37][0] +
                mat_A[153][1] * mat_B[45][0] +
                mat_A[153][2] * mat_B[53][0] +
                mat_A[153][3] * mat_B[61][0] +
                mat_A[154][0] * mat_B[69][0] +
                mat_A[154][1] * mat_B[77][0] +
                mat_A[154][2] * mat_B[85][0] +
                mat_A[154][3] * mat_B[93][0] +
                mat_A[155][0] * mat_B[101][0] +
                mat_A[155][1] * mat_B[109][0] +
                mat_A[155][2] * mat_B[117][0] +
                mat_A[155][3] * mat_B[125][0] +
                mat_A[156][0] * mat_B[133][0] +
                mat_A[156][1] * mat_B[141][0] +
                mat_A[156][2] * mat_B[149][0] +
                mat_A[156][3] * mat_B[157][0] +
                mat_A[157][0] * mat_B[165][0] +
                mat_A[157][1] * mat_B[173][0] +
                mat_A[157][2] * mat_B[181][0] +
                mat_A[157][3] * mat_B[189][0] +
                mat_A[158][0] * mat_B[197][0] +
                mat_A[158][1] * mat_B[205][0] +
                mat_A[158][2] * mat_B[213][0] +
                mat_A[158][3] * mat_B[221][0] +
                mat_A[159][0] * mat_B[229][0] +
                mat_A[159][1] * mat_B[237][0] +
                mat_A[159][2] * mat_B[245][0] +
                mat_A[159][3] * mat_B[253][0];
    mat_C[157][1] <=
                mat_A[152][0] * mat_B[5][1] +
                mat_A[152][1] * mat_B[13][1] +
                mat_A[152][2] * mat_B[21][1] +
                mat_A[152][3] * mat_B[29][1] +
                mat_A[153][0] * mat_B[37][1] +
                mat_A[153][1] * mat_B[45][1] +
                mat_A[153][2] * mat_B[53][1] +
                mat_A[153][3] * mat_B[61][1] +
                mat_A[154][0] * mat_B[69][1] +
                mat_A[154][1] * mat_B[77][1] +
                mat_A[154][2] * mat_B[85][1] +
                mat_A[154][3] * mat_B[93][1] +
                mat_A[155][0] * mat_B[101][1] +
                mat_A[155][1] * mat_B[109][1] +
                mat_A[155][2] * mat_B[117][1] +
                mat_A[155][3] * mat_B[125][1] +
                mat_A[156][0] * mat_B[133][1] +
                mat_A[156][1] * mat_B[141][1] +
                mat_A[156][2] * mat_B[149][1] +
                mat_A[156][3] * mat_B[157][1] +
                mat_A[157][0] * mat_B[165][1] +
                mat_A[157][1] * mat_B[173][1] +
                mat_A[157][2] * mat_B[181][1] +
                mat_A[157][3] * mat_B[189][1] +
                mat_A[158][0] * mat_B[197][1] +
                mat_A[158][1] * mat_B[205][1] +
                mat_A[158][2] * mat_B[213][1] +
                mat_A[158][3] * mat_B[221][1] +
                mat_A[159][0] * mat_B[229][1] +
                mat_A[159][1] * mat_B[237][1] +
                mat_A[159][2] * mat_B[245][1] +
                mat_A[159][3] * mat_B[253][1];
    mat_C[157][2] <=
                mat_A[152][0] * mat_B[5][2] +
                mat_A[152][1] * mat_B[13][2] +
                mat_A[152][2] * mat_B[21][2] +
                mat_A[152][3] * mat_B[29][2] +
                mat_A[153][0] * mat_B[37][2] +
                mat_A[153][1] * mat_B[45][2] +
                mat_A[153][2] * mat_B[53][2] +
                mat_A[153][3] * mat_B[61][2] +
                mat_A[154][0] * mat_B[69][2] +
                mat_A[154][1] * mat_B[77][2] +
                mat_A[154][2] * mat_B[85][2] +
                mat_A[154][3] * mat_B[93][2] +
                mat_A[155][0] * mat_B[101][2] +
                mat_A[155][1] * mat_B[109][2] +
                mat_A[155][2] * mat_B[117][2] +
                mat_A[155][3] * mat_B[125][2] +
                mat_A[156][0] * mat_B[133][2] +
                mat_A[156][1] * mat_B[141][2] +
                mat_A[156][2] * mat_B[149][2] +
                mat_A[156][3] * mat_B[157][2] +
                mat_A[157][0] * mat_B[165][2] +
                mat_A[157][1] * mat_B[173][2] +
                mat_A[157][2] * mat_B[181][2] +
                mat_A[157][3] * mat_B[189][2] +
                mat_A[158][0] * mat_B[197][2] +
                mat_A[158][1] * mat_B[205][2] +
                mat_A[158][2] * mat_B[213][2] +
                mat_A[158][3] * mat_B[221][2] +
                mat_A[159][0] * mat_B[229][2] +
                mat_A[159][1] * mat_B[237][2] +
                mat_A[159][2] * mat_B[245][2] +
                mat_A[159][3] * mat_B[253][2];
    mat_C[157][3] <=
                mat_A[152][0] * mat_B[5][3] +
                mat_A[152][1] * mat_B[13][3] +
                mat_A[152][2] * mat_B[21][3] +
                mat_A[152][3] * mat_B[29][3] +
                mat_A[153][0] * mat_B[37][3] +
                mat_A[153][1] * mat_B[45][3] +
                mat_A[153][2] * mat_B[53][3] +
                mat_A[153][3] * mat_B[61][3] +
                mat_A[154][0] * mat_B[69][3] +
                mat_A[154][1] * mat_B[77][3] +
                mat_A[154][2] * mat_B[85][3] +
                mat_A[154][3] * mat_B[93][3] +
                mat_A[155][0] * mat_B[101][3] +
                mat_A[155][1] * mat_B[109][3] +
                mat_A[155][2] * mat_B[117][3] +
                mat_A[155][3] * mat_B[125][3] +
                mat_A[156][0] * mat_B[133][3] +
                mat_A[156][1] * mat_B[141][3] +
                mat_A[156][2] * mat_B[149][3] +
                mat_A[156][3] * mat_B[157][3] +
                mat_A[157][0] * mat_B[165][3] +
                mat_A[157][1] * mat_B[173][3] +
                mat_A[157][2] * mat_B[181][3] +
                mat_A[157][3] * mat_B[189][3] +
                mat_A[158][0] * mat_B[197][3] +
                mat_A[158][1] * mat_B[205][3] +
                mat_A[158][2] * mat_B[213][3] +
                mat_A[158][3] * mat_B[221][3] +
                mat_A[159][0] * mat_B[229][3] +
                mat_A[159][1] * mat_B[237][3] +
                mat_A[159][2] * mat_B[245][3] +
                mat_A[159][3] * mat_B[253][3];
    mat_C[158][0] <=
                mat_A[152][0] * mat_B[6][0] +
                mat_A[152][1] * mat_B[14][0] +
                mat_A[152][2] * mat_B[22][0] +
                mat_A[152][3] * mat_B[30][0] +
                mat_A[153][0] * mat_B[38][0] +
                mat_A[153][1] * mat_B[46][0] +
                mat_A[153][2] * mat_B[54][0] +
                mat_A[153][3] * mat_B[62][0] +
                mat_A[154][0] * mat_B[70][0] +
                mat_A[154][1] * mat_B[78][0] +
                mat_A[154][2] * mat_B[86][0] +
                mat_A[154][3] * mat_B[94][0] +
                mat_A[155][0] * mat_B[102][0] +
                mat_A[155][1] * mat_B[110][0] +
                mat_A[155][2] * mat_B[118][0] +
                mat_A[155][3] * mat_B[126][0] +
                mat_A[156][0] * mat_B[134][0] +
                mat_A[156][1] * mat_B[142][0] +
                mat_A[156][2] * mat_B[150][0] +
                mat_A[156][3] * mat_B[158][0] +
                mat_A[157][0] * mat_B[166][0] +
                mat_A[157][1] * mat_B[174][0] +
                mat_A[157][2] * mat_B[182][0] +
                mat_A[157][3] * mat_B[190][0] +
                mat_A[158][0] * mat_B[198][0] +
                mat_A[158][1] * mat_B[206][0] +
                mat_A[158][2] * mat_B[214][0] +
                mat_A[158][3] * mat_B[222][0] +
                mat_A[159][0] * mat_B[230][0] +
                mat_A[159][1] * mat_B[238][0] +
                mat_A[159][2] * mat_B[246][0] +
                mat_A[159][3] * mat_B[254][0];
    mat_C[158][1] <=
                mat_A[152][0] * mat_B[6][1] +
                mat_A[152][1] * mat_B[14][1] +
                mat_A[152][2] * mat_B[22][1] +
                mat_A[152][3] * mat_B[30][1] +
                mat_A[153][0] * mat_B[38][1] +
                mat_A[153][1] * mat_B[46][1] +
                mat_A[153][2] * mat_B[54][1] +
                mat_A[153][3] * mat_B[62][1] +
                mat_A[154][0] * mat_B[70][1] +
                mat_A[154][1] * mat_B[78][1] +
                mat_A[154][2] * mat_B[86][1] +
                mat_A[154][3] * mat_B[94][1] +
                mat_A[155][0] * mat_B[102][1] +
                mat_A[155][1] * mat_B[110][1] +
                mat_A[155][2] * mat_B[118][1] +
                mat_A[155][3] * mat_B[126][1] +
                mat_A[156][0] * mat_B[134][1] +
                mat_A[156][1] * mat_B[142][1] +
                mat_A[156][2] * mat_B[150][1] +
                mat_A[156][3] * mat_B[158][1] +
                mat_A[157][0] * mat_B[166][1] +
                mat_A[157][1] * mat_B[174][1] +
                mat_A[157][2] * mat_B[182][1] +
                mat_A[157][3] * mat_B[190][1] +
                mat_A[158][0] * mat_B[198][1] +
                mat_A[158][1] * mat_B[206][1] +
                mat_A[158][2] * mat_B[214][1] +
                mat_A[158][3] * mat_B[222][1] +
                mat_A[159][0] * mat_B[230][1] +
                mat_A[159][1] * mat_B[238][1] +
                mat_A[159][2] * mat_B[246][1] +
                mat_A[159][3] * mat_B[254][1];
    mat_C[158][2] <=
                mat_A[152][0] * mat_B[6][2] +
                mat_A[152][1] * mat_B[14][2] +
                mat_A[152][2] * mat_B[22][2] +
                mat_A[152][3] * mat_B[30][2] +
                mat_A[153][0] * mat_B[38][2] +
                mat_A[153][1] * mat_B[46][2] +
                mat_A[153][2] * mat_B[54][2] +
                mat_A[153][3] * mat_B[62][2] +
                mat_A[154][0] * mat_B[70][2] +
                mat_A[154][1] * mat_B[78][2] +
                mat_A[154][2] * mat_B[86][2] +
                mat_A[154][3] * mat_B[94][2] +
                mat_A[155][0] * mat_B[102][2] +
                mat_A[155][1] * mat_B[110][2] +
                mat_A[155][2] * mat_B[118][2] +
                mat_A[155][3] * mat_B[126][2] +
                mat_A[156][0] * mat_B[134][2] +
                mat_A[156][1] * mat_B[142][2] +
                mat_A[156][2] * mat_B[150][2] +
                mat_A[156][3] * mat_B[158][2] +
                mat_A[157][0] * mat_B[166][2] +
                mat_A[157][1] * mat_B[174][2] +
                mat_A[157][2] * mat_B[182][2] +
                mat_A[157][3] * mat_B[190][2] +
                mat_A[158][0] * mat_B[198][2] +
                mat_A[158][1] * mat_B[206][2] +
                mat_A[158][2] * mat_B[214][2] +
                mat_A[158][3] * mat_B[222][2] +
                mat_A[159][0] * mat_B[230][2] +
                mat_A[159][1] * mat_B[238][2] +
                mat_A[159][2] * mat_B[246][2] +
                mat_A[159][3] * mat_B[254][2];
    mat_C[158][3] <=
                mat_A[152][0] * mat_B[6][3] +
                mat_A[152][1] * mat_B[14][3] +
                mat_A[152][2] * mat_B[22][3] +
                mat_A[152][3] * mat_B[30][3] +
                mat_A[153][0] * mat_B[38][3] +
                mat_A[153][1] * mat_B[46][3] +
                mat_A[153][2] * mat_B[54][3] +
                mat_A[153][3] * mat_B[62][3] +
                mat_A[154][0] * mat_B[70][3] +
                mat_A[154][1] * mat_B[78][3] +
                mat_A[154][2] * mat_B[86][3] +
                mat_A[154][3] * mat_B[94][3] +
                mat_A[155][0] * mat_B[102][3] +
                mat_A[155][1] * mat_B[110][3] +
                mat_A[155][2] * mat_B[118][3] +
                mat_A[155][3] * mat_B[126][3] +
                mat_A[156][0] * mat_B[134][3] +
                mat_A[156][1] * mat_B[142][3] +
                mat_A[156][2] * mat_B[150][3] +
                mat_A[156][3] * mat_B[158][3] +
                mat_A[157][0] * mat_B[166][3] +
                mat_A[157][1] * mat_B[174][3] +
                mat_A[157][2] * mat_B[182][3] +
                mat_A[157][3] * mat_B[190][3] +
                mat_A[158][0] * mat_B[198][3] +
                mat_A[158][1] * mat_B[206][3] +
                mat_A[158][2] * mat_B[214][3] +
                mat_A[158][3] * mat_B[222][3] +
                mat_A[159][0] * mat_B[230][3] +
                mat_A[159][1] * mat_B[238][3] +
                mat_A[159][2] * mat_B[246][3] +
                mat_A[159][3] * mat_B[254][3];
    mat_C[159][0] <=
                mat_A[152][0] * mat_B[7][0] +
                mat_A[152][1] * mat_B[15][0] +
                mat_A[152][2] * mat_B[23][0] +
                mat_A[152][3] * mat_B[31][0] +
                mat_A[153][0] * mat_B[39][0] +
                mat_A[153][1] * mat_B[47][0] +
                mat_A[153][2] * mat_B[55][0] +
                mat_A[153][3] * mat_B[63][0] +
                mat_A[154][0] * mat_B[71][0] +
                mat_A[154][1] * mat_B[79][0] +
                mat_A[154][2] * mat_B[87][0] +
                mat_A[154][3] * mat_B[95][0] +
                mat_A[155][0] * mat_B[103][0] +
                mat_A[155][1] * mat_B[111][0] +
                mat_A[155][2] * mat_B[119][0] +
                mat_A[155][3] * mat_B[127][0] +
                mat_A[156][0] * mat_B[135][0] +
                mat_A[156][1] * mat_B[143][0] +
                mat_A[156][2] * mat_B[151][0] +
                mat_A[156][3] * mat_B[159][0] +
                mat_A[157][0] * mat_B[167][0] +
                mat_A[157][1] * mat_B[175][0] +
                mat_A[157][2] * mat_B[183][0] +
                mat_A[157][3] * mat_B[191][0] +
                mat_A[158][0] * mat_B[199][0] +
                mat_A[158][1] * mat_B[207][0] +
                mat_A[158][2] * mat_B[215][0] +
                mat_A[158][3] * mat_B[223][0] +
                mat_A[159][0] * mat_B[231][0] +
                mat_A[159][1] * mat_B[239][0] +
                mat_A[159][2] * mat_B[247][0] +
                mat_A[159][3] * mat_B[255][0];
    mat_C[159][1] <=
                mat_A[152][0] * mat_B[7][1] +
                mat_A[152][1] * mat_B[15][1] +
                mat_A[152][2] * mat_B[23][1] +
                mat_A[152][3] * mat_B[31][1] +
                mat_A[153][0] * mat_B[39][1] +
                mat_A[153][1] * mat_B[47][1] +
                mat_A[153][2] * mat_B[55][1] +
                mat_A[153][3] * mat_B[63][1] +
                mat_A[154][0] * mat_B[71][1] +
                mat_A[154][1] * mat_B[79][1] +
                mat_A[154][2] * mat_B[87][1] +
                mat_A[154][3] * mat_B[95][1] +
                mat_A[155][0] * mat_B[103][1] +
                mat_A[155][1] * mat_B[111][1] +
                mat_A[155][2] * mat_B[119][1] +
                mat_A[155][3] * mat_B[127][1] +
                mat_A[156][0] * mat_B[135][1] +
                mat_A[156][1] * mat_B[143][1] +
                mat_A[156][2] * mat_B[151][1] +
                mat_A[156][3] * mat_B[159][1] +
                mat_A[157][0] * mat_B[167][1] +
                mat_A[157][1] * mat_B[175][1] +
                mat_A[157][2] * mat_B[183][1] +
                mat_A[157][3] * mat_B[191][1] +
                mat_A[158][0] * mat_B[199][1] +
                mat_A[158][1] * mat_B[207][1] +
                mat_A[158][2] * mat_B[215][1] +
                mat_A[158][3] * mat_B[223][1] +
                mat_A[159][0] * mat_B[231][1] +
                mat_A[159][1] * mat_B[239][1] +
                mat_A[159][2] * mat_B[247][1] +
                mat_A[159][3] * mat_B[255][1];
    mat_C[159][2] <=
                mat_A[152][0] * mat_B[7][2] +
                mat_A[152][1] * mat_B[15][2] +
                mat_A[152][2] * mat_B[23][2] +
                mat_A[152][3] * mat_B[31][2] +
                mat_A[153][0] * mat_B[39][2] +
                mat_A[153][1] * mat_B[47][2] +
                mat_A[153][2] * mat_B[55][2] +
                mat_A[153][3] * mat_B[63][2] +
                mat_A[154][0] * mat_B[71][2] +
                mat_A[154][1] * mat_B[79][2] +
                mat_A[154][2] * mat_B[87][2] +
                mat_A[154][3] * mat_B[95][2] +
                mat_A[155][0] * mat_B[103][2] +
                mat_A[155][1] * mat_B[111][2] +
                mat_A[155][2] * mat_B[119][2] +
                mat_A[155][3] * mat_B[127][2] +
                mat_A[156][0] * mat_B[135][2] +
                mat_A[156][1] * mat_B[143][2] +
                mat_A[156][2] * mat_B[151][2] +
                mat_A[156][3] * mat_B[159][2] +
                mat_A[157][0] * mat_B[167][2] +
                mat_A[157][1] * mat_B[175][2] +
                mat_A[157][2] * mat_B[183][2] +
                mat_A[157][3] * mat_B[191][2] +
                mat_A[158][0] * mat_B[199][2] +
                mat_A[158][1] * mat_B[207][2] +
                mat_A[158][2] * mat_B[215][2] +
                mat_A[158][3] * mat_B[223][2] +
                mat_A[159][0] * mat_B[231][2] +
                mat_A[159][1] * mat_B[239][2] +
                mat_A[159][2] * mat_B[247][2] +
                mat_A[159][3] * mat_B[255][2];
    mat_C[159][3] <=
                mat_A[152][0] * mat_B[7][3] +
                mat_A[152][1] * mat_B[15][3] +
                mat_A[152][2] * mat_B[23][3] +
                mat_A[152][3] * mat_B[31][3] +
                mat_A[153][0] * mat_B[39][3] +
                mat_A[153][1] * mat_B[47][3] +
                mat_A[153][2] * mat_B[55][3] +
                mat_A[153][3] * mat_B[63][3] +
                mat_A[154][0] * mat_B[71][3] +
                mat_A[154][1] * mat_B[79][3] +
                mat_A[154][2] * mat_B[87][3] +
                mat_A[154][3] * mat_B[95][3] +
                mat_A[155][0] * mat_B[103][3] +
                mat_A[155][1] * mat_B[111][3] +
                mat_A[155][2] * mat_B[119][3] +
                mat_A[155][3] * mat_B[127][3] +
                mat_A[156][0] * mat_B[135][3] +
                mat_A[156][1] * mat_B[143][3] +
                mat_A[156][2] * mat_B[151][3] +
                mat_A[156][3] * mat_B[159][3] +
                mat_A[157][0] * mat_B[167][3] +
                mat_A[157][1] * mat_B[175][3] +
                mat_A[157][2] * mat_B[183][3] +
                mat_A[157][3] * mat_B[191][3] +
                mat_A[158][0] * mat_B[199][3] +
                mat_A[158][1] * mat_B[207][3] +
                mat_A[158][2] * mat_B[215][3] +
                mat_A[158][3] * mat_B[223][3] +
                mat_A[159][0] * mat_B[231][3] +
                mat_A[159][1] * mat_B[239][3] +
                mat_A[159][2] * mat_B[247][3] +
                mat_A[159][3] * mat_B[255][3];
    mat_C[160][0] <=
                mat_A[160][0] * mat_B[0][0] +
                mat_A[160][1] * mat_B[8][0] +
                mat_A[160][2] * mat_B[16][0] +
                mat_A[160][3] * mat_B[24][0] +
                mat_A[161][0] * mat_B[32][0] +
                mat_A[161][1] * mat_B[40][0] +
                mat_A[161][2] * mat_B[48][0] +
                mat_A[161][3] * mat_B[56][0] +
                mat_A[162][0] * mat_B[64][0] +
                mat_A[162][1] * mat_B[72][0] +
                mat_A[162][2] * mat_B[80][0] +
                mat_A[162][3] * mat_B[88][0] +
                mat_A[163][0] * mat_B[96][0] +
                mat_A[163][1] * mat_B[104][0] +
                mat_A[163][2] * mat_B[112][0] +
                mat_A[163][3] * mat_B[120][0] +
                mat_A[164][0] * mat_B[128][0] +
                mat_A[164][1] * mat_B[136][0] +
                mat_A[164][2] * mat_B[144][0] +
                mat_A[164][3] * mat_B[152][0] +
                mat_A[165][0] * mat_B[160][0] +
                mat_A[165][1] * mat_B[168][0] +
                mat_A[165][2] * mat_B[176][0] +
                mat_A[165][3] * mat_B[184][0] +
                mat_A[166][0] * mat_B[192][0] +
                mat_A[166][1] * mat_B[200][0] +
                mat_A[166][2] * mat_B[208][0] +
                mat_A[166][3] * mat_B[216][0] +
                mat_A[167][0] * mat_B[224][0] +
                mat_A[167][1] * mat_B[232][0] +
                mat_A[167][2] * mat_B[240][0] +
                mat_A[167][3] * mat_B[248][0];
    mat_C[160][1] <=
                mat_A[160][0] * mat_B[0][1] +
                mat_A[160][1] * mat_B[8][1] +
                mat_A[160][2] * mat_B[16][1] +
                mat_A[160][3] * mat_B[24][1] +
                mat_A[161][0] * mat_B[32][1] +
                mat_A[161][1] * mat_B[40][1] +
                mat_A[161][2] * mat_B[48][1] +
                mat_A[161][3] * mat_B[56][1] +
                mat_A[162][0] * mat_B[64][1] +
                mat_A[162][1] * mat_B[72][1] +
                mat_A[162][2] * mat_B[80][1] +
                mat_A[162][3] * mat_B[88][1] +
                mat_A[163][0] * mat_B[96][1] +
                mat_A[163][1] * mat_B[104][1] +
                mat_A[163][2] * mat_B[112][1] +
                mat_A[163][3] * mat_B[120][1] +
                mat_A[164][0] * mat_B[128][1] +
                mat_A[164][1] * mat_B[136][1] +
                mat_A[164][2] * mat_B[144][1] +
                mat_A[164][3] * mat_B[152][1] +
                mat_A[165][0] * mat_B[160][1] +
                mat_A[165][1] * mat_B[168][1] +
                mat_A[165][2] * mat_B[176][1] +
                mat_A[165][3] * mat_B[184][1] +
                mat_A[166][0] * mat_B[192][1] +
                mat_A[166][1] * mat_B[200][1] +
                mat_A[166][2] * mat_B[208][1] +
                mat_A[166][3] * mat_B[216][1] +
                mat_A[167][0] * mat_B[224][1] +
                mat_A[167][1] * mat_B[232][1] +
                mat_A[167][2] * mat_B[240][1] +
                mat_A[167][3] * mat_B[248][1];
    mat_C[160][2] <=
                mat_A[160][0] * mat_B[0][2] +
                mat_A[160][1] * mat_B[8][2] +
                mat_A[160][2] * mat_B[16][2] +
                mat_A[160][3] * mat_B[24][2] +
                mat_A[161][0] * mat_B[32][2] +
                mat_A[161][1] * mat_B[40][2] +
                mat_A[161][2] * mat_B[48][2] +
                mat_A[161][3] * mat_B[56][2] +
                mat_A[162][0] * mat_B[64][2] +
                mat_A[162][1] * mat_B[72][2] +
                mat_A[162][2] * mat_B[80][2] +
                mat_A[162][3] * mat_B[88][2] +
                mat_A[163][0] * mat_B[96][2] +
                mat_A[163][1] * mat_B[104][2] +
                mat_A[163][2] * mat_B[112][2] +
                mat_A[163][3] * mat_B[120][2] +
                mat_A[164][0] * mat_B[128][2] +
                mat_A[164][1] * mat_B[136][2] +
                mat_A[164][2] * mat_B[144][2] +
                mat_A[164][3] * mat_B[152][2] +
                mat_A[165][0] * mat_B[160][2] +
                mat_A[165][1] * mat_B[168][2] +
                mat_A[165][2] * mat_B[176][2] +
                mat_A[165][3] * mat_B[184][2] +
                mat_A[166][0] * mat_B[192][2] +
                mat_A[166][1] * mat_B[200][2] +
                mat_A[166][2] * mat_B[208][2] +
                mat_A[166][3] * mat_B[216][2] +
                mat_A[167][0] * mat_B[224][2] +
                mat_A[167][1] * mat_B[232][2] +
                mat_A[167][2] * mat_B[240][2] +
                mat_A[167][3] * mat_B[248][2];
    mat_C[160][3] <=
                mat_A[160][0] * mat_B[0][3] +
                mat_A[160][1] * mat_B[8][3] +
                mat_A[160][2] * mat_B[16][3] +
                mat_A[160][3] * mat_B[24][3] +
                mat_A[161][0] * mat_B[32][3] +
                mat_A[161][1] * mat_B[40][3] +
                mat_A[161][2] * mat_B[48][3] +
                mat_A[161][3] * mat_B[56][3] +
                mat_A[162][0] * mat_B[64][3] +
                mat_A[162][1] * mat_B[72][3] +
                mat_A[162][2] * mat_B[80][3] +
                mat_A[162][3] * mat_B[88][3] +
                mat_A[163][0] * mat_B[96][3] +
                mat_A[163][1] * mat_B[104][3] +
                mat_A[163][2] * mat_B[112][3] +
                mat_A[163][3] * mat_B[120][3] +
                mat_A[164][0] * mat_B[128][3] +
                mat_A[164][1] * mat_B[136][3] +
                mat_A[164][2] * mat_B[144][3] +
                mat_A[164][3] * mat_B[152][3] +
                mat_A[165][0] * mat_B[160][3] +
                mat_A[165][1] * mat_B[168][3] +
                mat_A[165][2] * mat_B[176][3] +
                mat_A[165][3] * mat_B[184][3] +
                mat_A[166][0] * mat_B[192][3] +
                mat_A[166][1] * mat_B[200][3] +
                mat_A[166][2] * mat_B[208][3] +
                mat_A[166][3] * mat_B[216][3] +
                mat_A[167][0] * mat_B[224][3] +
                mat_A[167][1] * mat_B[232][3] +
                mat_A[167][2] * mat_B[240][3] +
                mat_A[167][3] * mat_B[248][3];
    mat_C[161][0] <=
                mat_A[160][0] * mat_B[1][0] +
                mat_A[160][1] * mat_B[9][0] +
                mat_A[160][2] * mat_B[17][0] +
                mat_A[160][3] * mat_B[25][0] +
                mat_A[161][0] * mat_B[33][0] +
                mat_A[161][1] * mat_B[41][0] +
                mat_A[161][2] * mat_B[49][0] +
                mat_A[161][3] * mat_B[57][0] +
                mat_A[162][0] * mat_B[65][0] +
                mat_A[162][1] * mat_B[73][0] +
                mat_A[162][2] * mat_B[81][0] +
                mat_A[162][3] * mat_B[89][0] +
                mat_A[163][0] * mat_B[97][0] +
                mat_A[163][1] * mat_B[105][0] +
                mat_A[163][2] * mat_B[113][0] +
                mat_A[163][3] * mat_B[121][0] +
                mat_A[164][0] * mat_B[129][0] +
                mat_A[164][1] * mat_B[137][0] +
                mat_A[164][2] * mat_B[145][0] +
                mat_A[164][3] * mat_B[153][0] +
                mat_A[165][0] * mat_B[161][0] +
                mat_A[165][1] * mat_B[169][0] +
                mat_A[165][2] * mat_B[177][0] +
                mat_A[165][3] * mat_B[185][0] +
                mat_A[166][0] * mat_B[193][0] +
                mat_A[166][1] * mat_B[201][0] +
                mat_A[166][2] * mat_B[209][0] +
                mat_A[166][3] * mat_B[217][0] +
                mat_A[167][0] * mat_B[225][0] +
                mat_A[167][1] * mat_B[233][0] +
                mat_A[167][2] * mat_B[241][0] +
                mat_A[167][3] * mat_B[249][0];
    mat_C[161][1] <=
                mat_A[160][0] * mat_B[1][1] +
                mat_A[160][1] * mat_B[9][1] +
                mat_A[160][2] * mat_B[17][1] +
                mat_A[160][3] * mat_B[25][1] +
                mat_A[161][0] * mat_B[33][1] +
                mat_A[161][1] * mat_B[41][1] +
                mat_A[161][2] * mat_B[49][1] +
                mat_A[161][3] * mat_B[57][1] +
                mat_A[162][0] * mat_B[65][1] +
                mat_A[162][1] * mat_B[73][1] +
                mat_A[162][2] * mat_B[81][1] +
                mat_A[162][3] * mat_B[89][1] +
                mat_A[163][0] * mat_B[97][1] +
                mat_A[163][1] * mat_B[105][1] +
                mat_A[163][2] * mat_B[113][1] +
                mat_A[163][3] * mat_B[121][1] +
                mat_A[164][0] * mat_B[129][1] +
                mat_A[164][1] * mat_B[137][1] +
                mat_A[164][2] * mat_B[145][1] +
                mat_A[164][3] * mat_B[153][1] +
                mat_A[165][0] * mat_B[161][1] +
                mat_A[165][1] * mat_B[169][1] +
                mat_A[165][2] * mat_B[177][1] +
                mat_A[165][3] * mat_B[185][1] +
                mat_A[166][0] * mat_B[193][1] +
                mat_A[166][1] * mat_B[201][1] +
                mat_A[166][2] * mat_B[209][1] +
                mat_A[166][3] * mat_B[217][1] +
                mat_A[167][0] * mat_B[225][1] +
                mat_A[167][1] * mat_B[233][1] +
                mat_A[167][2] * mat_B[241][1] +
                mat_A[167][3] * mat_B[249][1];
    mat_C[161][2] <=
                mat_A[160][0] * mat_B[1][2] +
                mat_A[160][1] * mat_B[9][2] +
                mat_A[160][2] * mat_B[17][2] +
                mat_A[160][3] * mat_B[25][2] +
                mat_A[161][0] * mat_B[33][2] +
                mat_A[161][1] * mat_B[41][2] +
                mat_A[161][2] * mat_B[49][2] +
                mat_A[161][3] * mat_B[57][2] +
                mat_A[162][0] * mat_B[65][2] +
                mat_A[162][1] * mat_B[73][2] +
                mat_A[162][2] * mat_B[81][2] +
                mat_A[162][3] * mat_B[89][2] +
                mat_A[163][0] * mat_B[97][2] +
                mat_A[163][1] * mat_B[105][2] +
                mat_A[163][2] * mat_B[113][2] +
                mat_A[163][3] * mat_B[121][2] +
                mat_A[164][0] * mat_B[129][2] +
                mat_A[164][1] * mat_B[137][2] +
                mat_A[164][2] * mat_B[145][2] +
                mat_A[164][3] * mat_B[153][2] +
                mat_A[165][0] * mat_B[161][2] +
                mat_A[165][1] * mat_B[169][2] +
                mat_A[165][2] * mat_B[177][2] +
                mat_A[165][3] * mat_B[185][2] +
                mat_A[166][0] * mat_B[193][2] +
                mat_A[166][1] * mat_B[201][2] +
                mat_A[166][2] * mat_B[209][2] +
                mat_A[166][3] * mat_B[217][2] +
                mat_A[167][0] * mat_B[225][2] +
                mat_A[167][1] * mat_B[233][2] +
                mat_A[167][2] * mat_B[241][2] +
                mat_A[167][3] * mat_B[249][2];
    mat_C[161][3] <=
                mat_A[160][0] * mat_B[1][3] +
                mat_A[160][1] * mat_B[9][3] +
                mat_A[160][2] * mat_B[17][3] +
                mat_A[160][3] * mat_B[25][3] +
                mat_A[161][0] * mat_B[33][3] +
                mat_A[161][1] * mat_B[41][3] +
                mat_A[161][2] * mat_B[49][3] +
                mat_A[161][3] * mat_B[57][3] +
                mat_A[162][0] * mat_B[65][3] +
                mat_A[162][1] * mat_B[73][3] +
                mat_A[162][2] * mat_B[81][3] +
                mat_A[162][3] * mat_B[89][3] +
                mat_A[163][0] * mat_B[97][3] +
                mat_A[163][1] * mat_B[105][3] +
                mat_A[163][2] * mat_B[113][3] +
                mat_A[163][3] * mat_B[121][3] +
                mat_A[164][0] * mat_B[129][3] +
                mat_A[164][1] * mat_B[137][3] +
                mat_A[164][2] * mat_B[145][3] +
                mat_A[164][3] * mat_B[153][3] +
                mat_A[165][0] * mat_B[161][3] +
                mat_A[165][1] * mat_B[169][3] +
                mat_A[165][2] * mat_B[177][3] +
                mat_A[165][3] * mat_B[185][3] +
                mat_A[166][0] * mat_B[193][3] +
                mat_A[166][1] * mat_B[201][3] +
                mat_A[166][2] * mat_B[209][3] +
                mat_A[166][3] * mat_B[217][3] +
                mat_A[167][0] * mat_B[225][3] +
                mat_A[167][1] * mat_B[233][3] +
                mat_A[167][2] * mat_B[241][3] +
                mat_A[167][3] * mat_B[249][3];
    mat_C[162][0] <=
                mat_A[160][0] * mat_B[2][0] +
                mat_A[160][1] * mat_B[10][0] +
                mat_A[160][2] * mat_B[18][0] +
                mat_A[160][3] * mat_B[26][0] +
                mat_A[161][0] * mat_B[34][0] +
                mat_A[161][1] * mat_B[42][0] +
                mat_A[161][2] * mat_B[50][0] +
                mat_A[161][3] * mat_B[58][0] +
                mat_A[162][0] * mat_B[66][0] +
                mat_A[162][1] * mat_B[74][0] +
                mat_A[162][2] * mat_B[82][0] +
                mat_A[162][3] * mat_B[90][0] +
                mat_A[163][0] * mat_B[98][0] +
                mat_A[163][1] * mat_B[106][0] +
                mat_A[163][2] * mat_B[114][0] +
                mat_A[163][3] * mat_B[122][0] +
                mat_A[164][0] * mat_B[130][0] +
                mat_A[164][1] * mat_B[138][0] +
                mat_A[164][2] * mat_B[146][0] +
                mat_A[164][3] * mat_B[154][0] +
                mat_A[165][0] * mat_B[162][0] +
                mat_A[165][1] * mat_B[170][0] +
                mat_A[165][2] * mat_B[178][0] +
                mat_A[165][3] * mat_B[186][0] +
                mat_A[166][0] * mat_B[194][0] +
                mat_A[166][1] * mat_B[202][0] +
                mat_A[166][2] * mat_B[210][0] +
                mat_A[166][3] * mat_B[218][0] +
                mat_A[167][0] * mat_B[226][0] +
                mat_A[167][1] * mat_B[234][0] +
                mat_A[167][2] * mat_B[242][0] +
                mat_A[167][3] * mat_B[250][0];
    mat_C[162][1] <=
                mat_A[160][0] * mat_B[2][1] +
                mat_A[160][1] * mat_B[10][1] +
                mat_A[160][2] * mat_B[18][1] +
                mat_A[160][3] * mat_B[26][1] +
                mat_A[161][0] * mat_B[34][1] +
                mat_A[161][1] * mat_B[42][1] +
                mat_A[161][2] * mat_B[50][1] +
                mat_A[161][3] * mat_B[58][1] +
                mat_A[162][0] * mat_B[66][1] +
                mat_A[162][1] * mat_B[74][1] +
                mat_A[162][2] * mat_B[82][1] +
                mat_A[162][3] * mat_B[90][1] +
                mat_A[163][0] * mat_B[98][1] +
                mat_A[163][1] * mat_B[106][1] +
                mat_A[163][2] * mat_B[114][1] +
                mat_A[163][3] * mat_B[122][1] +
                mat_A[164][0] * mat_B[130][1] +
                mat_A[164][1] * mat_B[138][1] +
                mat_A[164][2] * mat_B[146][1] +
                mat_A[164][3] * mat_B[154][1] +
                mat_A[165][0] * mat_B[162][1] +
                mat_A[165][1] * mat_B[170][1] +
                mat_A[165][2] * mat_B[178][1] +
                mat_A[165][3] * mat_B[186][1] +
                mat_A[166][0] * mat_B[194][1] +
                mat_A[166][1] * mat_B[202][1] +
                mat_A[166][2] * mat_B[210][1] +
                mat_A[166][3] * mat_B[218][1] +
                mat_A[167][0] * mat_B[226][1] +
                mat_A[167][1] * mat_B[234][1] +
                mat_A[167][2] * mat_B[242][1] +
                mat_A[167][3] * mat_B[250][1];
    mat_C[162][2] <=
                mat_A[160][0] * mat_B[2][2] +
                mat_A[160][1] * mat_B[10][2] +
                mat_A[160][2] * mat_B[18][2] +
                mat_A[160][3] * mat_B[26][2] +
                mat_A[161][0] * mat_B[34][2] +
                mat_A[161][1] * mat_B[42][2] +
                mat_A[161][2] * mat_B[50][2] +
                mat_A[161][3] * mat_B[58][2] +
                mat_A[162][0] * mat_B[66][2] +
                mat_A[162][1] * mat_B[74][2] +
                mat_A[162][2] * mat_B[82][2] +
                mat_A[162][3] * mat_B[90][2] +
                mat_A[163][0] * mat_B[98][2] +
                mat_A[163][1] * mat_B[106][2] +
                mat_A[163][2] * mat_B[114][2] +
                mat_A[163][3] * mat_B[122][2] +
                mat_A[164][0] * mat_B[130][2] +
                mat_A[164][1] * mat_B[138][2] +
                mat_A[164][2] * mat_B[146][2] +
                mat_A[164][3] * mat_B[154][2] +
                mat_A[165][0] * mat_B[162][2] +
                mat_A[165][1] * mat_B[170][2] +
                mat_A[165][2] * mat_B[178][2] +
                mat_A[165][3] * mat_B[186][2] +
                mat_A[166][0] * mat_B[194][2] +
                mat_A[166][1] * mat_B[202][2] +
                mat_A[166][2] * mat_B[210][2] +
                mat_A[166][3] * mat_B[218][2] +
                mat_A[167][0] * mat_B[226][2] +
                mat_A[167][1] * mat_B[234][2] +
                mat_A[167][2] * mat_B[242][2] +
                mat_A[167][3] * mat_B[250][2];
    mat_C[162][3] <=
                mat_A[160][0] * mat_B[2][3] +
                mat_A[160][1] * mat_B[10][3] +
                mat_A[160][2] * mat_B[18][3] +
                mat_A[160][3] * mat_B[26][3] +
                mat_A[161][0] * mat_B[34][3] +
                mat_A[161][1] * mat_B[42][3] +
                mat_A[161][2] * mat_B[50][3] +
                mat_A[161][3] * mat_B[58][3] +
                mat_A[162][0] * mat_B[66][3] +
                mat_A[162][1] * mat_B[74][3] +
                mat_A[162][2] * mat_B[82][3] +
                mat_A[162][3] * mat_B[90][3] +
                mat_A[163][0] * mat_B[98][3] +
                mat_A[163][1] * mat_B[106][3] +
                mat_A[163][2] * mat_B[114][3] +
                mat_A[163][3] * mat_B[122][3] +
                mat_A[164][0] * mat_B[130][3] +
                mat_A[164][1] * mat_B[138][3] +
                mat_A[164][2] * mat_B[146][3] +
                mat_A[164][3] * mat_B[154][3] +
                mat_A[165][0] * mat_B[162][3] +
                mat_A[165][1] * mat_B[170][3] +
                mat_A[165][2] * mat_B[178][3] +
                mat_A[165][3] * mat_B[186][3] +
                mat_A[166][0] * mat_B[194][3] +
                mat_A[166][1] * mat_B[202][3] +
                mat_A[166][2] * mat_B[210][3] +
                mat_A[166][3] * mat_B[218][3] +
                mat_A[167][0] * mat_B[226][3] +
                mat_A[167][1] * mat_B[234][3] +
                mat_A[167][2] * mat_B[242][3] +
                mat_A[167][3] * mat_B[250][3];
    mat_C[163][0] <=
                mat_A[160][0] * mat_B[3][0] +
                mat_A[160][1] * mat_B[11][0] +
                mat_A[160][2] * mat_B[19][0] +
                mat_A[160][3] * mat_B[27][0] +
                mat_A[161][0] * mat_B[35][0] +
                mat_A[161][1] * mat_B[43][0] +
                mat_A[161][2] * mat_B[51][0] +
                mat_A[161][3] * mat_B[59][0] +
                mat_A[162][0] * mat_B[67][0] +
                mat_A[162][1] * mat_B[75][0] +
                mat_A[162][2] * mat_B[83][0] +
                mat_A[162][3] * mat_B[91][0] +
                mat_A[163][0] * mat_B[99][0] +
                mat_A[163][1] * mat_B[107][0] +
                mat_A[163][2] * mat_B[115][0] +
                mat_A[163][3] * mat_B[123][0] +
                mat_A[164][0] * mat_B[131][0] +
                mat_A[164][1] * mat_B[139][0] +
                mat_A[164][2] * mat_B[147][0] +
                mat_A[164][3] * mat_B[155][0] +
                mat_A[165][0] * mat_B[163][0] +
                mat_A[165][1] * mat_B[171][0] +
                mat_A[165][2] * mat_B[179][0] +
                mat_A[165][3] * mat_B[187][0] +
                mat_A[166][0] * mat_B[195][0] +
                mat_A[166][1] * mat_B[203][0] +
                mat_A[166][2] * mat_B[211][0] +
                mat_A[166][3] * mat_B[219][0] +
                mat_A[167][0] * mat_B[227][0] +
                mat_A[167][1] * mat_B[235][0] +
                mat_A[167][2] * mat_B[243][0] +
                mat_A[167][3] * mat_B[251][0];
    mat_C[163][1] <=
                mat_A[160][0] * mat_B[3][1] +
                mat_A[160][1] * mat_B[11][1] +
                mat_A[160][2] * mat_B[19][1] +
                mat_A[160][3] * mat_B[27][1] +
                mat_A[161][0] * mat_B[35][1] +
                mat_A[161][1] * mat_B[43][1] +
                mat_A[161][2] * mat_B[51][1] +
                mat_A[161][3] * mat_B[59][1] +
                mat_A[162][0] * mat_B[67][1] +
                mat_A[162][1] * mat_B[75][1] +
                mat_A[162][2] * mat_B[83][1] +
                mat_A[162][3] * mat_B[91][1] +
                mat_A[163][0] * mat_B[99][1] +
                mat_A[163][1] * mat_B[107][1] +
                mat_A[163][2] * mat_B[115][1] +
                mat_A[163][3] * mat_B[123][1] +
                mat_A[164][0] * mat_B[131][1] +
                mat_A[164][1] * mat_B[139][1] +
                mat_A[164][2] * mat_B[147][1] +
                mat_A[164][3] * mat_B[155][1] +
                mat_A[165][0] * mat_B[163][1] +
                mat_A[165][1] * mat_B[171][1] +
                mat_A[165][2] * mat_B[179][1] +
                mat_A[165][3] * mat_B[187][1] +
                mat_A[166][0] * mat_B[195][1] +
                mat_A[166][1] * mat_B[203][1] +
                mat_A[166][2] * mat_B[211][1] +
                mat_A[166][3] * mat_B[219][1] +
                mat_A[167][0] * mat_B[227][1] +
                mat_A[167][1] * mat_B[235][1] +
                mat_A[167][2] * mat_B[243][1] +
                mat_A[167][3] * mat_B[251][1];
    mat_C[163][2] <=
                mat_A[160][0] * mat_B[3][2] +
                mat_A[160][1] * mat_B[11][2] +
                mat_A[160][2] * mat_B[19][2] +
                mat_A[160][3] * mat_B[27][2] +
                mat_A[161][0] * mat_B[35][2] +
                mat_A[161][1] * mat_B[43][2] +
                mat_A[161][2] * mat_B[51][2] +
                mat_A[161][3] * mat_B[59][2] +
                mat_A[162][0] * mat_B[67][2] +
                mat_A[162][1] * mat_B[75][2] +
                mat_A[162][2] * mat_B[83][2] +
                mat_A[162][3] * mat_B[91][2] +
                mat_A[163][0] * mat_B[99][2] +
                mat_A[163][1] * mat_B[107][2] +
                mat_A[163][2] * mat_B[115][2] +
                mat_A[163][3] * mat_B[123][2] +
                mat_A[164][0] * mat_B[131][2] +
                mat_A[164][1] * mat_B[139][2] +
                mat_A[164][2] * mat_B[147][2] +
                mat_A[164][3] * mat_B[155][2] +
                mat_A[165][0] * mat_B[163][2] +
                mat_A[165][1] * mat_B[171][2] +
                mat_A[165][2] * mat_B[179][2] +
                mat_A[165][3] * mat_B[187][2] +
                mat_A[166][0] * mat_B[195][2] +
                mat_A[166][1] * mat_B[203][2] +
                mat_A[166][2] * mat_B[211][2] +
                mat_A[166][3] * mat_B[219][2] +
                mat_A[167][0] * mat_B[227][2] +
                mat_A[167][1] * mat_B[235][2] +
                mat_A[167][2] * mat_B[243][2] +
                mat_A[167][3] * mat_B[251][2];
    mat_C[163][3] <=
                mat_A[160][0] * mat_B[3][3] +
                mat_A[160][1] * mat_B[11][3] +
                mat_A[160][2] * mat_B[19][3] +
                mat_A[160][3] * mat_B[27][3] +
                mat_A[161][0] * mat_B[35][3] +
                mat_A[161][1] * mat_B[43][3] +
                mat_A[161][2] * mat_B[51][3] +
                mat_A[161][3] * mat_B[59][3] +
                mat_A[162][0] * mat_B[67][3] +
                mat_A[162][1] * mat_B[75][3] +
                mat_A[162][2] * mat_B[83][3] +
                mat_A[162][3] * mat_B[91][3] +
                mat_A[163][0] * mat_B[99][3] +
                mat_A[163][1] * mat_B[107][3] +
                mat_A[163][2] * mat_B[115][3] +
                mat_A[163][3] * mat_B[123][3] +
                mat_A[164][0] * mat_B[131][3] +
                mat_A[164][1] * mat_B[139][3] +
                mat_A[164][2] * mat_B[147][3] +
                mat_A[164][3] * mat_B[155][3] +
                mat_A[165][0] * mat_B[163][3] +
                mat_A[165][1] * mat_B[171][3] +
                mat_A[165][2] * mat_B[179][3] +
                mat_A[165][3] * mat_B[187][3] +
                mat_A[166][0] * mat_B[195][3] +
                mat_A[166][1] * mat_B[203][3] +
                mat_A[166][2] * mat_B[211][3] +
                mat_A[166][3] * mat_B[219][3] +
                mat_A[167][0] * mat_B[227][3] +
                mat_A[167][1] * mat_B[235][3] +
                mat_A[167][2] * mat_B[243][3] +
                mat_A[167][3] * mat_B[251][3];
    mat_C[164][0] <=
                mat_A[160][0] * mat_B[4][0] +
                mat_A[160][1] * mat_B[12][0] +
                mat_A[160][2] * mat_B[20][0] +
                mat_A[160][3] * mat_B[28][0] +
                mat_A[161][0] * mat_B[36][0] +
                mat_A[161][1] * mat_B[44][0] +
                mat_A[161][2] * mat_B[52][0] +
                mat_A[161][3] * mat_B[60][0] +
                mat_A[162][0] * mat_B[68][0] +
                mat_A[162][1] * mat_B[76][0] +
                mat_A[162][2] * mat_B[84][0] +
                mat_A[162][3] * mat_B[92][0] +
                mat_A[163][0] * mat_B[100][0] +
                mat_A[163][1] * mat_B[108][0] +
                mat_A[163][2] * mat_B[116][0] +
                mat_A[163][3] * mat_B[124][0] +
                mat_A[164][0] * mat_B[132][0] +
                mat_A[164][1] * mat_B[140][0] +
                mat_A[164][2] * mat_B[148][0] +
                mat_A[164][3] * mat_B[156][0] +
                mat_A[165][0] * mat_B[164][0] +
                mat_A[165][1] * mat_B[172][0] +
                mat_A[165][2] * mat_B[180][0] +
                mat_A[165][3] * mat_B[188][0] +
                mat_A[166][0] * mat_B[196][0] +
                mat_A[166][1] * mat_B[204][0] +
                mat_A[166][2] * mat_B[212][0] +
                mat_A[166][3] * mat_B[220][0] +
                mat_A[167][0] * mat_B[228][0] +
                mat_A[167][1] * mat_B[236][0] +
                mat_A[167][2] * mat_B[244][0] +
                mat_A[167][3] * mat_B[252][0];
    mat_C[164][1] <=
                mat_A[160][0] * mat_B[4][1] +
                mat_A[160][1] * mat_B[12][1] +
                mat_A[160][2] * mat_B[20][1] +
                mat_A[160][3] * mat_B[28][1] +
                mat_A[161][0] * mat_B[36][1] +
                mat_A[161][1] * mat_B[44][1] +
                mat_A[161][2] * mat_B[52][1] +
                mat_A[161][3] * mat_B[60][1] +
                mat_A[162][0] * mat_B[68][1] +
                mat_A[162][1] * mat_B[76][1] +
                mat_A[162][2] * mat_B[84][1] +
                mat_A[162][3] * mat_B[92][1] +
                mat_A[163][0] * mat_B[100][1] +
                mat_A[163][1] * mat_B[108][1] +
                mat_A[163][2] * mat_B[116][1] +
                mat_A[163][3] * mat_B[124][1] +
                mat_A[164][0] * mat_B[132][1] +
                mat_A[164][1] * mat_B[140][1] +
                mat_A[164][2] * mat_B[148][1] +
                mat_A[164][3] * mat_B[156][1] +
                mat_A[165][0] * mat_B[164][1] +
                mat_A[165][1] * mat_B[172][1] +
                mat_A[165][2] * mat_B[180][1] +
                mat_A[165][3] * mat_B[188][1] +
                mat_A[166][0] * mat_B[196][1] +
                mat_A[166][1] * mat_B[204][1] +
                mat_A[166][2] * mat_B[212][1] +
                mat_A[166][3] * mat_B[220][1] +
                mat_A[167][0] * mat_B[228][1] +
                mat_A[167][1] * mat_B[236][1] +
                mat_A[167][2] * mat_B[244][1] +
                mat_A[167][3] * mat_B[252][1];
    mat_C[164][2] <=
                mat_A[160][0] * mat_B[4][2] +
                mat_A[160][1] * mat_B[12][2] +
                mat_A[160][2] * mat_B[20][2] +
                mat_A[160][3] * mat_B[28][2] +
                mat_A[161][0] * mat_B[36][2] +
                mat_A[161][1] * mat_B[44][2] +
                mat_A[161][2] * mat_B[52][2] +
                mat_A[161][3] * mat_B[60][2] +
                mat_A[162][0] * mat_B[68][2] +
                mat_A[162][1] * mat_B[76][2] +
                mat_A[162][2] * mat_B[84][2] +
                mat_A[162][3] * mat_B[92][2] +
                mat_A[163][0] * mat_B[100][2] +
                mat_A[163][1] * mat_B[108][2] +
                mat_A[163][2] * mat_B[116][2] +
                mat_A[163][3] * mat_B[124][2] +
                mat_A[164][0] * mat_B[132][2] +
                mat_A[164][1] * mat_B[140][2] +
                mat_A[164][2] * mat_B[148][2] +
                mat_A[164][3] * mat_B[156][2] +
                mat_A[165][0] * mat_B[164][2] +
                mat_A[165][1] * mat_B[172][2] +
                mat_A[165][2] * mat_B[180][2] +
                mat_A[165][3] * mat_B[188][2] +
                mat_A[166][0] * mat_B[196][2] +
                mat_A[166][1] * mat_B[204][2] +
                mat_A[166][2] * mat_B[212][2] +
                mat_A[166][3] * mat_B[220][2] +
                mat_A[167][0] * mat_B[228][2] +
                mat_A[167][1] * mat_B[236][2] +
                mat_A[167][2] * mat_B[244][2] +
                mat_A[167][3] * mat_B[252][2];
    mat_C[164][3] <=
                mat_A[160][0] * mat_B[4][3] +
                mat_A[160][1] * mat_B[12][3] +
                mat_A[160][2] * mat_B[20][3] +
                mat_A[160][3] * mat_B[28][3] +
                mat_A[161][0] * mat_B[36][3] +
                mat_A[161][1] * mat_B[44][3] +
                mat_A[161][2] * mat_B[52][3] +
                mat_A[161][3] * mat_B[60][3] +
                mat_A[162][0] * mat_B[68][3] +
                mat_A[162][1] * mat_B[76][3] +
                mat_A[162][2] * mat_B[84][3] +
                mat_A[162][3] * mat_B[92][3] +
                mat_A[163][0] * mat_B[100][3] +
                mat_A[163][1] * mat_B[108][3] +
                mat_A[163][2] * mat_B[116][3] +
                mat_A[163][3] * mat_B[124][3] +
                mat_A[164][0] * mat_B[132][3] +
                mat_A[164][1] * mat_B[140][3] +
                mat_A[164][2] * mat_B[148][3] +
                mat_A[164][3] * mat_B[156][3] +
                mat_A[165][0] * mat_B[164][3] +
                mat_A[165][1] * mat_B[172][3] +
                mat_A[165][2] * mat_B[180][3] +
                mat_A[165][3] * mat_B[188][3] +
                mat_A[166][0] * mat_B[196][3] +
                mat_A[166][1] * mat_B[204][3] +
                mat_A[166][2] * mat_B[212][3] +
                mat_A[166][3] * mat_B[220][3] +
                mat_A[167][0] * mat_B[228][3] +
                mat_A[167][1] * mat_B[236][3] +
                mat_A[167][2] * mat_B[244][3] +
                mat_A[167][3] * mat_B[252][3];
    mat_C[165][0] <=
                mat_A[160][0] * mat_B[5][0] +
                mat_A[160][1] * mat_B[13][0] +
                mat_A[160][2] * mat_B[21][0] +
                mat_A[160][3] * mat_B[29][0] +
                mat_A[161][0] * mat_B[37][0] +
                mat_A[161][1] * mat_B[45][0] +
                mat_A[161][2] * mat_B[53][0] +
                mat_A[161][3] * mat_B[61][0] +
                mat_A[162][0] * mat_B[69][0] +
                mat_A[162][1] * mat_B[77][0] +
                mat_A[162][2] * mat_B[85][0] +
                mat_A[162][3] * mat_B[93][0] +
                mat_A[163][0] * mat_B[101][0] +
                mat_A[163][1] * mat_B[109][0] +
                mat_A[163][2] * mat_B[117][0] +
                mat_A[163][3] * mat_B[125][0] +
                mat_A[164][0] * mat_B[133][0] +
                mat_A[164][1] * mat_B[141][0] +
                mat_A[164][2] * mat_B[149][0] +
                mat_A[164][3] * mat_B[157][0] +
                mat_A[165][0] * mat_B[165][0] +
                mat_A[165][1] * mat_B[173][0] +
                mat_A[165][2] * mat_B[181][0] +
                mat_A[165][3] * mat_B[189][0] +
                mat_A[166][0] * mat_B[197][0] +
                mat_A[166][1] * mat_B[205][0] +
                mat_A[166][2] * mat_B[213][0] +
                mat_A[166][3] * mat_B[221][0] +
                mat_A[167][0] * mat_B[229][0] +
                mat_A[167][1] * mat_B[237][0] +
                mat_A[167][2] * mat_B[245][0] +
                mat_A[167][3] * mat_B[253][0];
    mat_C[165][1] <=
                mat_A[160][0] * mat_B[5][1] +
                mat_A[160][1] * mat_B[13][1] +
                mat_A[160][2] * mat_B[21][1] +
                mat_A[160][3] * mat_B[29][1] +
                mat_A[161][0] * mat_B[37][1] +
                mat_A[161][1] * mat_B[45][1] +
                mat_A[161][2] * mat_B[53][1] +
                mat_A[161][3] * mat_B[61][1] +
                mat_A[162][0] * mat_B[69][1] +
                mat_A[162][1] * mat_B[77][1] +
                mat_A[162][2] * mat_B[85][1] +
                mat_A[162][3] * mat_B[93][1] +
                mat_A[163][0] * mat_B[101][1] +
                mat_A[163][1] * mat_B[109][1] +
                mat_A[163][2] * mat_B[117][1] +
                mat_A[163][3] * mat_B[125][1] +
                mat_A[164][0] * mat_B[133][1] +
                mat_A[164][1] * mat_B[141][1] +
                mat_A[164][2] * mat_B[149][1] +
                mat_A[164][3] * mat_B[157][1] +
                mat_A[165][0] * mat_B[165][1] +
                mat_A[165][1] * mat_B[173][1] +
                mat_A[165][2] * mat_B[181][1] +
                mat_A[165][3] * mat_B[189][1] +
                mat_A[166][0] * mat_B[197][1] +
                mat_A[166][1] * mat_B[205][1] +
                mat_A[166][2] * mat_B[213][1] +
                mat_A[166][3] * mat_B[221][1] +
                mat_A[167][0] * mat_B[229][1] +
                mat_A[167][1] * mat_B[237][1] +
                mat_A[167][2] * mat_B[245][1] +
                mat_A[167][3] * mat_B[253][1];
    mat_C[165][2] <=
                mat_A[160][0] * mat_B[5][2] +
                mat_A[160][1] * mat_B[13][2] +
                mat_A[160][2] * mat_B[21][2] +
                mat_A[160][3] * mat_B[29][2] +
                mat_A[161][0] * mat_B[37][2] +
                mat_A[161][1] * mat_B[45][2] +
                mat_A[161][2] * mat_B[53][2] +
                mat_A[161][3] * mat_B[61][2] +
                mat_A[162][0] * mat_B[69][2] +
                mat_A[162][1] * mat_B[77][2] +
                mat_A[162][2] * mat_B[85][2] +
                mat_A[162][3] * mat_B[93][2] +
                mat_A[163][0] * mat_B[101][2] +
                mat_A[163][1] * mat_B[109][2] +
                mat_A[163][2] * mat_B[117][2] +
                mat_A[163][3] * mat_B[125][2] +
                mat_A[164][0] * mat_B[133][2] +
                mat_A[164][1] * mat_B[141][2] +
                mat_A[164][2] * mat_B[149][2] +
                mat_A[164][3] * mat_B[157][2] +
                mat_A[165][0] * mat_B[165][2] +
                mat_A[165][1] * mat_B[173][2] +
                mat_A[165][2] * mat_B[181][2] +
                mat_A[165][3] * mat_B[189][2] +
                mat_A[166][0] * mat_B[197][2] +
                mat_A[166][1] * mat_B[205][2] +
                mat_A[166][2] * mat_B[213][2] +
                mat_A[166][3] * mat_B[221][2] +
                mat_A[167][0] * mat_B[229][2] +
                mat_A[167][1] * mat_B[237][2] +
                mat_A[167][2] * mat_B[245][2] +
                mat_A[167][3] * mat_B[253][2];
    mat_C[165][3] <=
                mat_A[160][0] * mat_B[5][3] +
                mat_A[160][1] * mat_B[13][3] +
                mat_A[160][2] * mat_B[21][3] +
                mat_A[160][3] * mat_B[29][3] +
                mat_A[161][0] * mat_B[37][3] +
                mat_A[161][1] * mat_B[45][3] +
                mat_A[161][2] * mat_B[53][3] +
                mat_A[161][3] * mat_B[61][3] +
                mat_A[162][0] * mat_B[69][3] +
                mat_A[162][1] * mat_B[77][3] +
                mat_A[162][2] * mat_B[85][3] +
                mat_A[162][3] * mat_B[93][3] +
                mat_A[163][0] * mat_B[101][3] +
                mat_A[163][1] * mat_B[109][3] +
                mat_A[163][2] * mat_B[117][3] +
                mat_A[163][3] * mat_B[125][3] +
                mat_A[164][0] * mat_B[133][3] +
                mat_A[164][1] * mat_B[141][3] +
                mat_A[164][2] * mat_B[149][3] +
                mat_A[164][3] * mat_B[157][3] +
                mat_A[165][0] * mat_B[165][3] +
                mat_A[165][1] * mat_B[173][3] +
                mat_A[165][2] * mat_B[181][3] +
                mat_A[165][3] * mat_B[189][3] +
                mat_A[166][0] * mat_B[197][3] +
                mat_A[166][1] * mat_B[205][3] +
                mat_A[166][2] * mat_B[213][3] +
                mat_A[166][3] * mat_B[221][3] +
                mat_A[167][0] * mat_B[229][3] +
                mat_A[167][1] * mat_B[237][3] +
                mat_A[167][2] * mat_B[245][3] +
                mat_A[167][3] * mat_B[253][3];
    mat_C[166][0] <=
                mat_A[160][0] * mat_B[6][0] +
                mat_A[160][1] * mat_B[14][0] +
                mat_A[160][2] * mat_B[22][0] +
                mat_A[160][3] * mat_B[30][0] +
                mat_A[161][0] * mat_B[38][0] +
                mat_A[161][1] * mat_B[46][0] +
                mat_A[161][2] * mat_B[54][0] +
                mat_A[161][3] * mat_B[62][0] +
                mat_A[162][0] * mat_B[70][0] +
                mat_A[162][1] * mat_B[78][0] +
                mat_A[162][2] * mat_B[86][0] +
                mat_A[162][3] * mat_B[94][0] +
                mat_A[163][0] * mat_B[102][0] +
                mat_A[163][1] * mat_B[110][0] +
                mat_A[163][2] * mat_B[118][0] +
                mat_A[163][3] * mat_B[126][0] +
                mat_A[164][0] * mat_B[134][0] +
                mat_A[164][1] * mat_B[142][0] +
                mat_A[164][2] * mat_B[150][0] +
                mat_A[164][3] * mat_B[158][0] +
                mat_A[165][0] * mat_B[166][0] +
                mat_A[165][1] * mat_B[174][0] +
                mat_A[165][2] * mat_B[182][0] +
                mat_A[165][3] * mat_B[190][0] +
                mat_A[166][0] * mat_B[198][0] +
                mat_A[166][1] * mat_B[206][0] +
                mat_A[166][2] * mat_B[214][0] +
                mat_A[166][3] * mat_B[222][0] +
                mat_A[167][0] * mat_B[230][0] +
                mat_A[167][1] * mat_B[238][0] +
                mat_A[167][2] * mat_B[246][0] +
                mat_A[167][3] * mat_B[254][0];
    mat_C[166][1] <=
                mat_A[160][0] * mat_B[6][1] +
                mat_A[160][1] * mat_B[14][1] +
                mat_A[160][2] * mat_B[22][1] +
                mat_A[160][3] * mat_B[30][1] +
                mat_A[161][0] * mat_B[38][1] +
                mat_A[161][1] * mat_B[46][1] +
                mat_A[161][2] * mat_B[54][1] +
                mat_A[161][3] * mat_B[62][1] +
                mat_A[162][0] * mat_B[70][1] +
                mat_A[162][1] * mat_B[78][1] +
                mat_A[162][2] * mat_B[86][1] +
                mat_A[162][3] * mat_B[94][1] +
                mat_A[163][0] * mat_B[102][1] +
                mat_A[163][1] * mat_B[110][1] +
                mat_A[163][2] * mat_B[118][1] +
                mat_A[163][3] * mat_B[126][1] +
                mat_A[164][0] * mat_B[134][1] +
                mat_A[164][1] * mat_B[142][1] +
                mat_A[164][2] * mat_B[150][1] +
                mat_A[164][3] * mat_B[158][1] +
                mat_A[165][0] * mat_B[166][1] +
                mat_A[165][1] * mat_B[174][1] +
                mat_A[165][2] * mat_B[182][1] +
                mat_A[165][3] * mat_B[190][1] +
                mat_A[166][0] * mat_B[198][1] +
                mat_A[166][1] * mat_B[206][1] +
                mat_A[166][2] * mat_B[214][1] +
                mat_A[166][3] * mat_B[222][1] +
                mat_A[167][0] * mat_B[230][1] +
                mat_A[167][1] * mat_B[238][1] +
                mat_A[167][2] * mat_B[246][1] +
                mat_A[167][3] * mat_B[254][1];
    mat_C[166][2] <=
                mat_A[160][0] * mat_B[6][2] +
                mat_A[160][1] * mat_B[14][2] +
                mat_A[160][2] * mat_B[22][2] +
                mat_A[160][3] * mat_B[30][2] +
                mat_A[161][0] * mat_B[38][2] +
                mat_A[161][1] * mat_B[46][2] +
                mat_A[161][2] * mat_B[54][2] +
                mat_A[161][3] * mat_B[62][2] +
                mat_A[162][0] * mat_B[70][2] +
                mat_A[162][1] * mat_B[78][2] +
                mat_A[162][2] * mat_B[86][2] +
                mat_A[162][3] * mat_B[94][2] +
                mat_A[163][0] * mat_B[102][2] +
                mat_A[163][1] * mat_B[110][2] +
                mat_A[163][2] * mat_B[118][2] +
                mat_A[163][3] * mat_B[126][2] +
                mat_A[164][0] * mat_B[134][2] +
                mat_A[164][1] * mat_B[142][2] +
                mat_A[164][2] * mat_B[150][2] +
                mat_A[164][3] * mat_B[158][2] +
                mat_A[165][0] * mat_B[166][2] +
                mat_A[165][1] * mat_B[174][2] +
                mat_A[165][2] * mat_B[182][2] +
                mat_A[165][3] * mat_B[190][2] +
                mat_A[166][0] * mat_B[198][2] +
                mat_A[166][1] * mat_B[206][2] +
                mat_A[166][2] * mat_B[214][2] +
                mat_A[166][3] * mat_B[222][2] +
                mat_A[167][0] * mat_B[230][2] +
                mat_A[167][1] * mat_B[238][2] +
                mat_A[167][2] * mat_B[246][2] +
                mat_A[167][3] * mat_B[254][2];
    mat_C[166][3] <=
                mat_A[160][0] * mat_B[6][3] +
                mat_A[160][1] * mat_B[14][3] +
                mat_A[160][2] * mat_B[22][3] +
                mat_A[160][3] * mat_B[30][3] +
                mat_A[161][0] * mat_B[38][3] +
                mat_A[161][1] * mat_B[46][3] +
                mat_A[161][2] * mat_B[54][3] +
                mat_A[161][3] * mat_B[62][3] +
                mat_A[162][0] * mat_B[70][3] +
                mat_A[162][1] * mat_B[78][3] +
                mat_A[162][2] * mat_B[86][3] +
                mat_A[162][3] * mat_B[94][3] +
                mat_A[163][0] * mat_B[102][3] +
                mat_A[163][1] * mat_B[110][3] +
                mat_A[163][2] * mat_B[118][3] +
                mat_A[163][3] * mat_B[126][3] +
                mat_A[164][0] * mat_B[134][3] +
                mat_A[164][1] * mat_B[142][3] +
                mat_A[164][2] * mat_B[150][3] +
                mat_A[164][3] * mat_B[158][3] +
                mat_A[165][0] * mat_B[166][3] +
                mat_A[165][1] * mat_B[174][3] +
                mat_A[165][2] * mat_B[182][3] +
                mat_A[165][3] * mat_B[190][3] +
                mat_A[166][0] * mat_B[198][3] +
                mat_A[166][1] * mat_B[206][3] +
                mat_A[166][2] * mat_B[214][3] +
                mat_A[166][3] * mat_B[222][3] +
                mat_A[167][0] * mat_B[230][3] +
                mat_A[167][1] * mat_B[238][3] +
                mat_A[167][2] * mat_B[246][3] +
                mat_A[167][3] * mat_B[254][3];
    mat_C[167][0] <=
                mat_A[160][0] * mat_B[7][0] +
                mat_A[160][1] * mat_B[15][0] +
                mat_A[160][2] * mat_B[23][0] +
                mat_A[160][3] * mat_B[31][0] +
                mat_A[161][0] * mat_B[39][0] +
                mat_A[161][1] * mat_B[47][0] +
                mat_A[161][2] * mat_B[55][0] +
                mat_A[161][3] * mat_B[63][0] +
                mat_A[162][0] * mat_B[71][0] +
                mat_A[162][1] * mat_B[79][0] +
                mat_A[162][2] * mat_B[87][0] +
                mat_A[162][3] * mat_B[95][0] +
                mat_A[163][0] * mat_B[103][0] +
                mat_A[163][1] * mat_B[111][0] +
                mat_A[163][2] * mat_B[119][0] +
                mat_A[163][3] * mat_B[127][0] +
                mat_A[164][0] * mat_B[135][0] +
                mat_A[164][1] * mat_B[143][0] +
                mat_A[164][2] * mat_B[151][0] +
                mat_A[164][3] * mat_B[159][0] +
                mat_A[165][0] * mat_B[167][0] +
                mat_A[165][1] * mat_B[175][0] +
                mat_A[165][2] * mat_B[183][0] +
                mat_A[165][3] * mat_B[191][0] +
                mat_A[166][0] * mat_B[199][0] +
                mat_A[166][1] * mat_B[207][0] +
                mat_A[166][2] * mat_B[215][0] +
                mat_A[166][3] * mat_B[223][0] +
                mat_A[167][0] * mat_B[231][0] +
                mat_A[167][1] * mat_B[239][0] +
                mat_A[167][2] * mat_B[247][0] +
                mat_A[167][3] * mat_B[255][0];
    mat_C[167][1] <=
                mat_A[160][0] * mat_B[7][1] +
                mat_A[160][1] * mat_B[15][1] +
                mat_A[160][2] * mat_B[23][1] +
                mat_A[160][3] * mat_B[31][1] +
                mat_A[161][0] * mat_B[39][1] +
                mat_A[161][1] * mat_B[47][1] +
                mat_A[161][2] * mat_B[55][1] +
                mat_A[161][3] * mat_B[63][1] +
                mat_A[162][0] * mat_B[71][1] +
                mat_A[162][1] * mat_B[79][1] +
                mat_A[162][2] * mat_B[87][1] +
                mat_A[162][3] * mat_B[95][1] +
                mat_A[163][0] * mat_B[103][1] +
                mat_A[163][1] * mat_B[111][1] +
                mat_A[163][2] * mat_B[119][1] +
                mat_A[163][3] * mat_B[127][1] +
                mat_A[164][0] * mat_B[135][1] +
                mat_A[164][1] * mat_B[143][1] +
                mat_A[164][2] * mat_B[151][1] +
                mat_A[164][3] * mat_B[159][1] +
                mat_A[165][0] * mat_B[167][1] +
                mat_A[165][1] * mat_B[175][1] +
                mat_A[165][2] * mat_B[183][1] +
                mat_A[165][3] * mat_B[191][1] +
                mat_A[166][0] * mat_B[199][1] +
                mat_A[166][1] * mat_B[207][1] +
                mat_A[166][2] * mat_B[215][1] +
                mat_A[166][3] * mat_B[223][1] +
                mat_A[167][0] * mat_B[231][1] +
                mat_A[167][1] * mat_B[239][1] +
                mat_A[167][2] * mat_B[247][1] +
                mat_A[167][3] * mat_B[255][1];
    mat_C[167][2] <=
                mat_A[160][0] * mat_B[7][2] +
                mat_A[160][1] * mat_B[15][2] +
                mat_A[160][2] * mat_B[23][2] +
                mat_A[160][3] * mat_B[31][2] +
                mat_A[161][0] * mat_B[39][2] +
                mat_A[161][1] * mat_B[47][2] +
                mat_A[161][2] * mat_B[55][2] +
                mat_A[161][3] * mat_B[63][2] +
                mat_A[162][0] * mat_B[71][2] +
                mat_A[162][1] * mat_B[79][2] +
                mat_A[162][2] * mat_B[87][2] +
                mat_A[162][3] * mat_B[95][2] +
                mat_A[163][0] * mat_B[103][2] +
                mat_A[163][1] * mat_B[111][2] +
                mat_A[163][2] * mat_B[119][2] +
                mat_A[163][3] * mat_B[127][2] +
                mat_A[164][0] * mat_B[135][2] +
                mat_A[164][1] * mat_B[143][2] +
                mat_A[164][2] * mat_B[151][2] +
                mat_A[164][3] * mat_B[159][2] +
                mat_A[165][0] * mat_B[167][2] +
                mat_A[165][1] * mat_B[175][2] +
                mat_A[165][2] * mat_B[183][2] +
                mat_A[165][3] * mat_B[191][2] +
                mat_A[166][0] * mat_B[199][2] +
                mat_A[166][1] * mat_B[207][2] +
                mat_A[166][2] * mat_B[215][2] +
                mat_A[166][3] * mat_B[223][2] +
                mat_A[167][0] * mat_B[231][2] +
                mat_A[167][1] * mat_B[239][2] +
                mat_A[167][2] * mat_B[247][2] +
                mat_A[167][3] * mat_B[255][2];
    mat_C[167][3] <=
                mat_A[160][0] * mat_B[7][3] +
                mat_A[160][1] * mat_B[15][3] +
                mat_A[160][2] * mat_B[23][3] +
                mat_A[160][3] * mat_B[31][3] +
                mat_A[161][0] * mat_B[39][3] +
                mat_A[161][1] * mat_B[47][3] +
                mat_A[161][2] * mat_B[55][3] +
                mat_A[161][3] * mat_B[63][3] +
                mat_A[162][0] * mat_B[71][3] +
                mat_A[162][1] * mat_B[79][3] +
                mat_A[162][2] * mat_B[87][3] +
                mat_A[162][3] * mat_B[95][3] +
                mat_A[163][0] * mat_B[103][3] +
                mat_A[163][1] * mat_B[111][3] +
                mat_A[163][2] * mat_B[119][3] +
                mat_A[163][3] * mat_B[127][3] +
                mat_A[164][0] * mat_B[135][3] +
                mat_A[164][1] * mat_B[143][3] +
                mat_A[164][2] * mat_B[151][3] +
                mat_A[164][3] * mat_B[159][3] +
                mat_A[165][0] * mat_B[167][3] +
                mat_A[165][1] * mat_B[175][3] +
                mat_A[165][2] * mat_B[183][3] +
                mat_A[165][3] * mat_B[191][3] +
                mat_A[166][0] * mat_B[199][3] +
                mat_A[166][1] * mat_B[207][3] +
                mat_A[166][2] * mat_B[215][3] +
                mat_A[166][3] * mat_B[223][3] +
                mat_A[167][0] * mat_B[231][3] +
                mat_A[167][1] * mat_B[239][3] +
                mat_A[167][2] * mat_B[247][3] +
                mat_A[167][3] * mat_B[255][3];
    mat_C[168][0] <=
                mat_A[168][0] * mat_B[0][0] +
                mat_A[168][1] * mat_B[8][0] +
                mat_A[168][2] * mat_B[16][0] +
                mat_A[168][3] * mat_B[24][0] +
                mat_A[169][0] * mat_B[32][0] +
                mat_A[169][1] * mat_B[40][0] +
                mat_A[169][2] * mat_B[48][0] +
                mat_A[169][3] * mat_B[56][0] +
                mat_A[170][0] * mat_B[64][0] +
                mat_A[170][1] * mat_B[72][0] +
                mat_A[170][2] * mat_B[80][0] +
                mat_A[170][3] * mat_B[88][0] +
                mat_A[171][0] * mat_B[96][0] +
                mat_A[171][1] * mat_B[104][0] +
                mat_A[171][2] * mat_B[112][0] +
                mat_A[171][3] * mat_B[120][0] +
                mat_A[172][0] * mat_B[128][0] +
                mat_A[172][1] * mat_B[136][0] +
                mat_A[172][2] * mat_B[144][0] +
                mat_A[172][3] * mat_B[152][0] +
                mat_A[173][0] * mat_B[160][0] +
                mat_A[173][1] * mat_B[168][0] +
                mat_A[173][2] * mat_B[176][0] +
                mat_A[173][3] * mat_B[184][0] +
                mat_A[174][0] * mat_B[192][0] +
                mat_A[174][1] * mat_B[200][0] +
                mat_A[174][2] * mat_B[208][0] +
                mat_A[174][3] * mat_B[216][0] +
                mat_A[175][0] * mat_B[224][0] +
                mat_A[175][1] * mat_B[232][0] +
                mat_A[175][2] * mat_B[240][0] +
                mat_A[175][3] * mat_B[248][0];
    mat_C[168][1] <=
                mat_A[168][0] * mat_B[0][1] +
                mat_A[168][1] * mat_B[8][1] +
                mat_A[168][2] * mat_B[16][1] +
                mat_A[168][3] * mat_B[24][1] +
                mat_A[169][0] * mat_B[32][1] +
                mat_A[169][1] * mat_B[40][1] +
                mat_A[169][2] * mat_B[48][1] +
                mat_A[169][3] * mat_B[56][1] +
                mat_A[170][0] * mat_B[64][1] +
                mat_A[170][1] * mat_B[72][1] +
                mat_A[170][2] * mat_B[80][1] +
                mat_A[170][3] * mat_B[88][1] +
                mat_A[171][0] * mat_B[96][1] +
                mat_A[171][1] * mat_B[104][1] +
                mat_A[171][2] * mat_B[112][1] +
                mat_A[171][3] * mat_B[120][1] +
                mat_A[172][0] * mat_B[128][1] +
                mat_A[172][1] * mat_B[136][1] +
                mat_A[172][2] * mat_B[144][1] +
                mat_A[172][3] * mat_B[152][1] +
                mat_A[173][0] * mat_B[160][1] +
                mat_A[173][1] * mat_B[168][1] +
                mat_A[173][2] * mat_B[176][1] +
                mat_A[173][3] * mat_B[184][1] +
                mat_A[174][0] * mat_B[192][1] +
                mat_A[174][1] * mat_B[200][1] +
                mat_A[174][2] * mat_B[208][1] +
                mat_A[174][3] * mat_B[216][1] +
                mat_A[175][0] * mat_B[224][1] +
                mat_A[175][1] * mat_B[232][1] +
                mat_A[175][2] * mat_B[240][1] +
                mat_A[175][3] * mat_B[248][1];
    mat_C[168][2] <=
                mat_A[168][0] * mat_B[0][2] +
                mat_A[168][1] * mat_B[8][2] +
                mat_A[168][2] * mat_B[16][2] +
                mat_A[168][3] * mat_B[24][2] +
                mat_A[169][0] * mat_B[32][2] +
                mat_A[169][1] * mat_B[40][2] +
                mat_A[169][2] * mat_B[48][2] +
                mat_A[169][3] * mat_B[56][2] +
                mat_A[170][0] * mat_B[64][2] +
                mat_A[170][1] * mat_B[72][2] +
                mat_A[170][2] * mat_B[80][2] +
                mat_A[170][3] * mat_B[88][2] +
                mat_A[171][0] * mat_B[96][2] +
                mat_A[171][1] * mat_B[104][2] +
                mat_A[171][2] * mat_B[112][2] +
                mat_A[171][3] * mat_B[120][2] +
                mat_A[172][0] * mat_B[128][2] +
                mat_A[172][1] * mat_B[136][2] +
                mat_A[172][2] * mat_B[144][2] +
                mat_A[172][3] * mat_B[152][2] +
                mat_A[173][0] * mat_B[160][2] +
                mat_A[173][1] * mat_B[168][2] +
                mat_A[173][2] * mat_B[176][2] +
                mat_A[173][3] * mat_B[184][2] +
                mat_A[174][0] * mat_B[192][2] +
                mat_A[174][1] * mat_B[200][2] +
                mat_A[174][2] * mat_B[208][2] +
                mat_A[174][3] * mat_B[216][2] +
                mat_A[175][0] * mat_B[224][2] +
                mat_A[175][1] * mat_B[232][2] +
                mat_A[175][2] * mat_B[240][2] +
                mat_A[175][3] * mat_B[248][2];
    mat_C[168][3] <=
                mat_A[168][0] * mat_B[0][3] +
                mat_A[168][1] * mat_B[8][3] +
                mat_A[168][2] * mat_B[16][3] +
                mat_A[168][3] * mat_B[24][3] +
                mat_A[169][0] * mat_B[32][3] +
                mat_A[169][1] * mat_B[40][3] +
                mat_A[169][2] * mat_B[48][3] +
                mat_A[169][3] * mat_B[56][3] +
                mat_A[170][0] * mat_B[64][3] +
                mat_A[170][1] * mat_B[72][3] +
                mat_A[170][2] * mat_B[80][3] +
                mat_A[170][3] * mat_B[88][3] +
                mat_A[171][0] * mat_B[96][3] +
                mat_A[171][1] * mat_B[104][3] +
                mat_A[171][2] * mat_B[112][3] +
                mat_A[171][3] * mat_B[120][3] +
                mat_A[172][0] * mat_B[128][3] +
                mat_A[172][1] * mat_B[136][3] +
                mat_A[172][2] * mat_B[144][3] +
                mat_A[172][3] * mat_B[152][3] +
                mat_A[173][0] * mat_B[160][3] +
                mat_A[173][1] * mat_B[168][3] +
                mat_A[173][2] * mat_B[176][3] +
                mat_A[173][3] * mat_B[184][3] +
                mat_A[174][0] * mat_B[192][3] +
                mat_A[174][1] * mat_B[200][3] +
                mat_A[174][2] * mat_B[208][3] +
                mat_A[174][3] * mat_B[216][3] +
                mat_A[175][0] * mat_B[224][3] +
                mat_A[175][1] * mat_B[232][3] +
                mat_A[175][2] * mat_B[240][3] +
                mat_A[175][3] * mat_B[248][3];
    mat_C[169][0] <=
                mat_A[168][0] * mat_B[1][0] +
                mat_A[168][1] * mat_B[9][0] +
                mat_A[168][2] * mat_B[17][0] +
                mat_A[168][3] * mat_B[25][0] +
                mat_A[169][0] * mat_B[33][0] +
                mat_A[169][1] * mat_B[41][0] +
                mat_A[169][2] * mat_B[49][0] +
                mat_A[169][3] * mat_B[57][0] +
                mat_A[170][0] * mat_B[65][0] +
                mat_A[170][1] * mat_B[73][0] +
                mat_A[170][2] * mat_B[81][0] +
                mat_A[170][3] * mat_B[89][0] +
                mat_A[171][0] * mat_B[97][0] +
                mat_A[171][1] * mat_B[105][0] +
                mat_A[171][2] * mat_B[113][0] +
                mat_A[171][3] * mat_B[121][0] +
                mat_A[172][0] * mat_B[129][0] +
                mat_A[172][1] * mat_B[137][0] +
                mat_A[172][2] * mat_B[145][0] +
                mat_A[172][3] * mat_B[153][0] +
                mat_A[173][0] * mat_B[161][0] +
                mat_A[173][1] * mat_B[169][0] +
                mat_A[173][2] * mat_B[177][0] +
                mat_A[173][3] * mat_B[185][0] +
                mat_A[174][0] * mat_B[193][0] +
                mat_A[174][1] * mat_B[201][0] +
                mat_A[174][2] * mat_B[209][0] +
                mat_A[174][3] * mat_B[217][0] +
                mat_A[175][0] * mat_B[225][0] +
                mat_A[175][1] * mat_B[233][0] +
                mat_A[175][2] * mat_B[241][0] +
                mat_A[175][3] * mat_B[249][0];
    mat_C[169][1] <=
                mat_A[168][0] * mat_B[1][1] +
                mat_A[168][1] * mat_B[9][1] +
                mat_A[168][2] * mat_B[17][1] +
                mat_A[168][3] * mat_B[25][1] +
                mat_A[169][0] * mat_B[33][1] +
                mat_A[169][1] * mat_B[41][1] +
                mat_A[169][2] * mat_B[49][1] +
                mat_A[169][3] * mat_B[57][1] +
                mat_A[170][0] * mat_B[65][1] +
                mat_A[170][1] * mat_B[73][1] +
                mat_A[170][2] * mat_B[81][1] +
                mat_A[170][3] * mat_B[89][1] +
                mat_A[171][0] * mat_B[97][1] +
                mat_A[171][1] * mat_B[105][1] +
                mat_A[171][2] * mat_B[113][1] +
                mat_A[171][3] * mat_B[121][1] +
                mat_A[172][0] * mat_B[129][1] +
                mat_A[172][1] * mat_B[137][1] +
                mat_A[172][2] * mat_B[145][1] +
                mat_A[172][3] * mat_B[153][1] +
                mat_A[173][0] * mat_B[161][1] +
                mat_A[173][1] * mat_B[169][1] +
                mat_A[173][2] * mat_B[177][1] +
                mat_A[173][3] * mat_B[185][1] +
                mat_A[174][0] * mat_B[193][1] +
                mat_A[174][1] * mat_B[201][1] +
                mat_A[174][2] * mat_B[209][1] +
                mat_A[174][3] * mat_B[217][1] +
                mat_A[175][0] * mat_B[225][1] +
                mat_A[175][1] * mat_B[233][1] +
                mat_A[175][2] * mat_B[241][1] +
                mat_A[175][3] * mat_B[249][1];
    mat_C[169][2] <=
                mat_A[168][0] * mat_B[1][2] +
                mat_A[168][1] * mat_B[9][2] +
                mat_A[168][2] * mat_B[17][2] +
                mat_A[168][3] * mat_B[25][2] +
                mat_A[169][0] * mat_B[33][2] +
                mat_A[169][1] * mat_B[41][2] +
                mat_A[169][2] * mat_B[49][2] +
                mat_A[169][3] * mat_B[57][2] +
                mat_A[170][0] * mat_B[65][2] +
                mat_A[170][1] * mat_B[73][2] +
                mat_A[170][2] * mat_B[81][2] +
                mat_A[170][3] * mat_B[89][2] +
                mat_A[171][0] * mat_B[97][2] +
                mat_A[171][1] * mat_B[105][2] +
                mat_A[171][2] * mat_B[113][2] +
                mat_A[171][3] * mat_B[121][2] +
                mat_A[172][0] * mat_B[129][2] +
                mat_A[172][1] * mat_B[137][2] +
                mat_A[172][2] * mat_B[145][2] +
                mat_A[172][3] * mat_B[153][2] +
                mat_A[173][0] * mat_B[161][2] +
                mat_A[173][1] * mat_B[169][2] +
                mat_A[173][2] * mat_B[177][2] +
                mat_A[173][3] * mat_B[185][2] +
                mat_A[174][0] * mat_B[193][2] +
                mat_A[174][1] * mat_B[201][2] +
                mat_A[174][2] * mat_B[209][2] +
                mat_A[174][3] * mat_B[217][2] +
                mat_A[175][0] * mat_B[225][2] +
                mat_A[175][1] * mat_B[233][2] +
                mat_A[175][2] * mat_B[241][2] +
                mat_A[175][3] * mat_B[249][2];
    mat_C[169][3] <=
                mat_A[168][0] * mat_B[1][3] +
                mat_A[168][1] * mat_B[9][3] +
                mat_A[168][2] * mat_B[17][3] +
                mat_A[168][3] * mat_B[25][3] +
                mat_A[169][0] * mat_B[33][3] +
                mat_A[169][1] * mat_B[41][3] +
                mat_A[169][2] * mat_B[49][3] +
                mat_A[169][3] * mat_B[57][3] +
                mat_A[170][0] * mat_B[65][3] +
                mat_A[170][1] * mat_B[73][3] +
                mat_A[170][2] * mat_B[81][3] +
                mat_A[170][3] * mat_B[89][3] +
                mat_A[171][0] * mat_B[97][3] +
                mat_A[171][1] * mat_B[105][3] +
                mat_A[171][2] * mat_B[113][3] +
                mat_A[171][3] * mat_B[121][3] +
                mat_A[172][0] * mat_B[129][3] +
                mat_A[172][1] * mat_B[137][3] +
                mat_A[172][2] * mat_B[145][3] +
                mat_A[172][3] * mat_B[153][3] +
                mat_A[173][0] * mat_B[161][3] +
                mat_A[173][1] * mat_B[169][3] +
                mat_A[173][2] * mat_B[177][3] +
                mat_A[173][3] * mat_B[185][3] +
                mat_A[174][0] * mat_B[193][3] +
                mat_A[174][1] * mat_B[201][3] +
                mat_A[174][2] * mat_B[209][3] +
                mat_A[174][3] * mat_B[217][3] +
                mat_A[175][0] * mat_B[225][3] +
                mat_A[175][1] * mat_B[233][3] +
                mat_A[175][2] * mat_B[241][3] +
                mat_A[175][3] * mat_B[249][3];
    mat_C[170][0] <=
                mat_A[168][0] * mat_B[2][0] +
                mat_A[168][1] * mat_B[10][0] +
                mat_A[168][2] * mat_B[18][0] +
                mat_A[168][3] * mat_B[26][0] +
                mat_A[169][0] * mat_B[34][0] +
                mat_A[169][1] * mat_B[42][0] +
                mat_A[169][2] * mat_B[50][0] +
                mat_A[169][3] * mat_B[58][0] +
                mat_A[170][0] * mat_B[66][0] +
                mat_A[170][1] * mat_B[74][0] +
                mat_A[170][2] * mat_B[82][0] +
                mat_A[170][3] * mat_B[90][0] +
                mat_A[171][0] * mat_B[98][0] +
                mat_A[171][1] * mat_B[106][0] +
                mat_A[171][2] * mat_B[114][0] +
                mat_A[171][3] * mat_B[122][0] +
                mat_A[172][0] * mat_B[130][0] +
                mat_A[172][1] * mat_B[138][0] +
                mat_A[172][2] * mat_B[146][0] +
                mat_A[172][3] * mat_B[154][0] +
                mat_A[173][0] * mat_B[162][0] +
                mat_A[173][1] * mat_B[170][0] +
                mat_A[173][2] * mat_B[178][0] +
                mat_A[173][3] * mat_B[186][0] +
                mat_A[174][0] * mat_B[194][0] +
                mat_A[174][1] * mat_B[202][0] +
                mat_A[174][2] * mat_B[210][0] +
                mat_A[174][3] * mat_B[218][0] +
                mat_A[175][0] * mat_B[226][0] +
                mat_A[175][1] * mat_B[234][0] +
                mat_A[175][2] * mat_B[242][0] +
                mat_A[175][3] * mat_B[250][0];
    mat_C[170][1] <=
                mat_A[168][0] * mat_B[2][1] +
                mat_A[168][1] * mat_B[10][1] +
                mat_A[168][2] * mat_B[18][1] +
                mat_A[168][3] * mat_B[26][1] +
                mat_A[169][0] * mat_B[34][1] +
                mat_A[169][1] * mat_B[42][1] +
                mat_A[169][2] * mat_B[50][1] +
                mat_A[169][3] * mat_B[58][1] +
                mat_A[170][0] * mat_B[66][1] +
                mat_A[170][1] * mat_B[74][1] +
                mat_A[170][2] * mat_B[82][1] +
                mat_A[170][3] * mat_B[90][1] +
                mat_A[171][0] * mat_B[98][1] +
                mat_A[171][1] * mat_B[106][1] +
                mat_A[171][2] * mat_B[114][1] +
                mat_A[171][3] * mat_B[122][1] +
                mat_A[172][0] * mat_B[130][1] +
                mat_A[172][1] * mat_B[138][1] +
                mat_A[172][2] * mat_B[146][1] +
                mat_A[172][3] * mat_B[154][1] +
                mat_A[173][0] * mat_B[162][1] +
                mat_A[173][1] * mat_B[170][1] +
                mat_A[173][2] * mat_B[178][1] +
                mat_A[173][3] * mat_B[186][1] +
                mat_A[174][0] * mat_B[194][1] +
                mat_A[174][1] * mat_B[202][1] +
                mat_A[174][2] * mat_B[210][1] +
                mat_A[174][3] * mat_B[218][1] +
                mat_A[175][0] * mat_B[226][1] +
                mat_A[175][1] * mat_B[234][1] +
                mat_A[175][2] * mat_B[242][1] +
                mat_A[175][3] * mat_B[250][1];
    mat_C[170][2] <=
                mat_A[168][0] * mat_B[2][2] +
                mat_A[168][1] * mat_B[10][2] +
                mat_A[168][2] * mat_B[18][2] +
                mat_A[168][3] * mat_B[26][2] +
                mat_A[169][0] * mat_B[34][2] +
                mat_A[169][1] * mat_B[42][2] +
                mat_A[169][2] * mat_B[50][2] +
                mat_A[169][3] * mat_B[58][2] +
                mat_A[170][0] * mat_B[66][2] +
                mat_A[170][1] * mat_B[74][2] +
                mat_A[170][2] * mat_B[82][2] +
                mat_A[170][3] * mat_B[90][2] +
                mat_A[171][0] * mat_B[98][2] +
                mat_A[171][1] * mat_B[106][2] +
                mat_A[171][2] * mat_B[114][2] +
                mat_A[171][3] * mat_B[122][2] +
                mat_A[172][0] * mat_B[130][2] +
                mat_A[172][1] * mat_B[138][2] +
                mat_A[172][2] * mat_B[146][2] +
                mat_A[172][3] * mat_B[154][2] +
                mat_A[173][0] * mat_B[162][2] +
                mat_A[173][1] * mat_B[170][2] +
                mat_A[173][2] * mat_B[178][2] +
                mat_A[173][3] * mat_B[186][2] +
                mat_A[174][0] * mat_B[194][2] +
                mat_A[174][1] * mat_B[202][2] +
                mat_A[174][2] * mat_B[210][2] +
                mat_A[174][3] * mat_B[218][2] +
                mat_A[175][0] * mat_B[226][2] +
                mat_A[175][1] * mat_B[234][2] +
                mat_A[175][2] * mat_B[242][2] +
                mat_A[175][3] * mat_B[250][2];
    mat_C[170][3] <=
                mat_A[168][0] * mat_B[2][3] +
                mat_A[168][1] * mat_B[10][3] +
                mat_A[168][2] * mat_B[18][3] +
                mat_A[168][3] * mat_B[26][3] +
                mat_A[169][0] * mat_B[34][3] +
                mat_A[169][1] * mat_B[42][3] +
                mat_A[169][2] * mat_B[50][3] +
                mat_A[169][3] * mat_B[58][3] +
                mat_A[170][0] * mat_B[66][3] +
                mat_A[170][1] * mat_B[74][3] +
                mat_A[170][2] * mat_B[82][3] +
                mat_A[170][3] * mat_B[90][3] +
                mat_A[171][0] * mat_B[98][3] +
                mat_A[171][1] * mat_B[106][3] +
                mat_A[171][2] * mat_B[114][3] +
                mat_A[171][3] * mat_B[122][3] +
                mat_A[172][0] * mat_B[130][3] +
                mat_A[172][1] * mat_B[138][3] +
                mat_A[172][2] * mat_B[146][3] +
                mat_A[172][3] * mat_B[154][3] +
                mat_A[173][0] * mat_B[162][3] +
                mat_A[173][1] * mat_B[170][3] +
                mat_A[173][2] * mat_B[178][3] +
                mat_A[173][3] * mat_B[186][3] +
                mat_A[174][0] * mat_B[194][3] +
                mat_A[174][1] * mat_B[202][3] +
                mat_A[174][2] * mat_B[210][3] +
                mat_A[174][3] * mat_B[218][3] +
                mat_A[175][0] * mat_B[226][3] +
                mat_A[175][1] * mat_B[234][3] +
                mat_A[175][2] * mat_B[242][3] +
                mat_A[175][3] * mat_B[250][3];
    mat_C[171][0] <=
                mat_A[168][0] * mat_B[3][0] +
                mat_A[168][1] * mat_B[11][0] +
                mat_A[168][2] * mat_B[19][0] +
                mat_A[168][3] * mat_B[27][0] +
                mat_A[169][0] * mat_B[35][0] +
                mat_A[169][1] * mat_B[43][0] +
                mat_A[169][2] * mat_B[51][0] +
                mat_A[169][3] * mat_B[59][0] +
                mat_A[170][0] * mat_B[67][0] +
                mat_A[170][1] * mat_B[75][0] +
                mat_A[170][2] * mat_B[83][0] +
                mat_A[170][3] * mat_B[91][0] +
                mat_A[171][0] * mat_B[99][0] +
                mat_A[171][1] * mat_B[107][0] +
                mat_A[171][2] * mat_B[115][0] +
                mat_A[171][3] * mat_B[123][0] +
                mat_A[172][0] * mat_B[131][0] +
                mat_A[172][1] * mat_B[139][0] +
                mat_A[172][2] * mat_B[147][0] +
                mat_A[172][3] * mat_B[155][0] +
                mat_A[173][0] * mat_B[163][0] +
                mat_A[173][1] * mat_B[171][0] +
                mat_A[173][2] * mat_B[179][0] +
                mat_A[173][3] * mat_B[187][0] +
                mat_A[174][0] * mat_B[195][0] +
                mat_A[174][1] * mat_B[203][0] +
                mat_A[174][2] * mat_B[211][0] +
                mat_A[174][3] * mat_B[219][0] +
                mat_A[175][0] * mat_B[227][0] +
                mat_A[175][1] * mat_B[235][0] +
                mat_A[175][2] * mat_B[243][0] +
                mat_A[175][3] * mat_B[251][0];
    mat_C[171][1] <=
                mat_A[168][0] * mat_B[3][1] +
                mat_A[168][1] * mat_B[11][1] +
                mat_A[168][2] * mat_B[19][1] +
                mat_A[168][3] * mat_B[27][1] +
                mat_A[169][0] * mat_B[35][1] +
                mat_A[169][1] * mat_B[43][1] +
                mat_A[169][2] * mat_B[51][1] +
                mat_A[169][3] * mat_B[59][1] +
                mat_A[170][0] * mat_B[67][1] +
                mat_A[170][1] * mat_B[75][1] +
                mat_A[170][2] * mat_B[83][1] +
                mat_A[170][3] * mat_B[91][1] +
                mat_A[171][0] * mat_B[99][1] +
                mat_A[171][1] * mat_B[107][1] +
                mat_A[171][2] * mat_B[115][1] +
                mat_A[171][3] * mat_B[123][1] +
                mat_A[172][0] * mat_B[131][1] +
                mat_A[172][1] * mat_B[139][1] +
                mat_A[172][2] * mat_B[147][1] +
                mat_A[172][3] * mat_B[155][1] +
                mat_A[173][0] * mat_B[163][1] +
                mat_A[173][1] * mat_B[171][1] +
                mat_A[173][2] * mat_B[179][1] +
                mat_A[173][3] * mat_B[187][1] +
                mat_A[174][0] * mat_B[195][1] +
                mat_A[174][1] * mat_B[203][1] +
                mat_A[174][2] * mat_B[211][1] +
                mat_A[174][3] * mat_B[219][1] +
                mat_A[175][0] * mat_B[227][1] +
                mat_A[175][1] * mat_B[235][1] +
                mat_A[175][2] * mat_B[243][1] +
                mat_A[175][3] * mat_B[251][1];
    mat_C[171][2] <=
                mat_A[168][0] * mat_B[3][2] +
                mat_A[168][1] * mat_B[11][2] +
                mat_A[168][2] * mat_B[19][2] +
                mat_A[168][3] * mat_B[27][2] +
                mat_A[169][0] * mat_B[35][2] +
                mat_A[169][1] * mat_B[43][2] +
                mat_A[169][2] * mat_B[51][2] +
                mat_A[169][3] * mat_B[59][2] +
                mat_A[170][0] * mat_B[67][2] +
                mat_A[170][1] * mat_B[75][2] +
                mat_A[170][2] * mat_B[83][2] +
                mat_A[170][3] * mat_B[91][2] +
                mat_A[171][0] * mat_B[99][2] +
                mat_A[171][1] * mat_B[107][2] +
                mat_A[171][2] * mat_B[115][2] +
                mat_A[171][3] * mat_B[123][2] +
                mat_A[172][0] * mat_B[131][2] +
                mat_A[172][1] * mat_B[139][2] +
                mat_A[172][2] * mat_B[147][2] +
                mat_A[172][3] * mat_B[155][2] +
                mat_A[173][0] * mat_B[163][2] +
                mat_A[173][1] * mat_B[171][2] +
                mat_A[173][2] * mat_B[179][2] +
                mat_A[173][3] * mat_B[187][2] +
                mat_A[174][0] * mat_B[195][2] +
                mat_A[174][1] * mat_B[203][2] +
                mat_A[174][2] * mat_B[211][2] +
                mat_A[174][3] * mat_B[219][2] +
                mat_A[175][0] * mat_B[227][2] +
                mat_A[175][1] * mat_B[235][2] +
                mat_A[175][2] * mat_B[243][2] +
                mat_A[175][3] * mat_B[251][2];
    mat_C[171][3] <=
                mat_A[168][0] * mat_B[3][3] +
                mat_A[168][1] * mat_B[11][3] +
                mat_A[168][2] * mat_B[19][3] +
                mat_A[168][3] * mat_B[27][3] +
                mat_A[169][0] * mat_B[35][3] +
                mat_A[169][1] * mat_B[43][3] +
                mat_A[169][2] * mat_B[51][3] +
                mat_A[169][3] * mat_B[59][3] +
                mat_A[170][0] * mat_B[67][3] +
                mat_A[170][1] * mat_B[75][3] +
                mat_A[170][2] * mat_B[83][3] +
                mat_A[170][3] * mat_B[91][3] +
                mat_A[171][0] * mat_B[99][3] +
                mat_A[171][1] * mat_B[107][3] +
                mat_A[171][2] * mat_B[115][3] +
                mat_A[171][3] * mat_B[123][3] +
                mat_A[172][0] * mat_B[131][3] +
                mat_A[172][1] * mat_B[139][3] +
                mat_A[172][2] * mat_B[147][3] +
                mat_A[172][3] * mat_B[155][3] +
                mat_A[173][0] * mat_B[163][3] +
                mat_A[173][1] * mat_B[171][3] +
                mat_A[173][2] * mat_B[179][3] +
                mat_A[173][3] * mat_B[187][3] +
                mat_A[174][0] * mat_B[195][3] +
                mat_A[174][1] * mat_B[203][3] +
                mat_A[174][2] * mat_B[211][3] +
                mat_A[174][3] * mat_B[219][3] +
                mat_A[175][0] * mat_B[227][3] +
                mat_A[175][1] * mat_B[235][3] +
                mat_A[175][2] * mat_B[243][3] +
                mat_A[175][3] * mat_B[251][3];
    mat_C[172][0] <=
                mat_A[168][0] * mat_B[4][0] +
                mat_A[168][1] * mat_B[12][0] +
                mat_A[168][2] * mat_B[20][0] +
                mat_A[168][3] * mat_B[28][0] +
                mat_A[169][0] * mat_B[36][0] +
                mat_A[169][1] * mat_B[44][0] +
                mat_A[169][2] * mat_B[52][0] +
                mat_A[169][3] * mat_B[60][0] +
                mat_A[170][0] * mat_B[68][0] +
                mat_A[170][1] * mat_B[76][0] +
                mat_A[170][2] * mat_B[84][0] +
                mat_A[170][3] * mat_B[92][0] +
                mat_A[171][0] * mat_B[100][0] +
                mat_A[171][1] * mat_B[108][0] +
                mat_A[171][2] * mat_B[116][0] +
                mat_A[171][3] * mat_B[124][0] +
                mat_A[172][0] * mat_B[132][0] +
                mat_A[172][1] * mat_B[140][0] +
                mat_A[172][2] * mat_B[148][0] +
                mat_A[172][3] * mat_B[156][0] +
                mat_A[173][0] * mat_B[164][0] +
                mat_A[173][1] * mat_B[172][0] +
                mat_A[173][2] * mat_B[180][0] +
                mat_A[173][3] * mat_B[188][0] +
                mat_A[174][0] * mat_B[196][0] +
                mat_A[174][1] * mat_B[204][0] +
                mat_A[174][2] * mat_B[212][0] +
                mat_A[174][3] * mat_B[220][0] +
                mat_A[175][0] * mat_B[228][0] +
                mat_A[175][1] * mat_B[236][0] +
                mat_A[175][2] * mat_B[244][0] +
                mat_A[175][3] * mat_B[252][0];
    mat_C[172][1] <=
                mat_A[168][0] * mat_B[4][1] +
                mat_A[168][1] * mat_B[12][1] +
                mat_A[168][2] * mat_B[20][1] +
                mat_A[168][3] * mat_B[28][1] +
                mat_A[169][0] * mat_B[36][1] +
                mat_A[169][1] * mat_B[44][1] +
                mat_A[169][2] * mat_B[52][1] +
                mat_A[169][3] * mat_B[60][1] +
                mat_A[170][0] * mat_B[68][1] +
                mat_A[170][1] * mat_B[76][1] +
                mat_A[170][2] * mat_B[84][1] +
                mat_A[170][3] * mat_B[92][1] +
                mat_A[171][0] * mat_B[100][1] +
                mat_A[171][1] * mat_B[108][1] +
                mat_A[171][2] * mat_B[116][1] +
                mat_A[171][3] * mat_B[124][1] +
                mat_A[172][0] * mat_B[132][1] +
                mat_A[172][1] * mat_B[140][1] +
                mat_A[172][2] * mat_B[148][1] +
                mat_A[172][3] * mat_B[156][1] +
                mat_A[173][0] * mat_B[164][1] +
                mat_A[173][1] * mat_B[172][1] +
                mat_A[173][2] * mat_B[180][1] +
                mat_A[173][3] * mat_B[188][1] +
                mat_A[174][0] * mat_B[196][1] +
                mat_A[174][1] * mat_B[204][1] +
                mat_A[174][2] * mat_B[212][1] +
                mat_A[174][3] * mat_B[220][1] +
                mat_A[175][0] * mat_B[228][1] +
                mat_A[175][1] * mat_B[236][1] +
                mat_A[175][2] * mat_B[244][1] +
                mat_A[175][3] * mat_B[252][1];
    mat_C[172][2] <=
                mat_A[168][0] * mat_B[4][2] +
                mat_A[168][1] * mat_B[12][2] +
                mat_A[168][2] * mat_B[20][2] +
                mat_A[168][3] * mat_B[28][2] +
                mat_A[169][0] * mat_B[36][2] +
                mat_A[169][1] * mat_B[44][2] +
                mat_A[169][2] * mat_B[52][2] +
                mat_A[169][3] * mat_B[60][2] +
                mat_A[170][0] * mat_B[68][2] +
                mat_A[170][1] * mat_B[76][2] +
                mat_A[170][2] * mat_B[84][2] +
                mat_A[170][3] * mat_B[92][2] +
                mat_A[171][0] * mat_B[100][2] +
                mat_A[171][1] * mat_B[108][2] +
                mat_A[171][2] * mat_B[116][2] +
                mat_A[171][3] * mat_B[124][2] +
                mat_A[172][0] * mat_B[132][2] +
                mat_A[172][1] * mat_B[140][2] +
                mat_A[172][2] * mat_B[148][2] +
                mat_A[172][3] * mat_B[156][2] +
                mat_A[173][0] * mat_B[164][2] +
                mat_A[173][1] * mat_B[172][2] +
                mat_A[173][2] * mat_B[180][2] +
                mat_A[173][3] * mat_B[188][2] +
                mat_A[174][0] * mat_B[196][2] +
                mat_A[174][1] * mat_B[204][2] +
                mat_A[174][2] * mat_B[212][2] +
                mat_A[174][3] * mat_B[220][2] +
                mat_A[175][0] * mat_B[228][2] +
                mat_A[175][1] * mat_B[236][2] +
                mat_A[175][2] * mat_B[244][2] +
                mat_A[175][3] * mat_B[252][2];
    mat_C[172][3] <=
                mat_A[168][0] * mat_B[4][3] +
                mat_A[168][1] * mat_B[12][3] +
                mat_A[168][2] * mat_B[20][3] +
                mat_A[168][3] * mat_B[28][3] +
                mat_A[169][0] * mat_B[36][3] +
                mat_A[169][1] * mat_B[44][3] +
                mat_A[169][2] * mat_B[52][3] +
                mat_A[169][3] * mat_B[60][3] +
                mat_A[170][0] * mat_B[68][3] +
                mat_A[170][1] * mat_B[76][3] +
                mat_A[170][2] * mat_B[84][3] +
                mat_A[170][3] * mat_B[92][3] +
                mat_A[171][0] * mat_B[100][3] +
                mat_A[171][1] * mat_B[108][3] +
                mat_A[171][2] * mat_B[116][3] +
                mat_A[171][3] * mat_B[124][3] +
                mat_A[172][0] * mat_B[132][3] +
                mat_A[172][1] * mat_B[140][3] +
                mat_A[172][2] * mat_B[148][3] +
                mat_A[172][3] * mat_B[156][3] +
                mat_A[173][0] * mat_B[164][3] +
                mat_A[173][1] * mat_B[172][3] +
                mat_A[173][2] * mat_B[180][3] +
                mat_A[173][3] * mat_B[188][3] +
                mat_A[174][0] * mat_B[196][3] +
                mat_A[174][1] * mat_B[204][3] +
                mat_A[174][2] * mat_B[212][3] +
                mat_A[174][3] * mat_B[220][3] +
                mat_A[175][0] * mat_B[228][3] +
                mat_A[175][1] * mat_B[236][3] +
                mat_A[175][2] * mat_B[244][3] +
                mat_A[175][3] * mat_B[252][3];
    mat_C[173][0] <=
                mat_A[168][0] * mat_B[5][0] +
                mat_A[168][1] * mat_B[13][0] +
                mat_A[168][2] * mat_B[21][0] +
                mat_A[168][3] * mat_B[29][0] +
                mat_A[169][0] * mat_B[37][0] +
                mat_A[169][1] * mat_B[45][0] +
                mat_A[169][2] * mat_B[53][0] +
                mat_A[169][3] * mat_B[61][0] +
                mat_A[170][0] * mat_B[69][0] +
                mat_A[170][1] * mat_B[77][0] +
                mat_A[170][2] * mat_B[85][0] +
                mat_A[170][3] * mat_B[93][0] +
                mat_A[171][0] * mat_B[101][0] +
                mat_A[171][1] * mat_B[109][0] +
                mat_A[171][2] * mat_B[117][0] +
                mat_A[171][3] * mat_B[125][0] +
                mat_A[172][0] * mat_B[133][0] +
                mat_A[172][1] * mat_B[141][0] +
                mat_A[172][2] * mat_B[149][0] +
                mat_A[172][3] * mat_B[157][0] +
                mat_A[173][0] * mat_B[165][0] +
                mat_A[173][1] * mat_B[173][0] +
                mat_A[173][2] * mat_B[181][0] +
                mat_A[173][3] * mat_B[189][0] +
                mat_A[174][0] * mat_B[197][0] +
                mat_A[174][1] * mat_B[205][0] +
                mat_A[174][2] * mat_B[213][0] +
                mat_A[174][3] * mat_B[221][0] +
                mat_A[175][0] * mat_B[229][0] +
                mat_A[175][1] * mat_B[237][0] +
                mat_A[175][2] * mat_B[245][0] +
                mat_A[175][3] * mat_B[253][0];
    mat_C[173][1] <=
                mat_A[168][0] * mat_B[5][1] +
                mat_A[168][1] * mat_B[13][1] +
                mat_A[168][2] * mat_B[21][1] +
                mat_A[168][3] * mat_B[29][1] +
                mat_A[169][0] * mat_B[37][1] +
                mat_A[169][1] * mat_B[45][1] +
                mat_A[169][2] * mat_B[53][1] +
                mat_A[169][3] * mat_B[61][1] +
                mat_A[170][0] * mat_B[69][1] +
                mat_A[170][1] * mat_B[77][1] +
                mat_A[170][2] * mat_B[85][1] +
                mat_A[170][3] * mat_B[93][1] +
                mat_A[171][0] * mat_B[101][1] +
                mat_A[171][1] * mat_B[109][1] +
                mat_A[171][2] * mat_B[117][1] +
                mat_A[171][3] * mat_B[125][1] +
                mat_A[172][0] * mat_B[133][1] +
                mat_A[172][1] * mat_B[141][1] +
                mat_A[172][2] * mat_B[149][1] +
                mat_A[172][3] * mat_B[157][1] +
                mat_A[173][0] * mat_B[165][1] +
                mat_A[173][1] * mat_B[173][1] +
                mat_A[173][2] * mat_B[181][1] +
                mat_A[173][3] * mat_B[189][1] +
                mat_A[174][0] * mat_B[197][1] +
                mat_A[174][1] * mat_B[205][1] +
                mat_A[174][2] * mat_B[213][1] +
                mat_A[174][3] * mat_B[221][1] +
                mat_A[175][0] * mat_B[229][1] +
                mat_A[175][1] * mat_B[237][1] +
                mat_A[175][2] * mat_B[245][1] +
                mat_A[175][3] * mat_B[253][1];
    mat_C[173][2] <=
                mat_A[168][0] * mat_B[5][2] +
                mat_A[168][1] * mat_B[13][2] +
                mat_A[168][2] * mat_B[21][2] +
                mat_A[168][3] * mat_B[29][2] +
                mat_A[169][0] * mat_B[37][2] +
                mat_A[169][1] * mat_B[45][2] +
                mat_A[169][2] * mat_B[53][2] +
                mat_A[169][3] * mat_B[61][2] +
                mat_A[170][0] * mat_B[69][2] +
                mat_A[170][1] * mat_B[77][2] +
                mat_A[170][2] * mat_B[85][2] +
                mat_A[170][3] * mat_B[93][2] +
                mat_A[171][0] * mat_B[101][2] +
                mat_A[171][1] * mat_B[109][2] +
                mat_A[171][2] * mat_B[117][2] +
                mat_A[171][3] * mat_B[125][2] +
                mat_A[172][0] * mat_B[133][2] +
                mat_A[172][1] * mat_B[141][2] +
                mat_A[172][2] * mat_B[149][2] +
                mat_A[172][3] * mat_B[157][2] +
                mat_A[173][0] * mat_B[165][2] +
                mat_A[173][1] * mat_B[173][2] +
                mat_A[173][2] * mat_B[181][2] +
                mat_A[173][3] * mat_B[189][2] +
                mat_A[174][0] * mat_B[197][2] +
                mat_A[174][1] * mat_B[205][2] +
                mat_A[174][2] * mat_B[213][2] +
                mat_A[174][3] * mat_B[221][2] +
                mat_A[175][0] * mat_B[229][2] +
                mat_A[175][1] * mat_B[237][2] +
                mat_A[175][2] * mat_B[245][2] +
                mat_A[175][3] * mat_B[253][2];
    mat_C[173][3] <=
                mat_A[168][0] * mat_B[5][3] +
                mat_A[168][1] * mat_B[13][3] +
                mat_A[168][2] * mat_B[21][3] +
                mat_A[168][3] * mat_B[29][3] +
                mat_A[169][0] * mat_B[37][3] +
                mat_A[169][1] * mat_B[45][3] +
                mat_A[169][2] * mat_B[53][3] +
                mat_A[169][3] * mat_B[61][3] +
                mat_A[170][0] * mat_B[69][3] +
                mat_A[170][1] * mat_B[77][3] +
                mat_A[170][2] * mat_B[85][3] +
                mat_A[170][3] * mat_B[93][3] +
                mat_A[171][0] * mat_B[101][3] +
                mat_A[171][1] * mat_B[109][3] +
                mat_A[171][2] * mat_B[117][3] +
                mat_A[171][3] * mat_B[125][3] +
                mat_A[172][0] * mat_B[133][3] +
                mat_A[172][1] * mat_B[141][3] +
                mat_A[172][2] * mat_B[149][3] +
                mat_A[172][3] * mat_B[157][3] +
                mat_A[173][0] * mat_B[165][3] +
                mat_A[173][1] * mat_B[173][3] +
                mat_A[173][2] * mat_B[181][3] +
                mat_A[173][3] * mat_B[189][3] +
                mat_A[174][0] * mat_B[197][3] +
                mat_A[174][1] * mat_B[205][3] +
                mat_A[174][2] * mat_B[213][3] +
                mat_A[174][3] * mat_B[221][3] +
                mat_A[175][0] * mat_B[229][3] +
                mat_A[175][1] * mat_B[237][3] +
                mat_A[175][2] * mat_B[245][3] +
                mat_A[175][3] * mat_B[253][3];
    mat_C[174][0] <=
                mat_A[168][0] * mat_B[6][0] +
                mat_A[168][1] * mat_B[14][0] +
                mat_A[168][2] * mat_B[22][0] +
                mat_A[168][3] * mat_B[30][0] +
                mat_A[169][0] * mat_B[38][0] +
                mat_A[169][1] * mat_B[46][0] +
                mat_A[169][2] * mat_B[54][0] +
                mat_A[169][3] * mat_B[62][0] +
                mat_A[170][0] * mat_B[70][0] +
                mat_A[170][1] * mat_B[78][0] +
                mat_A[170][2] * mat_B[86][0] +
                mat_A[170][3] * mat_B[94][0] +
                mat_A[171][0] * mat_B[102][0] +
                mat_A[171][1] * mat_B[110][0] +
                mat_A[171][2] * mat_B[118][0] +
                mat_A[171][3] * mat_B[126][0] +
                mat_A[172][0] * mat_B[134][0] +
                mat_A[172][1] * mat_B[142][0] +
                mat_A[172][2] * mat_B[150][0] +
                mat_A[172][3] * mat_B[158][0] +
                mat_A[173][0] * mat_B[166][0] +
                mat_A[173][1] * mat_B[174][0] +
                mat_A[173][2] * mat_B[182][0] +
                mat_A[173][3] * mat_B[190][0] +
                mat_A[174][0] * mat_B[198][0] +
                mat_A[174][1] * mat_B[206][0] +
                mat_A[174][2] * mat_B[214][0] +
                mat_A[174][3] * mat_B[222][0] +
                mat_A[175][0] * mat_B[230][0] +
                mat_A[175][1] * mat_B[238][0] +
                mat_A[175][2] * mat_B[246][0] +
                mat_A[175][3] * mat_B[254][0];
    mat_C[174][1] <=
                mat_A[168][0] * mat_B[6][1] +
                mat_A[168][1] * mat_B[14][1] +
                mat_A[168][2] * mat_B[22][1] +
                mat_A[168][3] * mat_B[30][1] +
                mat_A[169][0] * mat_B[38][1] +
                mat_A[169][1] * mat_B[46][1] +
                mat_A[169][2] * mat_B[54][1] +
                mat_A[169][3] * mat_B[62][1] +
                mat_A[170][0] * mat_B[70][1] +
                mat_A[170][1] * mat_B[78][1] +
                mat_A[170][2] * mat_B[86][1] +
                mat_A[170][3] * mat_B[94][1] +
                mat_A[171][0] * mat_B[102][1] +
                mat_A[171][1] * mat_B[110][1] +
                mat_A[171][2] * mat_B[118][1] +
                mat_A[171][3] * mat_B[126][1] +
                mat_A[172][0] * mat_B[134][1] +
                mat_A[172][1] * mat_B[142][1] +
                mat_A[172][2] * mat_B[150][1] +
                mat_A[172][3] * mat_B[158][1] +
                mat_A[173][0] * mat_B[166][1] +
                mat_A[173][1] * mat_B[174][1] +
                mat_A[173][2] * mat_B[182][1] +
                mat_A[173][3] * mat_B[190][1] +
                mat_A[174][0] * mat_B[198][1] +
                mat_A[174][1] * mat_B[206][1] +
                mat_A[174][2] * mat_B[214][1] +
                mat_A[174][3] * mat_B[222][1] +
                mat_A[175][0] * mat_B[230][1] +
                mat_A[175][1] * mat_B[238][1] +
                mat_A[175][2] * mat_B[246][1] +
                mat_A[175][3] * mat_B[254][1];
    mat_C[174][2] <=
                mat_A[168][0] * mat_B[6][2] +
                mat_A[168][1] * mat_B[14][2] +
                mat_A[168][2] * mat_B[22][2] +
                mat_A[168][3] * mat_B[30][2] +
                mat_A[169][0] * mat_B[38][2] +
                mat_A[169][1] * mat_B[46][2] +
                mat_A[169][2] * mat_B[54][2] +
                mat_A[169][3] * mat_B[62][2] +
                mat_A[170][0] * mat_B[70][2] +
                mat_A[170][1] * mat_B[78][2] +
                mat_A[170][2] * mat_B[86][2] +
                mat_A[170][3] * mat_B[94][2] +
                mat_A[171][0] * mat_B[102][2] +
                mat_A[171][1] * mat_B[110][2] +
                mat_A[171][2] * mat_B[118][2] +
                mat_A[171][3] * mat_B[126][2] +
                mat_A[172][0] * mat_B[134][2] +
                mat_A[172][1] * mat_B[142][2] +
                mat_A[172][2] * mat_B[150][2] +
                mat_A[172][3] * mat_B[158][2] +
                mat_A[173][0] * mat_B[166][2] +
                mat_A[173][1] * mat_B[174][2] +
                mat_A[173][2] * mat_B[182][2] +
                mat_A[173][3] * mat_B[190][2] +
                mat_A[174][0] * mat_B[198][2] +
                mat_A[174][1] * mat_B[206][2] +
                mat_A[174][2] * mat_B[214][2] +
                mat_A[174][3] * mat_B[222][2] +
                mat_A[175][0] * mat_B[230][2] +
                mat_A[175][1] * mat_B[238][2] +
                mat_A[175][2] * mat_B[246][2] +
                mat_A[175][3] * mat_B[254][2];
    mat_C[174][3] <=
                mat_A[168][0] * mat_B[6][3] +
                mat_A[168][1] * mat_B[14][3] +
                mat_A[168][2] * mat_B[22][3] +
                mat_A[168][3] * mat_B[30][3] +
                mat_A[169][0] * mat_B[38][3] +
                mat_A[169][1] * mat_B[46][3] +
                mat_A[169][2] * mat_B[54][3] +
                mat_A[169][3] * mat_B[62][3] +
                mat_A[170][0] * mat_B[70][3] +
                mat_A[170][1] * mat_B[78][3] +
                mat_A[170][2] * mat_B[86][3] +
                mat_A[170][3] * mat_B[94][3] +
                mat_A[171][0] * mat_B[102][3] +
                mat_A[171][1] * mat_B[110][3] +
                mat_A[171][2] * mat_B[118][3] +
                mat_A[171][3] * mat_B[126][3] +
                mat_A[172][0] * mat_B[134][3] +
                mat_A[172][1] * mat_B[142][3] +
                mat_A[172][2] * mat_B[150][3] +
                mat_A[172][3] * mat_B[158][3] +
                mat_A[173][0] * mat_B[166][3] +
                mat_A[173][1] * mat_B[174][3] +
                mat_A[173][2] * mat_B[182][3] +
                mat_A[173][3] * mat_B[190][3] +
                mat_A[174][0] * mat_B[198][3] +
                mat_A[174][1] * mat_B[206][3] +
                mat_A[174][2] * mat_B[214][3] +
                mat_A[174][3] * mat_B[222][3] +
                mat_A[175][0] * mat_B[230][3] +
                mat_A[175][1] * mat_B[238][3] +
                mat_A[175][2] * mat_B[246][3] +
                mat_A[175][3] * mat_B[254][3];
    mat_C[175][0] <=
                mat_A[168][0] * mat_B[7][0] +
                mat_A[168][1] * mat_B[15][0] +
                mat_A[168][2] * mat_B[23][0] +
                mat_A[168][3] * mat_B[31][0] +
                mat_A[169][0] * mat_B[39][0] +
                mat_A[169][1] * mat_B[47][0] +
                mat_A[169][2] * mat_B[55][0] +
                mat_A[169][3] * mat_B[63][0] +
                mat_A[170][0] * mat_B[71][0] +
                mat_A[170][1] * mat_B[79][0] +
                mat_A[170][2] * mat_B[87][0] +
                mat_A[170][3] * mat_B[95][0] +
                mat_A[171][0] * mat_B[103][0] +
                mat_A[171][1] * mat_B[111][0] +
                mat_A[171][2] * mat_B[119][0] +
                mat_A[171][3] * mat_B[127][0] +
                mat_A[172][0] * mat_B[135][0] +
                mat_A[172][1] * mat_B[143][0] +
                mat_A[172][2] * mat_B[151][0] +
                mat_A[172][3] * mat_B[159][0] +
                mat_A[173][0] * mat_B[167][0] +
                mat_A[173][1] * mat_B[175][0] +
                mat_A[173][2] * mat_B[183][0] +
                mat_A[173][3] * mat_B[191][0] +
                mat_A[174][0] * mat_B[199][0] +
                mat_A[174][1] * mat_B[207][0] +
                mat_A[174][2] * mat_B[215][0] +
                mat_A[174][3] * mat_B[223][0] +
                mat_A[175][0] * mat_B[231][0] +
                mat_A[175][1] * mat_B[239][0] +
                mat_A[175][2] * mat_B[247][0] +
                mat_A[175][3] * mat_B[255][0];
    mat_C[175][1] <=
                mat_A[168][0] * mat_B[7][1] +
                mat_A[168][1] * mat_B[15][1] +
                mat_A[168][2] * mat_B[23][1] +
                mat_A[168][3] * mat_B[31][1] +
                mat_A[169][0] * mat_B[39][1] +
                mat_A[169][1] * mat_B[47][1] +
                mat_A[169][2] * mat_B[55][1] +
                mat_A[169][3] * mat_B[63][1] +
                mat_A[170][0] * mat_B[71][1] +
                mat_A[170][1] * mat_B[79][1] +
                mat_A[170][2] * mat_B[87][1] +
                mat_A[170][3] * mat_B[95][1] +
                mat_A[171][0] * mat_B[103][1] +
                mat_A[171][1] * mat_B[111][1] +
                mat_A[171][2] * mat_B[119][1] +
                mat_A[171][3] * mat_B[127][1] +
                mat_A[172][0] * mat_B[135][1] +
                mat_A[172][1] * mat_B[143][1] +
                mat_A[172][2] * mat_B[151][1] +
                mat_A[172][3] * mat_B[159][1] +
                mat_A[173][0] * mat_B[167][1] +
                mat_A[173][1] * mat_B[175][1] +
                mat_A[173][2] * mat_B[183][1] +
                mat_A[173][3] * mat_B[191][1] +
                mat_A[174][0] * mat_B[199][1] +
                mat_A[174][1] * mat_B[207][1] +
                mat_A[174][2] * mat_B[215][1] +
                mat_A[174][3] * mat_B[223][1] +
                mat_A[175][0] * mat_B[231][1] +
                mat_A[175][1] * mat_B[239][1] +
                mat_A[175][2] * mat_B[247][1] +
                mat_A[175][3] * mat_B[255][1];
    mat_C[175][2] <=
                mat_A[168][0] * mat_B[7][2] +
                mat_A[168][1] * mat_B[15][2] +
                mat_A[168][2] * mat_B[23][2] +
                mat_A[168][3] * mat_B[31][2] +
                mat_A[169][0] * mat_B[39][2] +
                mat_A[169][1] * mat_B[47][2] +
                mat_A[169][2] * mat_B[55][2] +
                mat_A[169][3] * mat_B[63][2] +
                mat_A[170][0] * mat_B[71][2] +
                mat_A[170][1] * mat_B[79][2] +
                mat_A[170][2] * mat_B[87][2] +
                mat_A[170][3] * mat_B[95][2] +
                mat_A[171][0] * mat_B[103][2] +
                mat_A[171][1] * mat_B[111][2] +
                mat_A[171][2] * mat_B[119][2] +
                mat_A[171][3] * mat_B[127][2] +
                mat_A[172][0] * mat_B[135][2] +
                mat_A[172][1] * mat_B[143][2] +
                mat_A[172][2] * mat_B[151][2] +
                mat_A[172][3] * mat_B[159][2] +
                mat_A[173][0] * mat_B[167][2] +
                mat_A[173][1] * mat_B[175][2] +
                mat_A[173][2] * mat_B[183][2] +
                mat_A[173][3] * mat_B[191][2] +
                mat_A[174][0] * mat_B[199][2] +
                mat_A[174][1] * mat_B[207][2] +
                mat_A[174][2] * mat_B[215][2] +
                mat_A[174][3] * mat_B[223][2] +
                mat_A[175][0] * mat_B[231][2] +
                mat_A[175][1] * mat_B[239][2] +
                mat_A[175][2] * mat_B[247][2] +
                mat_A[175][3] * mat_B[255][2];
    mat_C[175][3] <=
                mat_A[168][0] * mat_B[7][3] +
                mat_A[168][1] * mat_B[15][3] +
                mat_A[168][2] * mat_B[23][3] +
                mat_A[168][3] * mat_B[31][3] +
                mat_A[169][0] * mat_B[39][3] +
                mat_A[169][1] * mat_B[47][3] +
                mat_A[169][2] * mat_B[55][3] +
                mat_A[169][3] * mat_B[63][3] +
                mat_A[170][0] * mat_B[71][3] +
                mat_A[170][1] * mat_B[79][3] +
                mat_A[170][2] * mat_B[87][3] +
                mat_A[170][3] * mat_B[95][3] +
                mat_A[171][0] * mat_B[103][3] +
                mat_A[171][1] * mat_B[111][3] +
                mat_A[171][2] * mat_B[119][3] +
                mat_A[171][3] * mat_B[127][3] +
                mat_A[172][0] * mat_B[135][3] +
                mat_A[172][1] * mat_B[143][3] +
                mat_A[172][2] * mat_B[151][3] +
                mat_A[172][3] * mat_B[159][3] +
                mat_A[173][0] * mat_B[167][3] +
                mat_A[173][1] * mat_B[175][3] +
                mat_A[173][2] * mat_B[183][3] +
                mat_A[173][3] * mat_B[191][3] +
                mat_A[174][0] * mat_B[199][3] +
                mat_A[174][1] * mat_B[207][3] +
                mat_A[174][2] * mat_B[215][3] +
                mat_A[174][3] * mat_B[223][3] +
                mat_A[175][0] * mat_B[231][3] +
                mat_A[175][1] * mat_B[239][3] +
                mat_A[175][2] * mat_B[247][3] +
                mat_A[175][3] * mat_B[255][3];
    mat_C[176][0] <=
                mat_A[176][0] * mat_B[0][0] +
                mat_A[176][1] * mat_B[8][0] +
                mat_A[176][2] * mat_B[16][0] +
                mat_A[176][3] * mat_B[24][0] +
                mat_A[177][0] * mat_B[32][0] +
                mat_A[177][1] * mat_B[40][0] +
                mat_A[177][2] * mat_B[48][0] +
                mat_A[177][3] * mat_B[56][0] +
                mat_A[178][0] * mat_B[64][0] +
                mat_A[178][1] * mat_B[72][0] +
                mat_A[178][2] * mat_B[80][0] +
                mat_A[178][3] * mat_B[88][0] +
                mat_A[179][0] * mat_B[96][0] +
                mat_A[179][1] * mat_B[104][0] +
                mat_A[179][2] * mat_B[112][0] +
                mat_A[179][3] * mat_B[120][0] +
                mat_A[180][0] * mat_B[128][0] +
                mat_A[180][1] * mat_B[136][0] +
                mat_A[180][2] * mat_B[144][0] +
                mat_A[180][3] * mat_B[152][0] +
                mat_A[181][0] * mat_B[160][0] +
                mat_A[181][1] * mat_B[168][0] +
                mat_A[181][2] * mat_B[176][0] +
                mat_A[181][3] * mat_B[184][0] +
                mat_A[182][0] * mat_B[192][0] +
                mat_A[182][1] * mat_B[200][0] +
                mat_A[182][2] * mat_B[208][0] +
                mat_A[182][3] * mat_B[216][0] +
                mat_A[183][0] * mat_B[224][0] +
                mat_A[183][1] * mat_B[232][0] +
                mat_A[183][2] * mat_B[240][0] +
                mat_A[183][3] * mat_B[248][0];
    mat_C[176][1] <=
                mat_A[176][0] * mat_B[0][1] +
                mat_A[176][1] * mat_B[8][1] +
                mat_A[176][2] * mat_B[16][1] +
                mat_A[176][3] * mat_B[24][1] +
                mat_A[177][0] * mat_B[32][1] +
                mat_A[177][1] * mat_B[40][1] +
                mat_A[177][2] * mat_B[48][1] +
                mat_A[177][3] * mat_B[56][1] +
                mat_A[178][0] * mat_B[64][1] +
                mat_A[178][1] * mat_B[72][1] +
                mat_A[178][2] * mat_B[80][1] +
                mat_A[178][3] * mat_B[88][1] +
                mat_A[179][0] * mat_B[96][1] +
                mat_A[179][1] * mat_B[104][1] +
                mat_A[179][2] * mat_B[112][1] +
                mat_A[179][3] * mat_B[120][1] +
                mat_A[180][0] * mat_B[128][1] +
                mat_A[180][1] * mat_B[136][1] +
                mat_A[180][2] * mat_B[144][1] +
                mat_A[180][3] * mat_B[152][1] +
                mat_A[181][0] * mat_B[160][1] +
                mat_A[181][1] * mat_B[168][1] +
                mat_A[181][2] * mat_B[176][1] +
                mat_A[181][3] * mat_B[184][1] +
                mat_A[182][0] * mat_B[192][1] +
                mat_A[182][1] * mat_B[200][1] +
                mat_A[182][2] * mat_B[208][1] +
                mat_A[182][3] * mat_B[216][1] +
                mat_A[183][0] * mat_B[224][1] +
                mat_A[183][1] * mat_B[232][1] +
                mat_A[183][2] * mat_B[240][1] +
                mat_A[183][3] * mat_B[248][1];
    mat_C[176][2] <=
                mat_A[176][0] * mat_B[0][2] +
                mat_A[176][1] * mat_B[8][2] +
                mat_A[176][2] * mat_B[16][2] +
                mat_A[176][3] * mat_B[24][2] +
                mat_A[177][0] * mat_B[32][2] +
                mat_A[177][1] * mat_B[40][2] +
                mat_A[177][2] * mat_B[48][2] +
                mat_A[177][3] * mat_B[56][2] +
                mat_A[178][0] * mat_B[64][2] +
                mat_A[178][1] * mat_B[72][2] +
                mat_A[178][2] * mat_B[80][2] +
                mat_A[178][3] * mat_B[88][2] +
                mat_A[179][0] * mat_B[96][2] +
                mat_A[179][1] * mat_B[104][2] +
                mat_A[179][2] * mat_B[112][2] +
                mat_A[179][3] * mat_B[120][2] +
                mat_A[180][0] * mat_B[128][2] +
                mat_A[180][1] * mat_B[136][2] +
                mat_A[180][2] * mat_B[144][2] +
                mat_A[180][3] * mat_B[152][2] +
                mat_A[181][0] * mat_B[160][2] +
                mat_A[181][1] * mat_B[168][2] +
                mat_A[181][2] * mat_B[176][2] +
                mat_A[181][3] * mat_B[184][2] +
                mat_A[182][0] * mat_B[192][2] +
                mat_A[182][1] * mat_B[200][2] +
                mat_A[182][2] * mat_B[208][2] +
                mat_A[182][3] * mat_B[216][2] +
                mat_A[183][0] * mat_B[224][2] +
                mat_A[183][1] * mat_B[232][2] +
                mat_A[183][2] * mat_B[240][2] +
                mat_A[183][3] * mat_B[248][2];
    mat_C[176][3] <=
                mat_A[176][0] * mat_B[0][3] +
                mat_A[176][1] * mat_B[8][3] +
                mat_A[176][2] * mat_B[16][3] +
                mat_A[176][3] * mat_B[24][3] +
                mat_A[177][0] * mat_B[32][3] +
                mat_A[177][1] * mat_B[40][3] +
                mat_A[177][2] * mat_B[48][3] +
                mat_A[177][3] * mat_B[56][3] +
                mat_A[178][0] * mat_B[64][3] +
                mat_A[178][1] * mat_B[72][3] +
                mat_A[178][2] * mat_B[80][3] +
                mat_A[178][3] * mat_B[88][3] +
                mat_A[179][0] * mat_B[96][3] +
                mat_A[179][1] * mat_B[104][3] +
                mat_A[179][2] * mat_B[112][3] +
                mat_A[179][3] * mat_B[120][3] +
                mat_A[180][0] * mat_B[128][3] +
                mat_A[180][1] * mat_B[136][3] +
                mat_A[180][2] * mat_B[144][3] +
                mat_A[180][3] * mat_B[152][3] +
                mat_A[181][0] * mat_B[160][3] +
                mat_A[181][1] * mat_B[168][3] +
                mat_A[181][2] * mat_B[176][3] +
                mat_A[181][3] * mat_B[184][3] +
                mat_A[182][0] * mat_B[192][3] +
                mat_A[182][1] * mat_B[200][3] +
                mat_A[182][2] * mat_B[208][3] +
                mat_A[182][3] * mat_B[216][3] +
                mat_A[183][0] * mat_B[224][3] +
                mat_A[183][1] * mat_B[232][3] +
                mat_A[183][2] * mat_B[240][3] +
                mat_A[183][3] * mat_B[248][3];
    mat_C[177][0] <=
                mat_A[176][0] * mat_B[1][0] +
                mat_A[176][1] * mat_B[9][0] +
                mat_A[176][2] * mat_B[17][0] +
                mat_A[176][3] * mat_B[25][0] +
                mat_A[177][0] * mat_B[33][0] +
                mat_A[177][1] * mat_B[41][0] +
                mat_A[177][2] * mat_B[49][0] +
                mat_A[177][3] * mat_B[57][0] +
                mat_A[178][0] * mat_B[65][0] +
                mat_A[178][1] * mat_B[73][0] +
                mat_A[178][2] * mat_B[81][0] +
                mat_A[178][3] * mat_B[89][0] +
                mat_A[179][0] * mat_B[97][0] +
                mat_A[179][1] * mat_B[105][0] +
                mat_A[179][2] * mat_B[113][0] +
                mat_A[179][3] * mat_B[121][0] +
                mat_A[180][0] * mat_B[129][0] +
                mat_A[180][1] * mat_B[137][0] +
                mat_A[180][2] * mat_B[145][0] +
                mat_A[180][3] * mat_B[153][0] +
                mat_A[181][0] * mat_B[161][0] +
                mat_A[181][1] * mat_B[169][0] +
                mat_A[181][2] * mat_B[177][0] +
                mat_A[181][3] * mat_B[185][0] +
                mat_A[182][0] * mat_B[193][0] +
                mat_A[182][1] * mat_B[201][0] +
                mat_A[182][2] * mat_B[209][0] +
                mat_A[182][3] * mat_B[217][0] +
                mat_A[183][0] * mat_B[225][0] +
                mat_A[183][1] * mat_B[233][0] +
                mat_A[183][2] * mat_B[241][0] +
                mat_A[183][3] * mat_B[249][0];
    mat_C[177][1] <=
                mat_A[176][0] * mat_B[1][1] +
                mat_A[176][1] * mat_B[9][1] +
                mat_A[176][2] * mat_B[17][1] +
                mat_A[176][3] * mat_B[25][1] +
                mat_A[177][0] * mat_B[33][1] +
                mat_A[177][1] * mat_B[41][1] +
                mat_A[177][2] * mat_B[49][1] +
                mat_A[177][3] * mat_B[57][1] +
                mat_A[178][0] * mat_B[65][1] +
                mat_A[178][1] * mat_B[73][1] +
                mat_A[178][2] * mat_B[81][1] +
                mat_A[178][3] * mat_B[89][1] +
                mat_A[179][0] * mat_B[97][1] +
                mat_A[179][1] * mat_B[105][1] +
                mat_A[179][2] * mat_B[113][1] +
                mat_A[179][3] * mat_B[121][1] +
                mat_A[180][0] * mat_B[129][1] +
                mat_A[180][1] * mat_B[137][1] +
                mat_A[180][2] * mat_B[145][1] +
                mat_A[180][3] * mat_B[153][1] +
                mat_A[181][0] * mat_B[161][1] +
                mat_A[181][1] * mat_B[169][1] +
                mat_A[181][2] * mat_B[177][1] +
                mat_A[181][3] * mat_B[185][1] +
                mat_A[182][0] * mat_B[193][1] +
                mat_A[182][1] * mat_B[201][1] +
                mat_A[182][2] * mat_B[209][1] +
                mat_A[182][3] * mat_B[217][1] +
                mat_A[183][0] * mat_B[225][1] +
                mat_A[183][1] * mat_B[233][1] +
                mat_A[183][2] * mat_B[241][1] +
                mat_A[183][3] * mat_B[249][1];
    mat_C[177][2] <=
                mat_A[176][0] * mat_B[1][2] +
                mat_A[176][1] * mat_B[9][2] +
                mat_A[176][2] * mat_B[17][2] +
                mat_A[176][3] * mat_B[25][2] +
                mat_A[177][0] * mat_B[33][2] +
                mat_A[177][1] * mat_B[41][2] +
                mat_A[177][2] * mat_B[49][2] +
                mat_A[177][3] * mat_B[57][2] +
                mat_A[178][0] * mat_B[65][2] +
                mat_A[178][1] * mat_B[73][2] +
                mat_A[178][2] * mat_B[81][2] +
                mat_A[178][3] * mat_B[89][2] +
                mat_A[179][0] * mat_B[97][2] +
                mat_A[179][1] * mat_B[105][2] +
                mat_A[179][2] * mat_B[113][2] +
                mat_A[179][3] * mat_B[121][2] +
                mat_A[180][0] * mat_B[129][2] +
                mat_A[180][1] * mat_B[137][2] +
                mat_A[180][2] * mat_B[145][2] +
                mat_A[180][3] * mat_B[153][2] +
                mat_A[181][0] * mat_B[161][2] +
                mat_A[181][1] * mat_B[169][2] +
                mat_A[181][2] * mat_B[177][2] +
                mat_A[181][3] * mat_B[185][2] +
                mat_A[182][0] * mat_B[193][2] +
                mat_A[182][1] * mat_B[201][2] +
                mat_A[182][2] * mat_B[209][2] +
                mat_A[182][3] * mat_B[217][2] +
                mat_A[183][0] * mat_B[225][2] +
                mat_A[183][1] * mat_B[233][2] +
                mat_A[183][2] * mat_B[241][2] +
                mat_A[183][3] * mat_B[249][2];
    mat_C[177][3] <=
                mat_A[176][0] * mat_B[1][3] +
                mat_A[176][1] * mat_B[9][3] +
                mat_A[176][2] * mat_B[17][3] +
                mat_A[176][3] * mat_B[25][3] +
                mat_A[177][0] * mat_B[33][3] +
                mat_A[177][1] * mat_B[41][3] +
                mat_A[177][2] * mat_B[49][3] +
                mat_A[177][3] * mat_B[57][3] +
                mat_A[178][0] * mat_B[65][3] +
                mat_A[178][1] * mat_B[73][3] +
                mat_A[178][2] * mat_B[81][3] +
                mat_A[178][3] * mat_B[89][3] +
                mat_A[179][0] * mat_B[97][3] +
                mat_A[179][1] * mat_B[105][3] +
                mat_A[179][2] * mat_B[113][3] +
                mat_A[179][3] * mat_B[121][3] +
                mat_A[180][0] * mat_B[129][3] +
                mat_A[180][1] * mat_B[137][3] +
                mat_A[180][2] * mat_B[145][3] +
                mat_A[180][3] * mat_B[153][3] +
                mat_A[181][0] * mat_B[161][3] +
                mat_A[181][1] * mat_B[169][3] +
                mat_A[181][2] * mat_B[177][3] +
                mat_A[181][3] * mat_B[185][3] +
                mat_A[182][0] * mat_B[193][3] +
                mat_A[182][1] * mat_B[201][3] +
                mat_A[182][2] * mat_B[209][3] +
                mat_A[182][3] * mat_B[217][3] +
                mat_A[183][0] * mat_B[225][3] +
                mat_A[183][1] * mat_B[233][3] +
                mat_A[183][2] * mat_B[241][3] +
                mat_A[183][3] * mat_B[249][3];
    mat_C[178][0] <=
                mat_A[176][0] * mat_B[2][0] +
                mat_A[176][1] * mat_B[10][0] +
                mat_A[176][2] * mat_B[18][0] +
                mat_A[176][3] * mat_B[26][0] +
                mat_A[177][0] * mat_B[34][0] +
                mat_A[177][1] * mat_B[42][0] +
                mat_A[177][2] * mat_B[50][0] +
                mat_A[177][3] * mat_B[58][0] +
                mat_A[178][0] * mat_B[66][0] +
                mat_A[178][1] * mat_B[74][0] +
                mat_A[178][2] * mat_B[82][0] +
                mat_A[178][3] * mat_B[90][0] +
                mat_A[179][0] * mat_B[98][0] +
                mat_A[179][1] * mat_B[106][0] +
                mat_A[179][2] * mat_B[114][0] +
                mat_A[179][3] * mat_B[122][0] +
                mat_A[180][0] * mat_B[130][0] +
                mat_A[180][1] * mat_B[138][0] +
                mat_A[180][2] * mat_B[146][0] +
                mat_A[180][3] * mat_B[154][0] +
                mat_A[181][0] * mat_B[162][0] +
                mat_A[181][1] * mat_B[170][0] +
                mat_A[181][2] * mat_B[178][0] +
                mat_A[181][3] * mat_B[186][0] +
                mat_A[182][0] * mat_B[194][0] +
                mat_A[182][1] * mat_B[202][0] +
                mat_A[182][2] * mat_B[210][0] +
                mat_A[182][3] * mat_B[218][0] +
                mat_A[183][0] * mat_B[226][0] +
                mat_A[183][1] * mat_B[234][0] +
                mat_A[183][2] * mat_B[242][0] +
                mat_A[183][3] * mat_B[250][0];
    mat_C[178][1] <=
                mat_A[176][0] * mat_B[2][1] +
                mat_A[176][1] * mat_B[10][1] +
                mat_A[176][2] * mat_B[18][1] +
                mat_A[176][3] * mat_B[26][1] +
                mat_A[177][0] * mat_B[34][1] +
                mat_A[177][1] * mat_B[42][1] +
                mat_A[177][2] * mat_B[50][1] +
                mat_A[177][3] * mat_B[58][1] +
                mat_A[178][0] * mat_B[66][1] +
                mat_A[178][1] * mat_B[74][1] +
                mat_A[178][2] * mat_B[82][1] +
                mat_A[178][3] * mat_B[90][1] +
                mat_A[179][0] * mat_B[98][1] +
                mat_A[179][1] * mat_B[106][1] +
                mat_A[179][2] * mat_B[114][1] +
                mat_A[179][3] * mat_B[122][1] +
                mat_A[180][0] * mat_B[130][1] +
                mat_A[180][1] * mat_B[138][1] +
                mat_A[180][2] * mat_B[146][1] +
                mat_A[180][3] * mat_B[154][1] +
                mat_A[181][0] * mat_B[162][1] +
                mat_A[181][1] * mat_B[170][1] +
                mat_A[181][2] * mat_B[178][1] +
                mat_A[181][3] * mat_B[186][1] +
                mat_A[182][0] * mat_B[194][1] +
                mat_A[182][1] * mat_B[202][1] +
                mat_A[182][2] * mat_B[210][1] +
                mat_A[182][3] * mat_B[218][1] +
                mat_A[183][0] * mat_B[226][1] +
                mat_A[183][1] * mat_B[234][1] +
                mat_A[183][2] * mat_B[242][1] +
                mat_A[183][3] * mat_B[250][1];
    mat_C[178][2] <=
                mat_A[176][0] * mat_B[2][2] +
                mat_A[176][1] * mat_B[10][2] +
                mat_A[176][2] * mat_B[18][2] +
                mat_A[176][3] * mat_B[26][2] +
                mat_A[177][0] * mat_B[34][2] +
                mat_A[177][1] * mat_B[42][2] +
                mat_A[177][2] * mat_B[50][2] +
                mat_A[177][3] * mat_B[58][2] +
                mat_A[178][0] * mat_B[66][2] +
                mat_A[178][1] * mat_B[74][2] +
                mat_A[178][2] * mat_B[82][2] +
                mat_A[178][3] * mat_B[90][2] +
                mat_A[179][0] * mat_B[98][2] +
                mat_A[179][1] * mat_B[106][2] +
                mat_A[179][2] * mat_B[114][2] +
                mat_A[179][3] * mat_B[122][2] +
                mat_A[180][0] * mat_B[130][2] +
                mat_A[180][1] * mat_B[138][2] +
                mat_A[180][2] * mat_B[146][2] +
                mat_A[180][3] * mat_B[154][2] +
                mat_A[181][0] * mat_B[162][2] +
                mat_A[181][1] * mat_B[170][2] +
                mat_A[181][2] * mat_B[178][2] +
                mat_A[181][3] * mat_B[186][2] +
                mat_A[182][0] * mat_B[194][2] +
                mat_A[182][1] * mat_B[202][2] +
                mat_A[182][2] * mat_B[210][2] +
                mat_A[182][3] * mat_B[218][2] +
                mat_A[183][0] * mat_B[226][2] +
                mat_A[183][1] * mat_B[234][2] +
                mat_A[183][2] * mat_B[242][2] +
                mat_A[183][3] * mat_B[250][2];
    mat_C[178][3] <=
                mat_A[176][0] * mat_B[2][3] +
                mat_A[176][1] * mat_B[10][3] +
                mat_A[176][2] * mat_B[18][3] +
                mat_A[176][3] * mat_B[26][3] +
                mat_A[177][0] * mat_B[34][3] +
                mat_A[177][1] * mat_B[42][3] +
                mat_A[177][2] * mat_B[50][3] +
                mat_A[177][3] * mat_B[58][3] +
                mat_A[178][0] * mat_B[66][3] +
                mat_A[178][1] * mat_B[74][3] +
                mat_A[178][2] * mat_B[82][3] +
                mat_A[178][3] * mat_B[90][3] +
                mat_A[179][0] * mat_B[98][3] +
                mat_A[179][1] * mat_B[106][3] +
                mat_A[179][2] * mat_B[114][3] +
                mat_A[179][3] * mat_B[122][3] +
                mat_A[180][0] * mat_B[130][3] +
                mat_A[180][1] * mat_B[138][3] +
                mat_A[180][2] * mat_B[146][3] +
                mat_A[180][3] * mat_B[154][3] +
                mat_A[181][0] * mat_B[162][3] +
                mat_A[181][1] * mat_B[170][3] +
                mat_A[181][2] * mat_B[178][3] +
                mat_A[181][3] * mat_B[186][3] +
                mat_A[182][0] * mat_B[194][3] +
                mat_A[182][1] * mat_B[202][3] +
                mat_A[182][2] * mat_B[210][3] +
                mat_A[182][3] * mat_B[218][3] +
                mat_A[183][0] * mat_B[226][3] +
                mat_A[183][1] * mat_B[234][3] +
                mat_A[183][2] * mat_B[242][3] +
                mat_A[183][3] * mat_B[250][3];
    mat_C[179][0] <=
                mat_A[176][0] * mat_B[3][0] +
                mat_A[176][1] * mat_B[11][0] +
                mat_A[176][2] * mat_B[19][0] +
                mat_A[176][3] * mat_B[27][0] +
                mat_A[177][0] * mat_B[35][0] +
                mat_A[177][1] * mat_B[43][0] +
                mat_A[177][2] * mat_B[51][0] +
                mat_A[177][3] * mat_B[59][0] +
                mat_A[178][0] * mat_B[67][0] +
                mat_A[178][1] * mat_B[75][0] +
                mat_A[178][2] * mat_B[83][0] +
                mat_A[178][3] * mat_B[91][0] +
                mat_A[179][0] * mat_B[99][0] +
                mat_A[179][1] * mat_B[107][0] +
                mat_A[179][2] * mat_B[115][0] +
                mat_A[179][3] * mat_B[123][0] +
                mat_A[180][0] * mat_B[131][0] +
                mat_A[180][1] * mat_B[139][0] +
                mat_A[180][2] * mat_B[147][0] +
                mat_A[180][3] * mat_B[155][0] +
                mat_A[181][0] * mat_B[163][0] +
                mat_A[181][1] * mat_B[171][0] +
                mat_A[181][2] * mat_B[179][0] +
                mat_A[181][3] * mat_B[187][0] +
                mat_A[182][0] * mat_B[195][0] +
                mat_A[182][1] * mat_B[203][0] +
                mat_A[182][2] * mat_B[211][0] +
                mat_A[182][3] * mat_B[219][0] +
                mat_A[183][0] * mat_B[227][0] +
                mat_A[183][1] * mat_B[235][0] +
                mat_A[183][2] * mat_B[243][0] +
                mat_A[183][3] * mat_B[251][0];
    mat_C[179][1] <=
                mat_A[176][0] * mat_B[3][1] +
                mat_A[176][1] * mat_B[11][1] +
                mat_A[176][2] * mat_B[19][1] +
                mat_A[176][3] * mat_B[27][1] +
                mat_A[177][0] * mat_B[35][1] +
                mat_A[177][1] * mat_B[43][1] +
                mat_A[177][2] * mat_B[51][1] +
                mat_A[177][3] * mat_B[59][1] +
                mat_A[178][0] * mat_B[67][1] +
                mat_A[178][1] * mat_B[75][1] +
                mat_A[178][2] * mat_B[83][1] +
                mat_A[178][3] * mat_B[91][1] +
                mat_A[179][0] * mat_B[99][1] +
                mat_A[179][1] * mat_B[107][1] +
                mat_A[179][2] * mat_B[115][1] +
                mat_A[179][3] * mat_B[123][1] +
                mat_A[180][0] * mat_B[131][1] +
                mat_A[180][1] * mat_B[139][1] +
                mat_A[180][2] * mat_B[147][1] +
                mat_A[180][3] * mat_B[155][1] +
                mat_A[181][0] * mat_B[163][1] +
                mat_A[181][1] * mat_B[171][1] +
                mat_A[181][2] * mat_B[179][1] +
                mat_A[181][3] * mat_B[187][1] +
                mat_A[182][0] * mat_B[195][1] +
                mat_A[182][1] * mat_B[203][1] +
                mat_A[182][2] * mat_B[211][1] +
                mat_A[182][3] * mat_B[219][1] +
                mat_A[183][0] * mat_B[227][1] +
                mat_A[183][1] * mat_B[235][1] +
                mat_A[183][2] * mat_B[243][1] +
                mat_A[183][3] * mat_B[251][1];
    mat_C[179][2] <=
                mat_A[176][0] * mat_B[3][2] +
                mat_A[176][1] * mat_B[11][2] +
                mat_A[176][2] * mat_B[19][2] +
                mat_A[176][3] * mat_B[27][2] +
                mat_A[177][0] * mat_B[35][2] +
                mat_A[177][1] * mat_B[43][2] +
                mat_A[177][2] * mat_B[51][2] +
                mat_A[177][3] * mat_B[59][2] +
                mat_A[178][0] * mat_B[67][2] +
                mat_A[178][1] * mat_B[75][2] +
                mat_A[178][2] * mat_B[83][2] +
                mat_A[178][3] * mat_B[91][2] +
                mat_A[179][0] * mat_B[99][2] +
                mat_A[179][1] * mat_B[107][2] +
                mat_A[179][2] * mat_B[115][2] +
                mat_A[179][3] * mat_B[123][2] +
                mat_A[180][0] * mat_B[131][2] +
                mat_A[180][1] * mat_B[139][2] +
                mat_A[180][2] * mat_B[147][2] +
                mat_A[180][3] * mat_B[155][2] +
                mat_A[181][0] * mat_B[163][2] +
                mat_A[181][1] * mat_B[171][2] +
                mat_A[181][2] * mat_B[179][2] +
                mat_A[181][3] * mat_B[187][2] +
                mat_A[182][0] * mat_B[195][2] +
                mat_A[182][1] * mat_B[203][2] +
                mat_A[182][2] * mat_B[211][2] +
                mat_A[182][3] * mat_B[219][2] +
                mat_A[183][0] * mat_B[227][2] +
                mat_A[183][1] * mat_B[235][2] +
                mat_A[183][2] * mat_B[243][2] +
                mat_A[183][3] * mat_B[251][2];
    mat_C[179][3] <=
                mat_A[176][0] * mat_B[3][3] +
                mat_A[176][1] * mat_B[11][3] +
                mat_A[176][2] * mat_B[19][3] +
                mat_A[176][3] * mat_B[27][3] +
                mat_A[177][0] * mat_B[35][3] +
                mat_A[177][1] * mat_B[43][3] +
                mat_A[177][2] * mat_B[51][3] +
                mat_A[177][3] * mat_B[59][3] +
                mat_A[178][0] * mat_B[67][3] +
                mat_A[178][1] * mat_B[75][3] +
                mat_A[178][2] * mat_B[83][3] +
                mat_A[178][3] * mat_B[91][3] +
                mat_A[179][0] * mat_B[99][3] +
                mat_A[179][1] * mat_B[107][3] +
                mat_A[179][2] * mat_B[115][3] +
                mat_A[179][3] * mat_B[123][3] +
                mat_A[180][0] * mat_B[131][3] +
                mat_A[180][1] * mat_B[139][3] +
                mat_A[180][2] * mat_B[147][3] +
                mat_A[180][3] * mat_B[155][3] +
                mat_A[181][0] * mat_B[163][3] +
                mat_A[181][1] * mat_B[171][3] +
                mat_A[181][2] * mat_B[179][3] +
                mat_A[181][3] * mat_B[187][3] +
                mat_A[182][0] * mat_B[195][3] +
                mat_A[182][1] * mat_B[203][3] +
                mat_A[182][2] * mat_B[211][3] +
                mat_A[182][3] * mat_B[219][3] +
                mat_A[183][0] * mat_B[227][3] +
                mat_A[183][1] * mat_B[235][3] +
                mat_A[183][2] * mat_B[243][3] +
                mat_A[183][3] * mat_B[251][3];
    mat_C[180][0] <=
                mat_A[176][0] * mat_B[4][0] +
                mat_A[176][1] * mat_B[12][0] +
                mat_A[176][2] * mat_B[20][0] +
                mat_A[176][3] * mat_B[28][0] +
                mat_A[177][0] * mat_B[36][0] +
                mat_A[177][1] * mat_B[44][0] +
                mat_A[177][2] * mat_B[52][0] +
                mat_A[177][3] * mat_B[60][0] +
                mat_A[178][0] * mat_B[68][0] +
                mat_A[178][1] * mat_B[76][0] +
                mat_A[178][2] * mat_B[84][0] +
                mat_A[178][3] * mat_B[92][0] +
                mat_A[179][0] * mat_B[100][0] +
                mat_A[179][1] * mat_B[108][0] +
                mat_A[179][2] * mat_B[116][0] +
                mat_A[179][3] * mat_B[124][0] +
                mat_A[180][0] * mat_B[132][0] +
                mat_A[180][1] * mat_B[140][0] +
                mat_A[180][2] * mat_B[148][0] +
                mat_A[180][3] * mat_B[156][0] +
                mat_A[181][0] * mat_B[164][0] +
                mat_A[181][1] * mat_B[172][0] +
                mat_A[181][2] * mat_B[180][0] +
                mat_A[181][3] * mat_B[188][0] +
                mat_A[182][0] * mat_B[196][0] +
                mat_A[182][1] * mat_B[204][0] +
                mat_A[182][2] * mat_B[212][0] +
                mat_A[182][3] * mat_B[220][0] +
                mat_A[183][0] * mat_B[228][0] +
                mat_A[183][1] * mat_B[236][0] +
                mat_A[183][2] * mat_B[244][0] +
                mat_A[183][3] * mat_B[252][0];
    mat_C[180][1] <=
                mat_A[176][0] * mat_B[4][1] +
                mat_A[176][1] * mat_B[12][1] +
                mat_A[176][2] * mat_B[20][1] +
                mat_A[176][3] * mat_B[28][1] +
                mat_A[177][0] * mat_B[36][1] +
                mat_A[177][1] * mat_B[44][1] +
                mat_A[177][2] * mat_B[52][1] +
                mat_A[177][3] * mat_B[60][1] +
                mat_A[178][0] * mat_B[68][1] +
                mat_A[178][1] * mat_B[76][1] +
                mat_A[178][2] * mat_B[84][1] +
                mat_A[178][3] * mat_B[92][1] +
                mat_A[179][0] * mat_B[100][1] +
                mat_A[179][1] * mat_B[108][1] +
                mat_A[179][2] * mat_B[116][1] +
                mat_A[179][3] * mat_B[124][1] +
                mat_A[180][0] * mat_B[132][1] +
                mat_A[180][1] * mat_B[140][1] +
                mat_A[180][2] * mat_B[148][1] +
                mat_A[180][3] * mat_B[156][1] +
                mat_A[181][0] * mat_B[164][1] +
                mat_A[181][1] * mat_B[172][1] +
                mat_A[181][2] * mat_B[180][1] +
                mat_A[181][3] * mat_B[188][1] +
                mat_A[182][0] * mat_B[196][1] +
                mat_A[182][1] * mat_B[204][1] +
                mat_A[182][2] * mat_B[212][1] +
                mat_A[182][3] * mat_B[220][1] +
                mat_A[183][0] * mat_B[228][1] +
                mat_A[183][1] * mat_B[236][1] +
                mat_A[183][2] * mat_B[244][1] +
                mat_A[183][3] * mat_B[252][1];
    mat_C[180][2] <=
                mat_A[176][0] * mat_B[4][2] +
                mat_A[176][1] * mat_B[12][2] +
                mat_A[176][2] * mat_B[20][2] +
                mat_A[176][3] * mat_B[28][2] +
                mat_A[177][0] * mat_B[36][2] +
                mat_A[177][1] * mat_B[44][2] +
                mat_A[177][2] * mat_B[52][2] +
                mat_A[177][3] * mat_B[60][2] +
                mat_A[178][0] * mat_B[68][2] +
                mat_A[178][1] * mat_B[76][2] +
                mat_A[178][2] * mat_B[84][2] +
                mat_A[178][3] * mat_B[92][2] +
                mat_A[179][0] * mat_B[100][2] +
                mat_A[179][1] * mat_B[108][2] +
                mat_A[179][2] * mat_B[116][2] +
                mat_A[179][3] * mat_B[124][2] +
                mat_A[180][0] * mat_B[132][2] +
                mat_A[180][1] * mat_B[140][2] +
                mat_A[180][2] * mat_B[148][2] +
                mat_A[180][3] * mat_B[156][2] +
                mat_A[181][0] * mat_B[164][2] +
                mat_A[181][1] * mat_B[172][2] +
                mat_A[181][2] * mat_B[180][2] +
                mat_A[181][3] * mat_B[188][2] +
                mat_A[182][0] * mat_B[196][2] +
                mat_A[182][1] * mat_B[204][2] +
                mat_A[182][2] * mat_B[212][2] +
                mat_A[182][3] * mat_B[220][2] +
                mat_A[183][0] * mat_B[228][2] +
                mat_A[183][1] * mat_B[236][2] +
                mat_A[183][2] * mat_B[244][2] +
                mat_A[183][3] * mat_B[252][2];
    mat_C[180][3] <=
                mat_A[176][0] * mat_B[4][3] +
                mat_A[176][1] * mat_B[12][3] +
                mat_A[176][2] * mat_B[20][3] +
                mat_A[176][3] * mat_B[28][3] +
                mat_A[177][0] * mat_B[36][3] +
                mat_A[177][1] * mat_B[44][3] +
                mat_A[177][2] * mat_B[52][3] +
                mat_A[177][3] * mat_B[60][3] +
                mat_A[178][0] * mat_B[68][3] +
                mat_A[178][1] * mat_B[76][3] +
                mat_A[178][2] * mat_B[84][3] +
                mat_A[178][3] * mat_B[92][3] +
                mat_A[179][0] * mat_B[100][3] +
                mat_A[179][1] * mat_B[108][3] +
                mat_A[179][2] * mat_B[116][3] +
                mat_A[179][3] * mat_B[124][3] +
                mat_A[180][0] * mat_B[132][3] +
                mat_A[180][1] * mat_B[140][3] +
                mat_A[180][2] * mat_B[148][3] +
                mat_A[180][3] * mat_B[156][3] +
                mat_A[181][0] * mat_B[164][3] +
                mat_A[181][1] * mat_B[172][3] +
                mat_A[181][2] * mat_B[180][3] +
                mat_A[181][3] * mat_B[188][3] +
                mat_A[182][0] * mat_B[196][3] +
                mat_A[182][1] * mat_B[204][3] +
                mat_A[182][2] * mat_B[212][3] +
                mat_A[182][3] * mat_B[220][3] +
                mat_A[183][0] * mat_B[228][3] +
                mat_A[183][1] * mat_B[236][3] +
                mat_A[183][2] * mat_B[244][3] +
                mat_A[183][3] * mat_B[252][3];
    mat_C[181][0] <=
                mat_A[176][0] * mat_B[5][0] +
                mat_A[176][1] * mat_B[13][0] +
                mat_A[176][2] * mat_B[21][0] +
                mat_A[176][3] * mat_B[29][0] +
                mat_A[177][0] * mat_B[37][0] +
                mat_A[177][1] * mat_B[45][0] +
                mat_A[177][2] * mat_B[53][0] +
                mat_A[177][3] * mat_B[61][0] +
                mat_A[178][0] * mat_B[69][0] +
                mat_A[178][1] * mat_B[77][0] +
                mat_A[178][2] * mat_B[85][0] +
                mat_A[178][3] * mat_B[93][0] +
                mat_A[179][0] * mat_B[101][0] +
                mat_A[179][1] * mat_B[109][0] +
                mat_A[179][2] * mat_B[117][0] +
                mat_A[179][3] * mat_B[125][0] +
                mat_A[180][0] * mat_B[133][0] +
                mat_A[180][1] * mat_B[141][0] +
                mat_A[180][2] * mat_B[149][0] +
                mat_A[180][3] * mat_B[157][0] +
                mat_A[181][0] * mat_B[165][0] +
                mat_A[181][1] * mat_B[173][0] +
                mat_A[181][2] * mat_B[181][0] +
                mat_A[181][3] * mat_B[189][0] +
                mat_A[182][0] * mat_B[197][0] +
                mat_A[182][1] * mat_B[205][0] +
                mat_A[182][2] * mat_B[213][0] +
                mat_A[182][3] * mat_B[221][0] +
                mat_A[183][0] * mat_B[229][0] +
                mat_A[183][1] * mat_B[237][0] +
                mat_A[183][2] * mat_B[245][0] +
                mat_A[183][3] * mat_B[253][0];
    mat_C[181][1] <=
                mat_A[176][0] * mat_B[5][1] +
                mat_A[176][1] * mat_B[13][1] +
                mat_A[176][2] * mat_B[21][1] +
                mat_A[176][3] * mat_B[29][1] +
                mat_A[177][0] * mat_B[37][1] +
                mat_A[177][1] * mat_B[45][1] +
                mat_A[177][2] * mat_B[53][1] +
                mat_A[177][3] * mat_B[61][1] +
                mat_A[178][0] * mat_B[69][1] +
                mat_A[178][1] * mat_B[77][1] +
                mat_A[178][2] * mat_B[85][1] +
                mat_A[178][3] * mat_B[93][1] +
                mat_A[179][0] * mat_B[101][1] +
                mat_A[179][1] * mat_B[109][1] +
                mat_A[179][2] * mat_B[117][1] +
                mat_A[179][3] * mat_B[125][1] +
                mat_A[180][0] * mat_B[133][1] +
                mat_A[180][1] * mat_B[141][1] +
                mat_A[180][2] * mat_B[149][1] +
                mat_A[180][3] * mat_B[157][1] +
                mat_A[181][0] * mat_B[165][1] +
                mat_A[181][1] * mat_B[173][1] +
                mat_A[181][2] * mat_B[181][1] +
                mat_A[181][3] * mat_B[189][1] +
                mat_A[182][0] * mat_B[197][1] +
                mat_A[182][1] * mat_B[205][1] +
                mat_A[182][2] * mat_B[213][1] +
                mat_A[182][3] * mat_B[221][1] +
                mat_A[183][0] * mat_B[229][1] +
                mat_A[183][1] * mat_B[237][1] +
                mat_A[183][2] * mat_B[245][1] +
                mat_A[183][3] * mat_B[253][1];
    mat_C[181][2] <=
                mat_A[176][0] * mat_B[5][2] +
                mat_A[176][1] * mat_B[13][2] +
                mat_A[176][2] * mat_B[21][2] +
                mat_A[176][3] * mat_B[29][2] +
                mat_A[177][0] * mat_B[37][2] +
                mat_A[177][1] * mat_B[45][2] +
                mat_A[177][2] * mat_B[53][2] +
                mat_A[177][3] * mat_B[61][2] +
                mat_A[178][0] * mat_B[69][2] +
                mat_A[178][1] * mat_B[77][2] +
                mat_A[178][2] * mat_B[85][2] +
                mat_A[178][3] * mat_B[93][2] +
                mat_A[179][0] * mat_B[101][2] +
                mat_A[179][1] * mat_B[109][2] +
                mat_A[179][2] * mat_B[117][2] +
                mat_A[179][3] * mat_B[125][2] +
                mat_A[180][0] * mat_B[133][2] +
                mat_A[180][1] * mat_B[141][2] +
                mat_A[180][2] * mat_B[149][2] +
                mat_A[180][3] * mat_B[157][2] +
                mat_A[181][0] * mat_B[165][2] +
                mat_A[181][1] * mat_B[173][2] +
                mat_A[181][2] * mat_B[181][2] +
                mat_A[181][3] * mat_B[189][2] +
                mat_A[182][0] * mat_B[197][2] +
                mat_A[182][1] * mat_B[205][2] +
                mat_A[182][2] * mat_B[213][2] +
                mat_A[182][3] * mat_B[221][2] +
                mat_A[183][0] * mat_B[229][2] +
                mat_A[183][1] * mat_B[237][2] +
                mat_A[183][2] * mat_B[245][2] +
                mat_A[183][3] * mat_B[253][2];
    mat_C[181][3] <=
                mat_A[176][0] * mat_B[5][3] +
                mat_A[176][1] * mat_B[13][3] +
                mat_A[176][2] * mat_B[21][3] +
                mat_A[176][3] * mat_B[29][3] +
                mat_A[177][0] * mat_B[37][3] +
                mat_A[177][1] * mat_B[45][3] +
                mat_A[177][2] * mat_B[53][3] +
                mat_A[177][3] * mat_B[61][3] +
                mat_A[178][0] * mat_B[69][3] +
                mat_A[178][1] * mat_B[77][3] +
                mat_A[178][2] * mat_B[85][3] +
                mat_A[178][3] * mat_B[93][3] +
                mat_A[179][0] * mat_B[101][3] +
                mat_A[179][1] * mat_B[109][3] +
                mat_A[179][2] * mat_B[117][3] +
                mat_A[179][3] * mat_B[125][3] +
                mat_A[180][0] * mat_B[133][3] +
                mat_A[180][1] * mat_B[141][3] +
                mat_A[180][2] * mat_B[149][3] +
                mat_A[180][3] * mat_B[157][3] +
                mat_A[181][0] * mat_B[165][3] +
                mat_A[181][1] * mat_B[173][3] +
                mat_A[181][2] * mat_B[181][3] +
                mat_A[181][3] * mat_B[189][3] +
                mat_A[182][0] * mat_B[197][3] +
                mat_A[182][1] * mat_B[205][3] +
                mat_A[182][2] * mat_B[213][3] +
                mat_A[182][3] * mat_B[221][3] +
                mat_A[183][0] * mat_B[229][3] +
                mat_A[183][1] * mat_B[237][3] +
                mat_A[183][2] * mat_B[245][3] +
                mat_A[183][3] * mat_B[253][3];
    mat_C[182][0] <=
                mat_A[176][0] * mat_B[6][0] +
                mat_A[176][1] * mat_B[14][0] +
                mat_A[176][2] * mat_B[22][0] +
                mat_A[176][3] * mat_B[30][0] +
                mat_A[177][0] * mat_B[38][0] +
                mat_A[177][1] * mat_B[46][0] +
                mat_A[177][2] * mat_B[54][0] +
                mat_A[177][3] * mat_B[62][0] +
                mat_A[178][0] * mat_B[70][0] +
                mat_A[178][1] * mat_B[78][0] +
                mat_A[178][2] * mat_B[86][0] +
                mat_A[178][3] * mat_B[94][0] +
                mat_A[179][0] * mat_B[102][0] +
                mat_A[179][1] * mat_B[110][0] +
                mat_A[179][2] * mat_B[118][0] +
                mat_A[179][3] * mat_B[126][0] +
                mat_A[180][0] * mat_B[134][0] +
                mat_A[180][1] * mat_B[142][0] +
                mat_A[180][2] * mat_B[150][0] +
                mat_A[180][3] * mat_B[158][0] +
                mat_A[181][0] * mat_B[166][0] +
                mat_A[181][1] * mat_B[174][0] +
                mat_A[181][2] * mat_B[182][0] +
                mat_A[181][3] * mat_B[190][0] +
                mat_A[182][0] * mat_B[198][0] +
                mat_A[182][1] * mat_B[206][0] +
                mat_A[182][2] * mat_B[214][0] +
                mat_A[182][3] * mat_B[222][0] +
                mat_A[183][0] * mat_B[230][0] +
                mat_A[183][1] * mat_B[238][0] +
                mat_A[183][2] * mat_B[246][0] +
                mat_A[183][3] * mat_B[254][0];
    mat_C[182][1] <=
                mat_A[176][0] * mat_B[6][1] +
                mat_A[176][1] * mat_B[14][1] +
                mat_A[176][2] * mat_B[22][1] +
                mat_A[176][3] * mat_B[30][1] +
                mat_A[177][0] * mat_B[38][1] +
                mat_A[177][1] * mat_B[46][1] +
                mat_A[177][2] * mat_B[54][1] +
                mat_A[177][3] * mat_B[62][1] +
                mat_A[178][0] * mat_B[70][1] +
                mat_A[178][1] * mat_B[78][1] +
                mat_A[178][2] * mat_B[86][1] +
                mat_A[178][3] * mat_B[94][1] +
                mat_A[179][0] * mat_B[102][1] +
                mat_A[179][1] * mat_B[110][1] +
                mat_A[179][2] * mat_B[118][1] +
                mat_A[179][3] * mat_B[126][1] +
                mat_A[180][0] * mat_B[134][1] +
                mat_A[180][1] * mat_B[142][1] +
                mat_A[180][2] * mat_B[150][1] +
                mat_A[180][3] * mat_B[158][1] +
                mat_A[181][0] * mat_B[166][1] +
                mat_A[181][1] * mat_B[174][1] +
                mat_A[181][2] * mat_B[182][1] +
                mat_A[181][3] * mat_B[190][1] +
                mat_A[182][0] * mat_B[198][1] +
                mat_A[182][1] * mat_B[206][1] +
                mat_A[182][2] * mat_B[214][1] +
                mat_A[182][3] * mat_B[222][1] +
                mat_A[183][0] * mat_B[230][1] +
                mat_A[183][1] * mat_B[238][1] +
                mat_A[183][2] * mat_B[246][1] +
                mat_A[183][3] * mat_B[254][1];
    mat_C[182][2] <=
                mat_A[176][0] * mat_B[6][2] +
                mat_A[176][1] * mat_B[14][2] +
                mat_A[176][2] * mat_B[22][2] +
                mat_A[176][3] * mat_B[30][2] +
                mat_A[177][0] * mat_B[38][2] +
                mat_A[177][1] * mat_B[46][2] +
                mat_A[177][2] * mat_B[54][2] +
                mat_A[177][3] * mat_B[62][2] +
                mat_A[178][0] * mat_B[70][2] +
                mat_A[178][1] * mat_B[78][2] +
                mat_A[178][2] * mat_B[86][2] +
                mat_A[178][3] * mat_B[94][2] +
                mat_A[179][0] * mat_B[102][2] +
                mat_A[179][1] * mat_B[110][2] +
                mat_A[179][2] * mat_B[118][2] +
                mat_A[179][3] * mat_B[126][2] +
                mat_A[180][0] * mat_B[134][2] +
                mat_A[180][1] * mat_B[142][2] +
                mat_A[180][2] * mat_B[150][2] +
                mat_A[180][3] * mat_B[158][2] +
                mat_A[181][0] * mat_B[166][2] +
                mat_A[181][1] * mat_B[174][2] +
                mat_A[181][2] * mat_B[182][2] +
                mat_A[181][3] * mat_B[190][2] +
                mat_A[182][0] * mat_B[198][2] +
                mat_A[182][1] * mat_B[206][2] +
                mat_A[182][2] * mat_B[214][2] +
                mat_A[182][3] * mat_B[222][2] +
                mat_A[183][0] * mat_B[230][2] +
                mat_A[183][1] * mat_B[238][2] +
                mat_A[183][2] * mat_B[246][2] +
                mat_A[183][3] * mat_B[254][2];
    mat_C[182][3] <=
                mat_A[176][0] * mat_B[6][3] +
                mat_A[176][1] * mat_B[14][3] +
                mat_A[176][2] * mat_B[22][3] +
                mat_A[176][3] * mat_B[30][3] +
                mat_A[177][0] * mat_B[38][3] +
                mat_A[177][1] * mat_B[46][3] +
                mat_A[177][2] * mat_B[54][3] +
                mat_A[177][3] * mat_B[62][3] +
                mat_A[178][0] * mat_B[70][3] +
                mat_A[178][1] * mat_B[78][3] +
                mat_A[178][2] * mat_B[86][3] +
                mat_A[178][3] * mat_B[94][3] +
                mat_A[179][0] * mat_B[102][3] +
                mat_A[179][1] * mat_B[110][3] +
                mat_A[179][2] * mat_B[118][3] +
                mat_A[179][3] * mat_B[126][3] +
                mat_A[180][0] * mat_B[134][3] +
                mat_A[180][1] * mat_B[142][3] +
                mat_A[180][2] * mat_B[150][3] +
                mat_A[180][3] * mat_B[158][3] +
                mat_A[181][0] * mat_B[166][3] +
                mat_A[181][1] * mat_B[174][3] +
                mat_A[181][2] * mat_B[182][3] +
                mat_A[181][3] * mat_B[190][3] +
                mat_A[182][0] * mat_B[198][3] +
                mat_A[182][1] * mat_B[206][3] +
                mat_A[182][2] * mat_B[214][3] +
                mat_A[182][3] * mat_B[222][3] +
                mat_A[183][0] * mat_B[230][3] +
                mat_A[183][1] * mat_B[238][3] +
                mat_A[183][2] * mat_B[246][3] +
                mat_A[183][3] * mat_B[254][3];
    mat_C[183][0] <=
                mat_A[176][0] * mat_B[7][0] +
                mat_A[176][1] * mat_B[15][0] +
                mat_A[176][2] * mat_B[23][0] +
                mat_A[176][3] * mat_B[31][0] +
                mat_A[177][0] * mat_B[39][0] +
                mat_A[177][1] * mat_B[47][0] +
                mat_A[177][2] * mat_B[55][0] +
                mat_A[177][3] * mat_B[63][0] +
                mat_A[178][0] * mat_B[71][0] +
                mat_A[178][1] * mat_B[79][0] +
                mat_A[178][2] * mat_B[87][0] +
                mat_A[178][3] * mat_B[95][0] +
                mat_A[179][0] * mat_B[103][0] +
                mat_A[179][1] * mat_B[111][0] +
                mat_A[179][2] * mat_B[119][0] +
                mat_A[179][3] * mat_B[127][0] +
                mat_A[180][0] * mat_B[135][0] +
                mat_A[180][1] * mat_B[143][0] +
                mat_A[180][2] * mat_B[151][0] +
                mat_A[180][3] * mat_B[159][0] +
                mat_A[181][0] * mat_B[167][0] +
                mat_A[181][1] * mat_B[175][0] +
                mat_A[181][2] * mat_B[183][0] +
                mat_A[181][3] * mat_B[191][0] +
                mat_A[182][0] * mat_B[199][0] +
                mat_A[182][1] * mat_B[207][0] +
                mat_A[182][2] * mat_B[215][0] +
                mat_A[182][3] * mat_B[223][0] +
                mat_A[183][0] * mat_B[231][0] +
                mat_A[183][1] * mat_B[239][0] +
                mat_A[183][2] * mat_B[247][0] +
                mat_A[183][3] * mat_B[255][0];
    mat_C[183][1] <=
                mat_A[176][0] * mat_B[7][1] +
                mat_A[176][1] * mat_B[15][1] +
                mat_A[176][2] * mat_B[23][1] +
                mat_A[176][3] * mat_B[31][1] +
                mat_A[177][0] * mat_B[39][1] +
                mat_A[177][1] * mat_B[47][1] +
                mat_A[177][2] * mat_B[55][1] +
                mat_A[177][3] * mat_B[63][1] +
                mat_A[178][0] * mat_B[71][1] +
                mat_A[178][1] * mat_B[79][1] +
                mat_A[178][2] * mat_B[87][1] +
                mat_A[178][3] * mat_B[95][1] +
                mat_A[179][0] * mat_B[103][1] +
                mat_A[179][1] * mat_B[111][1] +
                mat_A[179][2] * mat_B[119][1] +
                mat_A[179][3] * mat_B[127][1] +
                mat_A[180][0] * mat_B[135][1] +
                mat_A[180][1] * mat_B[143][1] +
                mat_A[180][2] * mat_B[151][1] +
                mat_A[180][3] * mat_B[159][1] +
                mat_A[181][0] * mat_B[167][1] +
                mat_A[181][1] * mat_B[175][1] +
                mat_A[181][2] * mat_B[183][1] +
                mat_A[181][3] * mat_B[191][1] +
                mat_A[182][0] * mat_B[199][1] +
                mat_A[182][1] * mat_B[207][1] +
                mat_A[182][2] * mat_B[215][1] +
                mat_A[182][3] * mat_B[223][1] +
                mat_A[183][0] * mat_B[231][1] +
                mat_A[183][1] * mat_B[239][1] +
                mat_A[183][2] * mat_B[247][1] +
                mat_A[183][3] * mat_B[255][1];
    mat_C[183][2] <=
                mat_A[176][0] * mat_B[7][2] +
                mat_A[176][1] * mat_B[15][2] +
                mat_A[176][2] * mat_B[23][2] +
                mat_A[176][3] * mat_B[31][2] +
                mat_A[177][0] * mat_B[39][2] +
                mat_A[177][1] * mat_B[47][2] +
                mat_A[177][2] * mat_B[55][2] +
                mat_A[177][3] * mat_B[63][2] +
                mat_A[178][0] * mat_B[71][2] +
                mat_A[178][1] * mat_B[79][2] +
                mat_A[178][2] * mat_B[87][2] +
                mat_A[178][3] * mat_B[95][2] +
                mat_A[179][0] * mat_B[103][2] +
                mat_A[179][1] * mat_B[111][2] +
                mat_A[179][2] * mat_B[119][2] +
                mat_A[179][3] * mat_B[127][2] +
                mat_A[180][0] * mat_B[135][2] +
                mat_A[180][1] * mat_B[143][2] +
                mat_A[180][2] * mat_B[151][2] +
                mat_A[180][3] * mat_B[159][2] +
                mat_A[181][0] * mat_B[167][2] +
                mat_A[181][1] * mat_B[175][2] +
                mat_A[181][2] * mat_B[183][2] +
                mat_A[181][3] * mat_B[191][2] +
                mat_A[182][0] * mat_B[199][2] +
                mat_A[182][1] * mat_B[207][2] +
                mat_A[182][2] * mat_B[215][2] +
                mat_A[182][3] * mat_B[223][2] +
                mat_A[183][0] * mat_B[231][2] +
                mat_A[183][1] * mat_B[239][2] +
                mat_A[183][2] * mat_B[247][2] +
                mat_A[183][3] * mat_B[255][2];
    mat_C[183][3] <=
                mat_A[176][0] * mat_B[7][3] +
                mat_A[176][1] * mat_B[15][3] +
                mat_A[176][2] * mat_B[23][3] +
                mat_A[176][3] * mat_B[31][3] +
                mat_A[177][0] * mat_B[39][3] +
                mat_A[177][1] * mat_B[47][3] +
                mat_A[177][2] * mat_B[55][3] +
                mat_A[177][3] * mat_B[63][3] +
                mat_A[178][0] * mat_B[71][3] +
                mat_A[178][1] * mat_B[79][3] +
                mat_A[178][2] * mat_B[87][3] +
                mat_A[178][3] * mat_B[95][3] +
                mat_A[179][0] * mat_B[103][3] +
                mat_A[179][1] * mat_B[111][3] +
                mat_A[179][2] * mat_B[119][3] +
                mat_A[179][3] * mat_B[127][3] +
                mat_A[180][0] * mat_B[135][3] +
                mat_A[180][1] * mat_B[143][3] +
                mat_A[180][2] * mat_B[151][3] +
                mat_A[180][3] * mat_B[159][3] +
                mat_A[181][0] * mat_B[167][3] +
                mat_A[181][1] * mat_B[175][3] +
                mat_A[181][2] * mat_B[183][3] +
                mat_A[181][3] * mat_B[191][3] +
                mat_A[182][0] * mat_B[199][3] +
                mat_A[182][1] * mat_B[207][3] +
                mat_A[182][2] * mat_B[215][3] +
                mat_A[182][3] * mat_B[223][3] +
                mat_A[183][0] * mat_B[231][3] +
                mat_A[183][1] * mat_B[239][3] +
                mat_A[183][2] * mat_B[247][3] +
                mat_A[183][3] * mat_B[255][3];
    mat_C[184][0] <=
                mat_A[184][0] * mat_B[0][0] +
                mat_A[184][1] * mat_B[8][0] +
                mat_A[184][2] * mat_B[16][0] +
                mat_A[184][3] * mat_B[24][0] +
                mat_A[185][0] * mat_B[32][0] +
                mat_A[185][1] * mat_B[40][0] +
                mat_A[185][2] * mat_B[48][0] +
                mat_A[185][3] * mat_B[56][0] +
                mat_A[186][0] * mat_B[64][0] +
                mat_A[186][1] * mat_B[72][0] +
                mat_A[186][2] * mat_B[80][0] +
                mat_A[186][3] * mat_B[88][0] +
                mat_A[187][0] * mat_B[96][0] +
                mat_A[187][1] * mat_B[104][0] +
                mat_A[187][2] * mat_B[112][0] +
                mat_A[187][3] * mat_B[120][0] +
                mat_A[188][0] * mat_B[128][0] +
                mat_A[188][1] * mat_B[136][0] +
                mat_A[188][2] * mat_B[144][0] +
                mat_A[188][3] * mat_B[152][0] +
                mat_A[189][0] * mat_B[160][0] +
                mat_A[189][1] * mat_B[168][0] +
                mat_A[189][2] * mat_B[176][0] +
                mat_A[189][3] * mat_B[184][0] +
                mat_A[190][0] * mat_B[192][0] +
                mat_A[190][1] * mat_B[200][0] +
                mat_A[190][2] * mat_B[208][0] +
                mat_A[190][3] * mat_B[216][0] +
                mat_A[191][0] * mat_B[224][0] +
                mat_A[191][1] * mat_B[232][0] +
                mat_A[191][2] * mat_B[240][0] +
                mat_A[191][3] * mat_B[248][0];
    mat_C[184][1] <=
                mat_A[184][0] * mat_B[0][1] +
                mat_A[184][1] * mat_B[8][1] +
                mat_A[184][2] * mat_B[16][1] +
                mat_A[184][3] * mat_B[24][1] +
                mat_A[185][0] * mat_B[32][1] +
                mat_A[185][1] * mat_B[40][1] +
                mat_A[185][2] * mat_B[48][1] +
                mat_A[185][3] * mat_B[56][1] +
                mat_A[186][0] * mat_B[64][1] +
                mat_A[186][1] * mat_B[72][1] +
                mat_A[186][2] * mat_B[80][1] +
                mat_A[186][3] * mat_B[88][1] +
                mat_A[187][0] * mat_B[96][1] +
                mat_A[187][1] * mat_B[104][1] +
                mat_A[187][2] * mat_B[112][1] +
                mat_A[187][3] * mat_B[120][1] +
                mat_A[188][0] * mat_B[128][1] +
                mat_A[188][1] * mat_B[136][1] +
                mat_A[188][2] * mat_B[144][1] +
                mat_A[188][3] * mat_B[152][1] +
                mat_A[189][0] * mat_B[160][1] +
                mat_A[189][1] * mat_B[168][1] +
                mat_A[189][2] * mat_B[176][1] +
                mat_A[189][3] * mat_B[184][1] +
                mat_A[190][0] * mat_B[192][1] +
                mat_A[190][1] * mat_B[200][1] +
                mat_A[190][2] * mat_B[208][1] +
                mat_A[190][3] * mat_B[216][1] +
                mat_A[191][0] * mat_B[224][1] +
                mat_A[191][1] * mat_B[232][1] +
                mat_A[191][2] * mat_B[240][1] +
                mat_A[191][3] * mat_B[248][1];
    mat_C[184][2] <=
                mat_A[184][0] * mat_B[0][2] +
                mat_A[184][1] * mat_B[8][2] +
                mat_A[184][2] * mat_B[16][2] +
                mat_A[184][3] * mat_B[24][2] +
                mat_A[185][0] * mat_B[32][2] +
                mat_A[185][1] * mat_B[40][2] +
                mat_A[185][2] * mat_B[48][2] +
                mat_A[185][3] * mat_B[56][2] +
                mat_A[186][0] * mat_B[64][2] +
                mat_A[186][1] * mat_B[72][2] +
                mat_A[186][2] * mat_B[80][2] +
                mat_A[186][3] * mat_B[88][2] +
                mat_A[187][0] * mat_B[96][2] +
                mat_A[187][1] * mat_B[104][2] +
                mat_A[187][2] * mat_B[112][2] +
                mat_A[187][3] * mat_B[120][2] +
                mat_A[188][0] * mat_B[128][2] +
                mat_A[188][1] * mat_B[136][2] +
                mat_A[188][2] * mat_B[144][2] +
                mat_A[188][3] * mat_B[152][2] +
                mat_A[189][0] * mat_B[160][2] +
                mat_A[189][1] * mat_B[168][2] +
                mat_A[189][2] * mat_B[176][2] +
                mat_A[189][3] * mat_B[184][2] +
                mat_A[190][0] * mat_B[192][2] +
                mat_A[190][1] * mat_B[200][2] +
                mat_A[190][2] * mat_B[208][2] +
                mat_A[190][3] * mat_B[216][2] +
                mat_A[191][0] * mat_B[224][2] +
                mat_A[191][1] * mat_B[232][2] +
                mat_A[191][2] * mat_B[240][2] +
                mat_A[191][3] * mat_B[248][2];
    mat_C[184][3] <=
                mat_A[184][0] * mat_B[0][3] +
                mat_A[184][1] * mat_B[8][3] +
                mat_A[184][2] * mat_B[16][3] +
                mat_A[184][3] * mat_B[24][3] +
                mat_A[185][0] * mat_B[32][3] +
                mat_A[185][1] * mat_B[40][3] +
                mat_A[185][2] * mat_B[48][3] +
                mat_A[185][3] * mat_B[56][3] +
                mat_A[186][0] * mat_B[64][3] +
                mat_A[186][1] * mat_B[72][3] +
                mat_A[186][2] * mat_B[80][3] +
                mat_A[186][3] * mat_B[88][3] +
                mat_A[187][0] * mat_B[96][3] +
                mat_A[187][1] * mat_B[104][3] +
                mat_A[187][2] * mat_B[112][3] +
                mat_A[187][3] * mat_B[120][3] +
                mat_A[188][0] * mat_B[128][3] +
                mat_A[188][1] * mat_B[136][3] +
                mat_A[188][2] * mat_B[144][3] +
                mat_A[188][3] * mat_B[152][3] +
                mat_A[189][0] * mat_B[160][3] +
                mat_A[189][1] * mat_B[168][3] +
                mat_A[189][2] * mat_B[176][3] +
                mat_A[189][3] * mat_B[184][3] +
                mat_A[190][0] * mat_B[192][3] +
                mat_A[190][1] * mat_B[200][3] +
                mat_A[190][2] * mat_B[208][3] +
                mat_A[190][3] * mat_B[216][3] +
                mat_A[191][0] * mat_B[224][3] +
                mat_A[191][1] * mat_B[232][3] +
                mat_A[191][2] * mat_B[240][3] +
                mat_A[191][3] * mat_B[248][3];
    mat_C[185][0] <=
                mat_A[184][0] * mat_B[1][0] +
                mat_A[184][1] * mat_B[9][0] +
                mat_A[184][2] * mat_B[17][0] +
                mat_A[184][3] * mat_B[25][0] +
                mat_A[185][0] * mat_B[33][0] +
                mat_A[185][1] * mat_B[41][0] +
                mat_A[185][2] * mat_B[49][0] +
                mat_A[185][3] * mat_B[57][0] +
                mat_A[186][0] * mat_B[65][0] +
                mat_A[186][1] * mat_B[73][0] +
                mat_A[186][2] * mat_B[81][0] +
                mat_A[186][3] * mat_B[89][0] +
                mat_A[187][0] * mat_B[97][0] +
                mat_A[187][1] * mat_B[105][0] +
                mat_A[187][2] * mat_B[113][0] +
                mat_A[187][3] * mat_B[121][0] +
                mat_A[188][0] * mat_B[129][0] +
                mat_A[188][1] * mat_B[137][0] +
                mat_A[188][2] * mat_B[145][0] +
                mat_A[188][3] * mat_B[153][0] +
                mat_A[189][0] * mat_B[161][0] +
                mat_A[189][1] * mat_B[169][0] +
                mat_A[189][2] * mat_B[177][0] +
                mat_A[189][3] * mat_B[185][0] +
                mat_A[190][0] * mat_B[193][0] +
                mat_A[190][1] * mat_B[201][0] +
                mat_A[190][2] * mat_B[209][0] +
                mat_A[190][3] * mat_B[217][0] +
                mat_A[191][0] * mat_B[225][0] +
                mat_A[191][1] * mat_B[233][0] +
                mat_A[191][2] * mat_B[241][0] +
                mat_A[191][3] * mat_B[249][0];
    mat_C[185][1] <=
                mat_A[184][0] * mat_B[1][1] +
                mat_A[184][1] * mat_B[9][1] +
                mat_A[184][2] * mat_B[17][1] +
                mat_A[184][3] * mat_B[25][1] +
                mat_A[185][0] * mat_B[33][1] +
                mat_A[185][1] * mat_B[41][1] +
                mat_A[185][2] * mat_B[49][1] +
                mat_A[185][3] * mat_B[57][1] +
                mat_A[186][0] * mat_B[65][1] +
                mat_A[186][1] * mat_B[73][1] +
                mat_A[186][2] * mat_B[81][1] +
                mat_A[186][3] * mat_B[89][1] +
                mat_A[187][0] * mat_B[97][1] +
                mat_A[187][1] * mat_B[105][1] +
                mat_A[187][2] * mat_B[113][1] +
                mat_A[187][3] * mat_B[121][1] +
                mat_A[188][0] * mat_B[129][1] +
                mat_A[188][1] * mat_B[137][1] +
                mat_A[188][2] * mat_B[145][1] +
                mat_A[188][3] * mat_B[153][1] +
                mat_A[189][0] * mat_B[161][1] +
                mat_A[189][1] * mat_B[169][1] +
                mat_A[189][2] * mat_B[177][1] +
                mat_A[189][3] * mat_B[185][1] +
                mat_A[190][0] * mat_B[193][1] +
                mat_A[190][1] * mat_B[201][1] +
                mat_A[190][2] * mat_B[209][1] +
                mat_A[190][3] * mat_B[217][1] +
                mat_A[191][0] * mat_B[225][1] +
                mat_A[191][1] * mat_B[233][1] +
                mat_A[191][2] * mat_B[241][1] +
                mat_A[191][3] * mat_B[249][1];
    mat_C[185][2] <=
                mat_A[184][0] * mat_B[1][2] +
                mat_A[184][1] * mat_B[9][2] +
                mat_A[184][2] * mat_B[17][2] +
                mat_A[184][3] * mat_B[25][2] +
                mat_A[185][0] * mat_B[33][2] +
                mat_A[185][1] * mat_B[41][2] +
                mat_A[185][2] * mat_B[49][2] +
                mat_A[185][3] * mat_B[57][2] +
                mat_A[186][0] * mat_B[65][2] +
                mat_A[186][1] * mat_B[73][2] +
                mat_A[186][2] * mat_B[81][2] +
                mat_A[186][3] * mat_B[89][2] +
                mat_A[187][0] * mat_B[97][2] +
                mat_A[187][1] * mat_B[105][2] +
                mat_A[187][2] * mat_B[113][2] +
                mat_A[187][3] * mat_B[121][2] +
                mat_A[188][0] * mat_B[129][2] +
                mat_A[188][1] * mat_B[137][2] +
                mat_A[188][2] * mat_B[145][2] +
                mat_A[188][3] * mat_B[153][2] +
                mat_A[189][0] * mat_B[161][2] +
                mat_A[189][1] * mat_B[169][2] +
                mat_A[189][2] * mat_B[177][2] +
                mat_A[189][3] * mat_B[185][2] +
                mat_A[190][0] * mat_B[193][2] +
                mat_A[190][1] * mat_B[201][2] +
                mat_A[190][2] * mat_B[209][2] +
                mat_A[190][3] * mat_B[217][2] +
                mat_A[191][0] * mat_B[225][2] +
                mat_A[191][1] * mat_B[233][2] +
                mat_A[191][2] * mat_B[241][2] +
                mat_A[191][3] * mat_B[249][2];
    mat_C[185][3] <=
                mat_A[184][0] * mat_B[1][3] +
                mat_A[184][1] * mat_B[9][3] +
                mat_A[184][2] * mat_B[17][3] +
                mat_A[184][3] * mat_B[25][3] +
                mat_A[185][0] * mat_B[33][3] +
                mat_A[185][1] * mat_B[41][3] +
                mat_A[185][2] * mat_B[49][3] +
                mat_A[185][3] * mat_B[57][3] +
                mat_A[186][0] * mat_B[65][3] +
                mat_A[186][1] * mat_B[73][3] +
                mat_A[186][2] * mat_B[81][3] +
                mat_A[186][3] * mat_B[89][3] +
                mat_A[187][0] * mat_B[97][3] +
                mat_A[187][1] * mat_B[105][3] +
                mat_A[187][2] * mat_B[113][3] +
                mat_A[187][3] * mat_B[121][3] +
                mat_A[188][0] * mat_B[129][3] +
                mat_A[188][1] * mat_B[137][3] +
                mat_A[188][2] * mat_B[145][3] +
                mat_A[188][3] * mat_B[153][3] +
                mat_A[189][0] * mat_B[161][3] +
                mat_A[189][1] * mat_B[169][3] +
                mat_A[189][2] * mat_B[177][3] +
                mat_A[189][3] * mat_B[185][3] +
                mat_A[190][0] * mat_B[193][3] +
                mat_A[190][1] * mat_B[201][3] +
                mat_A[190][2] * mat_B[209][3] +
                mat_A[190][3] * mat_B[217][3] +
                mat_A[191][0] * mat_B[225][3] +
                mat_A[191][1] * mat_B[233][3] +
                mat_A[191][2] * mat_B[241][3] +
                mat_A[191][3] * mat_B[249][3];
    mat_C[186][0] <=
                mat_A[184][0] * mat_B[2][0] +
                mat_A[184][1] * mat_B[10][0] +
                mat_A[184][2] * mat_B[18][0] +
                mat_A[184][3] * mat_B[26][0] +
                mat_A[185][0] * mat_B[34][0] +
                mat_A[185][1] * mat_B[42][0] +
                mat_A[185][2] * mat_B[50][0] +
                mat_A[185][3] * mat_B[58][0] +
                mat_A[186][0] * mat_B[66][0] +
                mat_A[186][1] * mat_B[74][0] +
                mat_A[186][2] * mat_B[82][0] +
                mat_A[186][3] * mat_B[90][0] +
                mat_A[187][0] * mat_B[98][0] +
                mat_A[187][1] * mat_B[106][0] +
                mat_A[187][2] * mat_B[114][0] +
                mat_A[187][3] * mat_B[122][0] +
                mat_A[188][0] * mat_B[130][0] +
                mat_A[188][1] * mat_B[138][0] +
                mat_A[188][2] * mat_B[146][0] +
                mat_A[188][3] * mat_B[154][0] +
                mat_A[189][0] * mat_B[162][0] +
                mat_A[189][1] * mat_B[170][0] +
                mat_A[189][2] * mat_B[178][0] +
                mat_A[189][3] * mat_B[186][0] +
                mat_A[190][0] * mat_B[194][0] +
                mat_A[190][1] * mat_B[202][0] +
                mat_A[190][2] * mat_B[210][0] +
                mat_A[190][3] * mat_B[218][0] +
                mat_A[191][0] * mat_B[226][0] +
                mat_A[191][1] * mat_B[234][0] +
                mat_A[191][2] * mat_B[242][0] +
                mat_A[191][3] * mat_B[250][0];
    mat_C[186][1] <=
                mat_A[184][0] * mat_B[2][1] +
                mat_A[184][1] * mat_B[10][1] +
                mat_A[184][2] * mat_B[18][1] +
                mat_A[184][3] * mat_B[26][1] +
                mat_A[185][0] * mat_B[34][1] +
                mat_A[185][1] * mat_B[42][1] +
                mat_A[185][2] * mat_B[50][1] +
                mat_A[185][3] * mat_B[58][1] +
                mat_A[186][0] * mat_B[66][1] +
                mat_A[186][1] * mat_B[74][1] +
                mat_A[186][2] * mat_B[82][1] +
                mat_A[186][3] * mat_B[90][1] +
                mat_A[187][0] * mat_B[98][1] +
                mat_A[187][1] * mat_B[106][1] +
                mat_A[187][2] * mat_B[114][1] +
                mat_A[187][3] * mat_B[122][1] +
                mat_A[188][0] * mat_B[130][1] +
                mat_A[188][1] * mat_B[138][1] +
                mat_A[188][2] * mat_B[146][1] +
                mat_A[188][3] * mat_B[154][1] +
                mat_A[189][0] * mat_B[162][1] +
                mat_A[189][1] * mat_B[170][1] +
                mat_A[189][2] * mat_B[178][1] +
                mat_A[189][3] * mat_B[186][1] +
                mat_A[190][0] * mat_B[194][1] +
                mat_A[190][1] * mat_B[202][1] +
                mat_A[190][2] * mat_B[210][1] +
                mat_A[190][3] * mat_B[218][1] +
                mat_A[191][0] * mat_B[226][1] +
                mat_A[191][1] * mat_B[234][1] +
                mat_A[191][2] * mat_B[242][1] +
                mat_A[191][3] * mat_B[250][1];
    mat_C[186][2] <=
                mat_A[184][0] * mat_B[2][2] +
                mat_A[184][1] * mat_B[10][2] +
                mat_A[184][2] * mat_B[18][2] +
                mat_A[184][3] * mat_B[26][2] +
                mat_A[185][0] * mat_B[34][2] +
                mat_A[185][1] * mat_B[42][2] +
                mat_A[185][2] * mat_B[50][2] +
                mat_A[185][3] * mat_B[58][2] +
                mat_A[186][0] * mat_B[66][2] +
                mat_A[186][1] * mat_B[74][2] +
                mat_A[186][2] * mat_B[82][2] +
                mat_A[186][3] * mat_B[90][2] +
                mat_A[187][0] * mat_B[98][2] +
                mat_A[187][1] * mat_B[106][2] +
                mat_A[187][2] * mat_B[114][2] +
                mat_A[187][3] * mat_B[122][2] +
                mat_A[188][0] * mat_B[130][2] +
                mat_A[188][1] * mat_B[138][2] +
                mat_A[188][2] * mat_B[146][2] +
                mat_A[188][3] * mat_B[154][2] +
                mat_A[189][0] * mat_B[162][2] +
                mat_A[189][1] * mat_B[170][2] +
                mat_A[189][2] * mat_B[178][2] +
                mat_A[189][3] * mat_B[186][2] +
                mat_A[190][0] * mat_B[194][2] +
                mat_A[190][1] * mat_B[202][2] +
                mat_A[190][2] * mat_B[210][2] +
                mat_A[190][3] * mat_B[218][2] +
                mat_A[191][0] * mat_B[226][2] +
                mat_A[191][1] * mat_B[234][2] +
                mat_A[191][2] * mat_B[242][2] +
                mat_A[191][3] * mat_B[250][2];
    mat_C[186][3] <=
                mat_A[184][0] * mat_B[2][3] +
                mat_A[184][1] * mat_B[10][3] +
                mat_A[184][2] * mat_B[18][3] +
                mat_A[184][3] * mat_B[26][3] +
                mat_A[185][0] * mat_B[34][3] +
                mat_A[185][1] * mat_B[42][3] +
                mat_A[185][2] * mat_B[50][3] +
                mat_A[185][3] * mat_B[58][3] +
                mat_A[186][0] * mat_B[66][3] +
                mat_A[186][1] * mat_B[74][3] +
                mat_A[186][2] * mat_B[82][3] +
                mat_A[186][3] * mat_B[90][3] +
                mat_A[187][0] * mat_B[98][3] +
                mat_A[187][1] * mat_B[106][3] +
                mat_A[187][2] * mat_B[114][3] +
                mat_A[187][3] * mat_B[122][3] +
                mat_A[188][0] * mat_B[130][3] +
                mat_A[188][1] * mat_B[138][3] +
                mat_A[188][2] * mat_B[146][3] +
                mat_A[188][3] * mat_B[154][3] +
                mat_A[189][0] * mat_B[162][3] +
                mat_A[189][1] * mat_B[170][3] +
                mat_A[189][2] * mat_B[178][3] +
                mat_A[189][3] * mat_B[186][3] +
                mat_A[190][0] * mat_B[194][3] +
                mat_A[190][1] * mat_B[202][3] +
                mat_A[190][2] * mat_B[210][3] +
                mat_A[190][3] * mat_B[218][3] +
                mat_A[191][0] * mat_B[226][3] +
                mat_A[191][1] * mat_B[234][3] +
                mat_A[191][2] * mat_B[242][3] +
                mat_A[191][3] * mat_B[250][3];
    mat_C[187][0] <=
                mat_A[184][0] * mat_B[3][0] +
                mat_A[184][1] * mat_B[11][0] +
                mat_A[184][2] * mat_B[19][0] +
                mat_A[184][3] * mat_B[27][0] +
                mat_A[185][0] * mat_B[35][0] +
                mat_A[185][1] * mat_B[43][0] +
                mat_A[185][2] * mat_B[51][0] +
                mat_A[185][3] * mat_B[59][0] +
                mat_A[186][0] * mat_B[67][0] +
                mat_A[186][1] * mat_B[75][0] +
                mat_A[186][2] * mat_B[83][0] +
                mat_A[186][3] * mat_B[91][0] +
                mat_A[187][0] * mat_B[99][0] +
                mat_A[187][1] * mat_B[107][0] +
                mat_A[187][2] * mat_B[115][0] +
                mat_A[187][3] * mat_B[123][0] +
                mat_A[188][0] * mat_B[131][0] +
                mat_A[188][1] * mat_B[139][0] +
                mat_A[188][2] * mat_B[147][0] +
                mat_A[188][3] * mat_B[155][0] +
                mat_A[189][0] * mat_B[163][0] +
                mat_A[189][1] * mat_B[171][0] +
                mat_A[189][2] * mat_B[179][0] +
                mat_A[189][3] * mat_B[187][0] +
                mat_A[190][0] * mat_B[195][0] +
                mat_A[190][1] * mat_B[203][0] +
                mat_A[190][2] * mat_B[211][0] +
                mat_A[190][3] * mat_B[219][0] +
                mat_A[191][0] * mat_B[227][0] +
                mat_A[191][1] * mat_B[235][0] +
                mat_A[191][2] * mat_B[243][0] +
                mat_A[191][3] * mat_B[251][0];
    mat_C[187][1] <=
                mat_A[184][0] * mat_B[3][1] +
                mat_A[184][1] * mat_B[11][1] +
                mat_A[184][2] * mat_B[19][1] +
                mat_A[184][3] * mat_B[27][1] +
                mat_A[185][0] * mat_B[35][1] +
                mat_A[185][1] * mat_B[43][1] +
                mat_A[185][2] * mat_B[51][1] +
                mat_A[185][3] * mat_B[59][1] +
                mat_A[186][0] * mat_B[67][1] +
                mat_A[186][1] * mat_B[75][1] +
                mat_A[186][2] * mat_B[83][1] +
                mat_A[186][3] * mat_B[91][1] +
                mat_A[187][0] * mat_B[99][1] +
                mat_A[187][1] * mat_B[107][1] +
                mat_A[187][2] * mat_B[115][1] +
                mat_A[187][3] * mat_B[123][1] +
                mat_A[188][0] * mat_B[131][1] +
                mat_A[188][1] * mat_B[139][1] +
                mat_A[188][2] * mat_B[147][1] +
                mat_A[188][3] * mat_B[155][1] +
                mat_A[189][0] * mat_B[163][1] +
                mat_A[189][1] * mat_B[171][1] +
                mat_A[189][2] * mat_B[179][1] +
                mat_A[189][3] * mat_B[187][1] +
                mat_A[190][0] * mat_B[195][1] +
                mat_A[190][1] * mat_B[203][1] +
                mat_A[190][2] * mat_B[211][1] +
                mat_A[190][3] * mat_B[219][1] +
                mat_A[191][0] * mat_B[227][1] +
                mat_A[191][1] * mat_B[235][1] +
                mat_A[191][2] * mat_B[243][1] +
                mat_A[191][3] * mat_B[251][1];
    mat_C[187][2] <=
                mat_A[184][0] * mat_B[3][2] +
                mat_A[184][1] * mat_B[11][2] +
                mat_A[184][2] * mat_B[19][2] +
                mat_A[184][3] * mat_B[27][2] +
                mat_A[185][0] * mat_B[35][2] +
                mat_A[185][1] * mat_B[43][2] +
                mat_A[185][2] * mat_B[51][2] +
                mat_A[185][3] * mat_B[59][2] +
                mat_A[186][0] * mat_B[67][2] +
                mat_A[186][1] * mat_B[75][2] +
                mat_A[186][2] * mat_B[83][2] +
                mat_A[186][3] * mat_B[91][2] +
                mat_A[187][0] * mat_B[99][2] +
                mat_A[187][1] * mat_B[107][2] +
                mat_A[187][2] * mat_B[115][2] +
                mat_A[187][3] * mat_B[123][2] +
                mat_A[188][0] * mat_B[131][2] +
                mat_A[188][1] * mat_B[139][2] +
                mat_A[188][2] * mat_B[147][2] +
                mat_A[188][3] * mat_B[155][2] +
                mat_A[189][0] * mat_B[163][2] +
                mat_A[189][1] * mat_B[171][2] +
                mat_A[189][2] * mat_B[179][2] +
                mat_A[189][3] * mat_B[187][2] +
                mat_A[190][0] * mat_B[195][2] +
                mat_A[190][1] * mat_B[203][2] +
                mat_A[190][2] * mat_B[211][2] +
                mat_A[190][3] * mat_B[219][2] +
                mat_A[191][0] * mat_B[227][2] +
                mat_A[191][1] * mat_B[235][2] +
                mat_A[191][2] * mat_B[243][2] +
                mat_A[191][3] * mat_B[251][2];
    mat_C[187][3] <=
                mat_A[184][0] * mat_B[3][3] +
                mat_A[184][1] * mat_B[11][3] +
                mat_A[184][2] * mat_B[19][3] +
                mat_A[184][3] * mat_B[27][3] +
                mat_A[185][0] * mat_B[35][3] +
                mat_A[185][1] * mat_B[43][3] +
                mat_A[185][2] * mat_B[51][3] +
                mat_A[185][3] * mat_B[59][3] +
                mat_A[186][0] * mat_B[67][3] +
                mat_A[186][1] * mat_B[75][3] +
                mat_A[186][2] * mat_B[83][3] +
                mat_A[186][3] * mat_B[91][3] +
                mat_A[187][0] * mat_B[99][3] +
                mat_A[187][1] * mat_B[107][3] +
                mat_A[187][2] * mat_B[115][3] +
                mat_A[187][3] * mat_B[123][3] +
                mat_A[188][0] * mat_B[131][3] +
                mat_A[188][1] * mat_B[139][3] +
                mat_A[188][2] * mat_B[147][3] +
                mat_A[188][3] * mat_B[155][3] +
                mat_A[189][0] * mat_B[163][3] +
                mat_A[189][1] * mat_B[171][3] +
                mat_A[189][2] * mat_B[179][3] +
                mat_A[189][3] * mat_B[187][3] +
                mat_A[190][0] * mat_B[195][3] +
                mat_A[190][1] * mat_B[203][3] +
                mat_A[190][2] * mat_B[211][3] +
                mat_A[190][3] * mat_B[219][3] +
                mat_A[191][0] * mat_B[227][3] +
                mat_A[191][1] * mat_B[235][3] +
                mat_A[191][2] * mat_B[243][3] +
                mat_A[191][3] * mat_B[251][3];
    mat_C[188][0] <=
                mat_A[184][0] * mat_B[4][0] +
                mat_A[184][1] * mat_B[12][0] +
                mat_A[184][2] * mat_B[20][0] +
                mat_A[184][3] * mat_B[28][0] +
                mat_A[185][0] * mat_B[36][0] +
                mat_A[185][1] * mat_B[44][0] +
                mat_A[185][2] * mat_B[52][0] +
                mat_A[185][3] * mat_B[60][0] +
                mat_A[186][0] * mat_B[68][0] +
                mat_A[186][1] * mat_B[76][0] +
                mat_A[186][2] * mat_B[84][0] +
                mat_A[186][3] * mat_B[92][0] +
                mat_A[187][0] * mat_B[100][0] +
                mat_A[187][1] * mat_B[108][0] +
                mat_A[187][2] * mat_B[116][0] +
                mat_A[187][3] * mat_B[124][0] +
                mat_A[188][0] * mat_B[132][0] +
                mat_A[188][1] * mat_B[140][0] +
                mat_A[188][2] * mat_B[148][0] +
                mat_A[188][3] * mat_B[156][0] +
                mat_A[189][0] * mat_B[164][0] +
                mat_A[189][1] * mat_B[172][0] +
                mat_A[189][2] * mat_B[180][0] +
                mat_A[189][3] * mat_B[188][0] +
                mat_A[190][0] * mat_B[196][0] +
                mat_A[190][1] * mat_B[204][0] +
                mat_A[190][2] * mat_B[212][0] +
                mat_A[190][3] * mat_B[220][0] +
                mat_A[191][0] * mat_B[228][0] +
                mat_A[191][1] * mat_B[236][0] +
                mat_A[191][2] * mat_B[244][0] +
                mat_A[191][3] * mat_B[252][0];
    mat_C[188][1] <=
                mat_A[184][0] * mat_B[4][1] +
                mat_A[184][1] * mat_B[12][1] +
                mat_A[184][2] * mat_B[20][1] +
                mat_A[184][3] * mat_B[28][1] +
                mat_A[185][0] * mat_B[36][1] +
                mat_A[185][1] * mat_B[44][1] +
                mat_A[185][2] * mat_B[52][1] +
                mat_A[185][3] * mat_B[60][1] +
                mat_A[186][0] * mat_B[68][1] +
                mat_A[186][1] * mat_B[76][1] +
                mat_A[186][2] * mat_B[84][1] +
                mat_A[186][3] * mat_B[92][1] +
                mat_A[187][0] * mat_B[100][1] +
                mat_A[187][1] * mat_B[108][1] +
                mat_A[187][2] * mat_B[116][1] +
                mat_A[187][3] * mat_B[124][1] +
                mat_A[188][0] * mat_B[132][1] +
                mat_A[188][1] * mat_B[140][1] +
                mat_A[188][2] * mat_B[148][1] +
                mat_A[188][3] * mat_B[156][1] +
                mat_A[189][0] * mat_B[164][1] +
                mat_A[189][1] * mat_B[172][1] +
                mat_A[189][2] * mat_B[180][1] +
                mat_A[189][3] * mat_B[188][1] +
                mat_A[190][0] * mat_B[196][1] +
                mat_A[190][1] * mat_B[204][1] +
                mat_A[190][2] * mat_B[212][1] +
                mat_A[190][3] * mat_B[220][1] +
                mat_A[191][0] * mat_B[228][1] +
                mat_A[191][1] * mat_B[236][1] +
                mat_A[191][2] * mat_B[244][1] +
                mat_A[191][3] * mat_B[252][1];
    mat_C[188][2] <=
                mat_A[184][0] * mat_B[4][2] +
                mat_A[184][1] * mat_B[12][2] +
                mat_A[184][2] * mat_B[20][2] +
                mat_A[184][3] * mat_B[28][2] +
                mat_A[185][0] * mat_B[36][2] +
                mat_A[185][1] * mat_B[44][2] +
                mat_A[185][2] * mat_B[52][2] +
                mat_A[185][3] * mat_B[60][2] +
                mat_A[186][0] * mat_B[68][2] +
                mat_A[186][1] * mat_B[76][2] +
                mat_A[186][2] * mat_B[84][2] +
                mat_A[186][3] * mat_B[92][2] +
                mat_A[187][0] * mat_B[100][2] +
                mat_A[187][1] * mat_B[108][2] +
                mat_A[187][2] * mat_B[116][2] +
                mat_A[187][3] * mat_B[124][2] +
                mat_A[188][0] * mat_B[132][2] +
                mat_A[188][1] * mat_B[140][2] +
                mat_A[188][2] * mat_B[148][2] +
                mat_A[188][3] * mat_B[156][2] +
                mat_A[189][0] * mat_B[164][2] +
                mat_A[189][1] * mat_B[172][2] +
                mat_A[189][2] * mat_B[180][2] +
                mat_A[189][3] * mat_B[188][2] +
                mat_A[190][0] * mat_B[196][2] +
                mat_A[190][1] * mat_B[204][2] +
                mat_A[190][2] * mat_B[212][2] +
                mat_A[190][3] * mat_B[220][2] +
                mat_A[191][0] * mat_B[228][2] +
                mat_A[191][1] * mat_B[236][2] +
                mat_A[191][2] * mat_B[244][2] +
                mat_A[191][3] * mat_B[252][2];
    mat_C[188][3] <=
                mat_A[184][0] * mat_B[4][3] +
                mat_A[184][1] * mat_B[12][3] +
                mat_A[184][2] * mat_B[20][3] +
                mat_A[184][3] * mat_B[28][3] +
                mat_A[185][0] * mat_B[36][3] +
                mat_A[185][1] * mat_B[44][3] +
                mat_A[185][2] * mat_B[52][3] +
                mat_A[185][3] * mat_B[60][3] +
                mat_A[186][0] * mat_B[68][3] +
                mat_A[186][1] * mat_B[76][3] +
                mat_A[186][2] * mat_B[84][3] +
                mat_A[186][3] * mat_B[92][3] +
                mat_A[187][0] * mat_B[100][3] +
                mat_A[187][1] * mat_B[108][3] +
                mat_A[187][2] * mat_B[116][3] +
                mat_A[187][3] * mat_B[124][3] +
                mat_A[188][0] * mat_B[132][3] +
                mat_A[188][1] * mat_B[140][3] +
                mat_A[188][2] * mat_B[148][3] +
                mat_A[188][3] * mat_B[156][3] +
                mat_A[189][0] * mat_B[164][3] +
                mat_A[189][1] * mat_B[172][3] +
                mat_A[189][2] * mat_B[180][3] +
                mat_A[189][3] * mat_B[188][3] +
                mat_A[190][0] * mat_B[196][3] +
                mat_A[190][1] * mat_B[204][3] +
                mat_A[190][2] * mat_B[212][3] +
                mat_A[190][3] * mat_B[220][3] +
                mat_A[191][0] * mat_B[228][3] +
                mat_A[191][1] * mat_B[236][3] +
                mat_A[191][2] * mat_B[244][3] +
                mat_A[191][3] * mat_B[252][3];
    mat_C[189][0] <=
                mat_A[184][0] * mat_B[5][0] +
                mat_A[184][1] * mat_B[13][0] +
                mat_A[184][2] * mat_B[21][0] +
                mat_A[184][3] * mat_B[29][0] +
                mat_A[185][0] * mat_B[37][0] +
                mat_A[185][1] * mat_B[45][0] +
                mat_A[185][2] * mat_B[53][0] +
                mat_A[185][3] * mat_B[61][0] +
                mat_A[186][0] * mat_B[69][0] +
                mat_A[186][1] * mat_B[77][0] +
                mat_A[186][2] * mat_B[85][0] +
                mat_A[186][3] * mat_B[93][0] +
                mat_A[187][0] * mat_B[101][0] +
                mat_A[187][1] * mat_B[109][0] +
                mat_A[187][2] * mat_B[117][0] +
                mat_A[187][3] * mat_B[125][0] +
                mat_A[188][0] * mat_B[133][0] +
                mat_A[188][1] * mat_B[141][0] +
                mat_A[188][2] * mat_B[149][0] +
                mat_A[188][3] * mat_B[157][0] +
                mat_A[189][0] * mat_B[165][0] +
                mat_A[189][1] * mat_B[173][0] +
                mat_A[189][2] * mat_B[181][0] +
                mat_A[189][3] * mat_B[189][0] +
                mat_A[190][0] * mat_B[197][0] +
                mat_A[190][1] * mat_B[205][0] +
                mat_A[190][2] * mat_B[213][0] +
                mat_A[190][3] * mat_B[221][0] +
                mat_A[191][0] * mat_B[229][0] +
                mat_A[191][1] * mat_B[237][0] +
                mat_A[191][2] * mat_B[245][0] +
                mat_A[191][3] * mat_B[253][0];
    mat_C[189][1] <=
                mat_A[184][0] * mat_B[5][1] +
                mat_A[184][1] * mat_B[13][1] +
                mat_A[184][2] * mat_B[21][1] +
                mat_A[184][3] * mat_B[29][1] +
                mat_A[185][0] * mat_B[37][1] +
                mat_A[185][1] * mat_B[45][1] +
                mat_A[185][2] * mat_B[53][1] +
                mat_A[185][3] * mat_B[61][1] +
                mat_A[186][0] * mat_B[69][1] +
                mat_A[186][1] * mat_B[77][1] +
                mat_A[186][2] * mat_B[85][1] +
                mat_A[186][3] * mat_B[93][1] +
                mat_A[187][0] * mat_B[101][1] +
                mat_A[187][1] * mat_B[109][1] +
                mat_A[187][2] * mat_B[117][1] +
                mat_A[187][3] * mat_B[125][1] +
                mat_A[188][0] * mat_B[133][1] +
                mat_A[188][1] * mat_B[141][1] +
                mat_A[188][2] * mat_B[149][1] +
                mat_A[188][3] * mat_B[157][1] +
                mat_A[189][0] * mat_B[165][1] +
                mat_A[189][1] * mat_B[173][1] +
                mat_A[189][2] * mat_B[181][1] +
                mat_A[189][3] * mat_B[189][1] +
                mat_A[190][0] * mat_B[197][1] +
                mat_A[190][1] * mat_B[205][1] +
                mat_A[190][2] * mat_B[213][1] +
                mat_A[190][3] * mat_B[221][1] +
                mat_A[191][0] * mat_B[229][1] +
                mat_A[191][1] * mat_B[237][1] +
                mat_A[191][2] * mat_B[245][1] +
                mat_A[191][3] * mat_B[253][1];
    mat_C[189][2] <=
                mat_A[184][0] * mat_B[5][2] +
                mat_A[184][1] * mat_B[13][2] +
                mat_A[184][2] * mat_B[21][2] +
                mat_A[184][3] * mat_B[29][2] +
                mat_A[185][0] * mat_B[37][2] +
                mat_A[185][1] * mat_B[45][2] +
                mat_A[185][2] * mat_B[53][2] +
                mat_A[185][3] * mat_B[61][2] +
                mat_A[186][0] * mat_B[69][2] +
                mat_A[186][1] * mat_B[77][2] +
                mat_A[186][2] * mat_B[85][2] +
                mat_A[186][3] * mat_B[93][2] +
                mat_A[187][0] * mat_B[101][2] +
                mat_A[187][1] * mat_B[109][2] +
                mat_A[187][2] * mat_B[117][2] +
                mat_A[187][3] * mat_B[125][2] +
                mat_A[188][0] * mat_B[133][2] +
                mat_A[188][1] * mat_B[141][2] +
                mat_A[188][2] * mat_B[149][2] +
                mat_A[188][3] * mat_B[157][2] +
                mat_A[189][0] * mat_B[165][2] +
                mat_A[189][1] * mat_B[173][2] +
                mat_A[189][2] * mat_B[181][2] +
                mat_A[189][3] * mat_B[189][2] +
                mat_A[190][0] * mat_B[197][2] +
                mat_A[190][1] * mat_B[205][2] +
                mat_A[190][2] * mat_B[213][2] +
                mat_A[190][3] * mat_B[221][2] +
                mat_A[191][0] * mat_B[229][2] +
                mat_A[191][1] * mat_B[237][2] +
                mat_A[191][2] * mat_B[245][2] +
                mat_A[191][3] * mat_B[253][2];
    mat_C[189][3] <=
                mat_A[184][0] * mat_B[5][3] +
                mat_A[184][1] * mat_B[13][3] +
                mat_A[184][2] * mat_B[21][3] +
                mat_A[184][3] * mat_B[29][3] +
                mat_A[185][0] * mat_B[37][3] +
                mat_A[185][1] * mat_B[45][3] +
                mat_A[185][2] * mat_B[53][3] +
                mat_A[185][3] * mat_B[61][3] +
                mat_A[186][0] * mat_B[69][3] +
                mat_A[186][1] * mat_B[77][3] +
                mat_A[186][2] * mat_B[85][3] +
                mat_A[186][3] * mat_B[93][3] +
                mat_A[187][0] * mat_B[101][3] +
                mat_A[187][1] * mat_B[109][3] +
                mat_A[187][2] * mat_B[117][3] +
                mat_A[187][3] * mat_B[125][3] +
                mat_A[188][0] * mat_B[133][3] +
                mat_A[188][1] * mat_B[141][3] +
                mat_A[188][2] * mat_B[149][3] +
                mat_A[188][3] * mat_B[157][3] +
                mat_A[189][0] * mat_B[165][3] +
                mat_A[189][1] * mat_B[173][3] +
                mat_A[189][2] * mat_B[181][3] +
                mat_A[189][3] * mat_B[189][3] +
                mat_A[190][0] * mat_B[197][3] +
                mat_A[190][1] * mat_B[205][3] +
                mat_A[190][2] * mat_B[213][3] +
                mat_A[190][3] * mat_B[221][3] +
                mat_A[191][0] * mat_B[229][3] +
                mat_A[191][1] * mat_B[237][3] +
                mat_A[191][2] * mat_B[245][3] +
                mat_A[191][3] * mat_B[253][3];
    mat_C[190][0] <=
                mat_A[184][0] * mat_B[6][0] +
                mat_A[184][1] * mat_B[14][0] +
                mat_A[184][2] * mat_B[22][0] +
                mat_A[184][3] * mat_B[30][0] +
                mat_A[185][0] * mat_B[38][0] +
                mat_A[185][1] * mat_B[46][0] +
                mat_A[185][2] * mat_B[54][0] +
                mat_A[185][3] * mat_B[62][0] +
                mat_A[186][0] * mat_B[70][0] +
                mat_A[186][1] * mat_B[78][0] +
                mat_A[186][2] * mat_B[86][0] +
                mat_A[186][3] * mat_B[94][0] +
                mat_A[187][0] * mat_B[102][0] +
                mat_A[187][1] * mat_B[110][0] +
                mat_A[187][2] * mat_B[118][0] +
                mat_A[187][3] * mat_B[126][0] +
                mat_A[188][0] * mat_B[134][0] +
                mat_A[188][1] * mat_B[142][0] +
                mat_A[188][2] * mat_B[150][0] +
                mat_A[188][3] * mat_B[158][0] +
                mat_A[189][0] * mat_B[166][0] +
                mat_A[189][1] * mat_B[174][0] +
                mat_A[189][2] * mat_B[182][0] +
                mat_A[189][3] * mat_B[190][0] +
                mat_A[190][0] * mat_B[198][0] +
                mat_A[190][1] * mat_B[206][0] +
                mat_A[190][2] * mat_B[214][0] +
                mat_A[190][3] * mat_B[222][0] +
                mat_A[191][0] * mat_B[230][0] +
                mat_A[191][1] * mat_B[238][0] +
                mat_A[191][2] * mat_B[246][0] +
                mat_A[191][3] * mat_B[254][0];
    mat_C[190][1] <=
                mat_A[184][0] * mat_B[6][1] +
                mat_A[184][1] * mat_B[14][1] +
                mat_A[184][2] * mat_B[22][1] +
                mat_A[184][3] * mat_B[30][1] +
                mat_A[185][0] * mat_B[38][1] +
                mat_A[185][1] * mat_B[46][1] +
                mat_A[185][2] * mat_B[54][1] +
                mat_A[185][3] * mat_B[62][1] +
                mat_A[186][0] * mat_B[70][1] +
                mat_A[186][1] * mat_B[78][1] +
                mat_A[186][2] * mat_B[86][1] +
                mat_A[186][3] * mat_B[94][1] +
                mat_A[187][0] * mat_B[102][1] +
                mat_A[187][1] * mat_B[110][1] +
                mat_A[187][2] * mat_B[118][1] +
                mat_A[187][3] * mat_B[126][1] +
                mat_A[188][0] * mat_B[134][1] +
                mat_A[188][1] * mat_B[142][1] +
                mat_A[188][2] * mat_B[150][1] +
                mat_A[188][3] * mat_B[158][1] +
                mat_A[189][0] * mat_B[166][1] +
                mat_A[189][1] * mat_B[174][1] +
                mat_A[189][2] * mat_B[182][1] +
                mat_A[189][3] * mat_B[190][1] +
                mat_A[190][0] * mat_B[198][1] +
                mat_A[190][1] * mat_B[206][1] +
                mat_A[190][2] * mat_B[214][1] +
                mat_A[190][3] * mat_B[222][1] +
                mat_A[191][0] * mat_B[230][1] +
                mat_A[191][1] * mat_B[238][1] +
                mat_A[191][2] * mat_B[246][1] +
                mat_A[191][3] * mat_B[254][1];
    mat_C[190][2] <=
                mat_A[184][0] * mat_B[6][2] +
                mat_A[184][1] * mat_B[14][2] +
                mat_A[184][2] * mat_B[22][2] +
                mat_A[184][3] * mat_B[30][2] +
                mat_A[185][0] * mat_B[38][2] +
                mat_A[185][1] * mat_B[46][2] +
                mat_A[185][2] * mat_B[54][2] +
                mat_A[185][3] * mat_B[62][2] +
                mat_A[186][0] * mat_B[70][2] +
                mat_A[186][1] * mat_B[78][2] +
                mat_A[186][2] * mat_B[86][2] +
                mat_A[186][3] * mat_B[94][2] +
                mat_A[187][0] * mat_B[102][2] +
                mat_A[187][1] * mat_B[110][2] +
                mat_A[187][2] * mat_B[118][2] +
                mat_A[187][3] * mat_B[126][2] +
                mat_A[188][0] * mat_B[134][2] +
                mat_A[188][1] * mat_B[142][2] +
                mat_A[188][2] * mat_B[150][2] +
                mat_A[188][3] * mat_B[158][2] +
                mat_A[189][0] * mat_B[166][2] +
                mat_A[189][1] * mat_B[174][2] +
                mat_A[189][2] * mat_B[182][2] +
                mat_A[189][3] * mat_B[190][2] +
                mat_A[190][0] * mat_B[198][2] +
                mat_A[190][1] * mat_B[206][2] +
                mat_A[190][2] * mat_B[214][2] +
                mat_A[190][3] * mat_B[222][2] +
                mat_A[191][0] * mat_B[230][2] +
                mat_A[191][1] * mat_B[238][2] +
                mat_A[191][2] * mat_B[246][2] +
                mat_A[191][3] * mat_B[254][2];
    mat_C[190][3] <=
                mat_A[184][0] * mat_B[6][3] +
                mat_A[184][1] * mat_B[14][3] +
                mat_A[184][2] * mat_B[22][3] +
                mat_A[184][3] * mat_B[30][3] +
                mat_A[185][0] * mat_B[38][3] +
                mat_A[185][1] * mat_B[46][3] +
                mat_A[185][2] * mat_B[54][3] +
                mat_A[185][3] * mat_B[62][3] +
                mat_A[186][0] * mat_B[70][3] +
                mat_A[186][1] * mat_B[78][3] +
                mat_A[186][2] * mat_B[86][3] +
                mat_A[186][3] * mat_B[94][3] +
                mat_A[187][0] * mat_B[102][3] +
                mat_A[187][1] * mat_B[110][3] +
                mat_A[187][2] * mat_B[118][3] +
                mat_A[187][3] * mat_B[126][3] +
                mat_A[188][0] * mat_B[134][3] +
                mat_A[188][1] * mat_B[142][3] +
                mat_A[188][2] * mat_B[150][3] +
                mat_A[188][3] * mat_B[158][3] +
                mat_A[189][0] * mat_B[166][3] +
                mat_A[189][1] * mat_B[174][3] +
                mat_A[189][2] * mat_B[182][3] +
                mat_A[189][3] * mat_B[190][3] +
                mat_A[190][0] * mat_B[198][3] +
                mat_A[190][1] * mat_B[206][3] +
                mat_A[190][2] * mat_B[214][3] +
                mat_A[190][3] * mat_B[222][3] +
                mat_A[191][0] * mat_B[230][3] +
                mat_A[191][1] * mat_B[238][3] +
                mat_A[191][2] * mat_B[246][3] +
                mat_A[191][3] * mat_B[254][3];
    mat_C[191][0] <=
                mat_A[184][0] * mat_B[7][0] +
                mat_A[184][1] * mat_B[15][0] +
                mat_A[184][2] * mat_B[23][0] +
                mat_A[184][3] * mat_B[31][0] +
                mat_A[185][0] * mat_B[39][0] +
                mat_A[185][1] * mat_B[47][0] +
                mat_A[185][2] * mat_B[55][0] +
                mat_A[185][3] * mat_B[63][0] +
                mat_A[186][0] * mat_B[71][0] +
                mat_A[186][1] * mat_B[79][0] +
                mat_A[186][2] * mat_B[87][0] +
                mat_A[186][3] * mat_B[95][0] +
                mat_A[187][0] * mat_B[103][0] +
                mat_A[187][1] * mat_B[111][0] +
                mat_A[187][2] * mat_B[119][0] +
                mat_A[187][3] * mat_B[127][0] +
                mat_A[188][0] * mat_B[135][0] +
                mat_A[188][1] * mat_B[143][0] +
                mat_A[188][2] * mat_B[151][0] +
                mat_A[188][3] * mat_B[159][0] +
                mat_A[189][0] * mat_B[167][0] +
                mat_A[189][1] * mat_B[175][0] +
                mat_A[189][2] * mat_B[183][0] +
                mat_A[189][3] * mat_B[191][0] +
                mat_A[190][0] * mat_B[199][0] +
                mat_A[190][1] * mat_B[207][0] +
                mat_A[190][2] * mat_B[215][0] +
                mat_A[190][3] * mat_B[223][0] +
                mat_A[191][0] * mat_B[231][0] +
                mat_A[191][1] * mat_B[239][0] +
                mat_A[191][2] * mat_B[247][0] +
                mat_A[191][3] * mat_B[255][0];
    mat_C[191][1] <=
                mat_A[184][0] * mat_B[7][1] +
                mat_A[184][1] * mat_B[15][1] +
                mat_A[184][2] * mat_B[23][1] +
                mat_A[184][3] * mat_B[31][1] +
                mat_A[185][0] * mat_B[39][1] +
                mat_A[185][1] * mat_B[47][1] +
                mat_A[185][2] * mat_B[55][1] +
                mat_A[185][3] * mat_B[63][1] +
                mat_A[186][0] * mat_B[71][1] +
                mat_A[186][1] * mat_B[79][1] +
                mat_A[186][2] * mat_B[87][1] +
                mat_A[186][3] * mat_B[95][1] +
                mat_A[187][0] * mat_B[103][1] +
                mat_A[187][1] * mat_B[111][1] +
                mat_A[187][2] * mat_B[119][1] +
                mat_A[187][3] * mat_B[127][1] +
                mat_A[188][0] * mat_B[135][1] +
                mat_A[188][1] * mat_B[143][1] +
                mat_A[188][2] * mat_B[151][1] +
                mat_A[188][3] * mat_B[159][1] +
                mat_A[189][0] * mat_B[167][1] +
                mat_A[189][1] * mat_B[175][1] +
                mat_A[189][2] * mat_B[183][1] +
                mat_A[189][3] * mat_B[191][1] +
                mat_A[190][0] * mat_B[199][1] +
                mat_A[190][1] * mat_B[207][1] +
                mat_A[190][2] * mat_B[215][1] +
                mat_A[190][3] * mat_B[223][1] +
                mat_A[191][0] * mat_B[231][1] +
                mat_A[191][1] * mat_B[239][1] +
                mat_A[191][2] * mat_B[247][1] +
                mat_A[191][3] * mat_B[255][1];
    mat_C[191][2] <=
                mat_A[184][0] * mat_B[7][2] +
                mat_A[184][1] * mat_B[15][2] +
                mat_A[184][2] * mat_B[23][2] +
                mat_A[184][3] * mat_B[31][2] +
                mat_A[185][0] * mat_B[39][2] +
                mat_A[185][1] * mat_B[47][2] +
                mat_A[185][2] * mat_B[55][2] +
                mat_A[185][3] * mat_B[63][2] +
                mat_A[186][0] * mat_B[71][2] +
                mat_A[186][1] * mat_B[79][2] +
                mat_A[186][2] * mat_B[87][2] +
                mat_A[186][3] * mat_B[95][2] +
                mat_A[187][0] * mat_B[103][2] +
                mat_A[187][1] * mat_B[111][2] +
                mat_A[187][2] * mat_B[119][2] +
                mat_A[187][3] * mat_B[127][2] +
                mat_A[188][0] * mat_B[135][2] +
                mat_A[188][1] * mat_B[143][2] +
                mat_A[188][2] * mat_B[151][2] +
                mat_A[188][3] * mat_B[159][2] +
                mat_A[189][0] * mat_B[167][2] +
                mat_A[189][1] * mat_B[175][2] +
                mat_A[189][2] * mat_B[183][2] +
                mat_A[189][3] * mat_B[191][2] +
                mat_A[190][0] * mat_B[199][2] +
                mat_A[190][1] * mat_B[207][2] +
                mat_A[190][2] * mat_B[215][2] +
                mat_A[190][3] * mat_B[223][2] +
                mat_A[191][0] * mat_B[231][2] +
                mat_A[191][1] * mat_B[239][2] +
                mat_A[191][2] * mat_B[247][2] +
                mat_A[191][3] * mat_B[255][2];
    mat_C[191][3] <=
                mat_A[184][0] * mat_B[7][3] +
                mat_A[184][1] * mat_B[15][3] +
                mat_A[184][2] * mat_B[23][3] +
                mat_A[184][3] * mat_B[31][3] +
                mat_A[185][0] * mat_B[39][3] +
                mat_A[185][1] * mat_B[47][3] +
                mat_A[185][2] * mat_B[55][3] +
                mat_A[185][3] * mat_B[63][3] +
                mat_A[186][0] * mat_B[71][3] +
                mat_A[186][1] * mat_B[79][3] +
                mat_A[186][2] * mat_B[87][3] +
                mat_A[186][3] * mat_B[95][3] +
                mat_A[187][0] * mat_B[103][3] +
                mat_A[187][1] * mat_B[111][3] +
                mat_A[187][2] * mat_B[119][3] +
                mat_A[187][3] * mat_B[127][3] +
                mat_A[188][0] * mat_B[135][3] +
                mat_A[188][1] * mat_B[143][3] +
                mat_A[188][2] * mat_B[151][3] +
                mat_A[188][3] * mat_B[159][3] +
                mat_A[189][0] * mat_B[167][3] +
                mat_A[189][1] * mat_B[175][3] +
                mat_A[189][2] * mat_B[183][3] +
                mat_A[189][3] * mat_B[191][3] +
                mat_A[190][0] * mat_B[199][3] +
                mat_A[190][1] * mat_B[207][3] +
                mat_A[190][2] * mat_B[215][3] +
                mat_A[190][3] * mat_B[223][3] +
                mat_A[191][0] * mat_B[231][3] +
                mat_A[191][1] * mat_B[239][3] +
                mat_A[191][2] * mat_B[247][3] +
                mat_A[191][3] * mat_B[255][3];
    mat_C[192][0] <=
                mat_A[192][0] * mat_B[0][0] +
                mat_A[192][1] * mat_B[8][0] +
                mat_A[192][2] * mat_B[16][0] +
                mat_A[192][3] * mat_B[24][0] +
                mat_A[193][0] * mat_B[32][0] +
                mat_A[193][1] * mat_B[40][0] +
                mat_A[193][2] * mat_B[48][0] +
                mat_A[193][3] * mat_B[56][0] +
                mat_A[194][0] * mat_B[64][0] +
                mat_A[194][1] * mat_B[72][0] +
                mat_A[194][2] * mat_B[80][0] +
                mat_A[194][3] * mat_B[88][0] +
                mat_A[195][0] * mat_B[96][0] +
                mat_A[195][1] * mat_B[104][0] +
                mat_A[195][2] * mat_B[112][0] +
                mat_A[195][3] * mat_B[120][0] +
                mat_A[196][0] * mat_B[128][0] +
                mat_A[196][1] * mat_B[136][0] +
                mat_A[196][2] * mat_B[144][0] +
                mat_A[196][3] * mat_B[152][0] +
                mat_A[197][0] * mat_B[160][0] +
                mat_A[197][1] * mat_B[168][0] +
                mat_A[197][2] * mat_B[176][0] +
                mat_A[197][3] * mat_B[184][0] +
                mat_A[198][0] * mat_B[192][0] +
                mat_A[198][1] * mat_B[200][0] +
                mat_A[198][2] * mat_B[208][0] +
                mat_A[198][3] * mat_B[216][0] +
                mat_A[199][0] * mat_B[224][0] +
                mat_A[199][1] * mat_B[232][0] +
                mat_A[199][2] * mat_B[240][0] +
                mat_A[199][3] * mat_B[248][0];
    mat_C[192][1] <=
                mat_A[192][0] * mat_B[0][1] +
                mat_A[192][1] * mat_B[8][1] +
                mat_A[192][2] * mat_B[16][1] +
                mat_A[192][3] * mat_B[24][1] +
                mat_A[193][0] * mat_B[32][1] +
                mat_A[193][1] * mat_B[40][1] +
                mat_A[193][2] * mat_B[48][1] +
                mat_A[193][3] * mat_B[56][1] +
                mat_A[194][0] * mat_B[64][1] +
                mat_A[194][1] * mat_B[72][1] +
                mat_A[194][2] * mat_B[80][1] +
                mat_A[194][3] * mat_B[88][1] +
                mat_A[195][0] * mat_B[96][1] +
                mat_A[195][1] * mat_B[104][1] +
                mat_A[195][2] * mat_B[112][1] +
                mat_A[195][3] * mat_B[120][1] +
                mat_A[196][0] * mat_B[128][1] +
                mat_A[196][1] * mat_B[136][1] +
                mat_A[196][2] * mat_B[144][1] +
                mat_A[196][3] * mat_B[152][1] +
                mat_A[197][0] * mat_B[160][1] +
                mat_A[197][1] * mat_B[168][1] +
                mat_A[197][2] * mat_B[176][1] +
                mat_A[197][3] * mat_B[184][1] +
                mat_A[198][0] * mat_B[192][1] +
                mat_A[198][1] * mat_B[200][1] +
                mat_A[198][2] * mat_B[208][1] +
                mat_A[198][3] * mat_B[216][1] +
                mat_A[199][0] * mat_B[224][1] +
                mat_A[199][1] * mat_B[232][1] +
                mat_A[199][2] * mat_B[240][1] +
                mat_A[199][3] * mat_B[248][1];
    mat_C[192][2] <=
                mat_A[192][0] * mat_B[0][2] +
                mat_A[192][1] * mat_B[8][2] +
                mat_A[192][2] * mat_B[16][2] +
                mat_A[192][3] * mat_B[24][2] +
                mat_A[193][0] * mat_B[32][2] +
                mat_A[193][1] * mat_B[40][2] +
                mat_A[193][2] * mat_B[48][2] +
                mat_A[193][3] * mat_B[56][2] +
                mat_A[194][0] * mat_B[64][2] +
                mat_A[194][1] * mat_B[72][2] +
                mat_A[194][2] * mat_B[80][2] +
                mat_A[194][3] * mat_B[88][2] +
                mat_A[195][0] * mat_B[96][2] +
                mat_A[195][1] * mat_B[104][2] +
                mat_A[195][2] * mat_B[112][2] +
                mat_A[195][3] * mat_B[120][2] +
                mat_A[196][0] * mat_B[128][2] +
                mat_A[196][1] * mat_B[136][2] +
                mat_A[196][2] * mat_B[144][2] +
                mat_A[196][3] * mat_B[152][2] +
                mat_A[197][0] * mat_B[160][2] +
                mat_A[197][1] * mat_B[168][2] +
                mat_A[197][2] * mat_B[176][2] +
                mat_A[197][3] * mat_B[184][2] +
                mat_A[198][0] * mat_B[192][2] +
                mat_A[198][1] * mat_B[200][2] +
                mat_A[198][2] * mat_B[208][2] +
                mat_A[198][3] * mat_B[216][2] +
                mat_A[199][0] * mat_B[224][2] +
                mat_A[199][1] * mat_B[232][2] +
                mat_A[199][2] * mat_B[240][2] +
                mat_A[199][3] * mat_B[248][2];
    mat_C[192][3] <=
                mat_A[192][0] * mat_B[0][3] +
                mat_A[192][1] * mat_B[8][3] +
                mat_A[192][2] * mat_B[16][3] +
                mat_A[192][3] * mat_B[24][3] +
                mat_A[193][0] * mat_B[32][3] +
                mat_A[193][1] * mat_B[40][3] +
                mat_A[193][2] * mat_B[48][3] +
                mat_A[193][3] * mat_B[56][3] +
                mat_A[194][0] * mat_B[64][3] +
                mat_A[194][1] * mat_B[72][3] +
                mat_A[194][2] * mat_B[80][3] +
                mat_A[194][3] * mat_B[88][3] +
                mat_A[195][0] * mat_B[96][3] +
                mat_A[195][1] * mat_B[104][3] +
                mat_A[195][2] * mat_B[112][3] +
                mat_A[195][3] * mat_B[120][3] +
                mat_A[196][0] * mat_B[128][3] +
                mat_A[196][1] * mat_B[136][3] +
                mat_A[196][2] * mat_B[144][3] +
                mat_A[196][3] * mat_B[152][3] +
                mat_A[197][0] * mat_B[160][3] +
                mat_A[197][1] * mat_B[168][3] +
                mat_A[197][2] * mat_B[176][3] +
                mat_A[197][3] * mat_B[184][3] +
                mat_A[198][0] * mat_B[192][3] +
                mat_A[198][1] * mat_B[200][3] +
                mat_A[198][2] * mat_B[208][3] +
                mat_A[198][3] * mat_B[216][3] +
                mat_A[199][0] * mat_B[224][3] +
                mat_A[199][1] * mat_B[232][3] +
                mat_A[199][2] * mat_B[240][3] +
                mat_A[199][3] * mat_B[248][3];
    mat_C[193][0] <=
                mat_A[192][0] * mat_B[1][0] +
                mat_A[192][1] * mat_B[9][0] +
                mat_A[192][2] * mat_B[17][0] +
                mat_A[192][3] * mat_B[25][0] +
                mat_A[193][0] * mat_B[33][0] +
                mat_A[193][1] * mat_B[41][0] +
                mat_A[193][2] * mat_B[49][0] +
                mat_A[193][3] * mat_B[57][0] +
                mat_A[194][0] * mat_B[65][0] +
                mat_A[194][1] * mat_B[73][0] +
                mat_A[194][2] * mat_B[81][0] +
                mat_A[194][3] * mat_B[89][0] +
                mat_A[195][0] * mat_B[97][0] +
                mat_A[195][1] * mat_B[105][0] +
                mat_A[195][2] * mat_B[113][0] +
                mat_A[195][3] * mat_B[121][0] +
                mat_A[196][0] * mat_B[129][0] +
                mat_A[196][1] * mat_B[137][0] +
                mat_A[196][2] * mat_B[145][0] +
                mat_A[196][3] * mat_B[153][0] +
                mat_A[197][0] * mat_B[161][0] +
                mat_A[197][1] * mat_B[169][0] +
                mat_A[197][2] * mat_B[177][0] +
                mat_A[197][3] * mat_B[185][0] +
                mat_A[198][0] * mat_B[193][0] +
                mat_A[198][1] * mat_B[201][0] +
                mat_A[198][2] * mat_B[209][0] +
                mat_A[198][3] * mat_B[217][0] +
                mat_A[199][0] * mat_B[225][0] +
                mat_A[199][1] * mat_B[233][0] +
                mat_A[199][2] * mat_B[241][0] +
                mat_A[199][3] * mat_B[249][0];
    mat_C[193][1] <=
                mat_A[192][0] * mat_B[1][1] +
                mat_A[192][1] * mat_B[9][1] +
                mat_A[192][2] * mat_B[17][1] +
                mat_A[192][3] * mat_B[25][1] +
                mat_A[193][0] * mat_B[33][1] +
                mat_A[193][1] * mat_B[41][1] +
                mat_A[193][2] * mat_B[49][1] +
                mat_A[193][3] * mat_B[57][1] +
                mat_A[194][0] * mat_B[65][1] +
                mat_A[194][1] * mat_B[73][1] +
                mat_A[194][2] * mat_B[81][1] +
                mat_A[194][3] * mat_B[89][1] +
                mat_A[195][0] * mat_B[97][1] +
                mat_A[195][1] * mat_B[105][1] +
                mat_A[195][2] * mat_B[113][1] +
                mat_A[195][3] * mat_B[121][1] +
                mat_A[196][0] * mat_B[129][1] +
                mat_A[196][1] * mat_B[137][1] +
                mat_A[196][2] * mat_B[145][1] +
                mat_A[196][3] * mat_B[153][1] +
                mat_A[197][0] * mat_B[161][1] +
                mat_A[197][1] * mat_B[169][1] +
                mat_A[197][2] * mat_B[177][1] +
                mat_A[197][3] * mat_B[185][1] +
                mat_A[198][0] * mat_B[193][1] +
                mat_A[198][1] * mat_B[201][1] +
                mat_A[198][2] * mat_B[209][1] +
                mat_A[198][3] * mat_B[217][1] +
                mat_A[199][0] * mat_B[225][1] +
                mat_A[199][1] * mat_B[233][1] +
                mat_A[199][2] * mat_B[241][1] +
                mat_A[199][3] * mat_B[249][1];
    mat_C[193][2] <=
                mat_A[192][0] * mat_B[1][2] +
                mat_A[192][1] * mat_B[9][2] +
                mat_A[192][2] * mat_B[17][2] +
                mat_A[192][3] * mat_B[25][2] +
                mat_A[193][0] * mat_B[33][2] +
                mat_A[193][1] * mat_B[41][2] +
                mat_A[193][2] * mat_B[49][2] +
                mat_A[193][3] * mat_B[57][2] +
                mat_A[194][0] * mat_B[65][2] +
                mat_A[194][1] * mat_B[73][2] +
                mat_A[194][2] * mat_B[81][2] +
                mat_A[194][3] * mat_B[89][2] +
                mat_A[195][0] * mat_B[97][2] +
                mat_A[195][1] * mat_B[105][2] +
                mat_A[195][2] * mat_B[113][2] +
                mat_A[195][3] * mat_B[121][2] +
                mat_A[196][0] * mat_B[129][2] +
                mat_A[196][1] * mat_B[137][2] +
                mat_A[196][2] * mat_B[145][2] +
                mat_A[196][3] * mat_B[153][2] +
                mat_A[197][0] * mat_B[161][2] +
                mat_A[197][1] * mat_B[169][2] +
                mat_A[197][2] * mat_B[177][2] +
                mat_A[197][3] * mat_B[185][2] +
                mat_A[198][0] * mat_B[193][2] +
                mat_A[198][1] * mat_B[201][2] +
                mat_A[198][2] * mat_B[209][2] +
                mat_A[198][3] * mat_B[217][2] +
                mat_A[199][0] * mat_B[225][2] +
                mat_A[199][1] * mat_B[233][2] +
                mat_A[199][2] * mat_B[241][2] +
                mat_A[199][3] * mat_B[249][2];
    mat_C[193][3] <=
                mat_A[192][0] * mat_B[1][3] +
                mat_A[192][1] * mat_B[9][3] +
                mat_A[192][2] * mat_B[17][3] +
                mat_A[192][3] * mat_B[25][3] +
                mat_A[193][0] * mat_B[33][3] +
                mat_A[193][1] * mat_B[41][3] +
                mat_A[193][2] * mat_B[49][3] +
                mat_A[193][3] * mat_B[57][3] +
                mat_A[194][0] * mat_B[65][3] +
                mat_A[194][1] * mat_B[73][3] +
                mat_A[194][2] * mat_B[81][3] +
                mat_A[194][3] * mat_B[89][3] +
                mat_A[195][0] * mat_B[97][3] +
                mat_A[195][1] * mat_B[105][3] +
                mat_A[195][2] * mat_B[113][3] +
                mat_A[195][3] * mat_B[121][3] +
                mat_A[196][0] * mat_B[129][3] +
                mat_A[196][1] * mat_B[137][3] +
                mat_A[196][2] * mat_B[145][3] +
                mat_A[196][3] * mat_B[153][3] +
                mat_A[197][0] * mat_B[161][3] +
                mat_A[197][1] * mat_B[169][3] +
                mat_A[197][2] * mat_B[177][3] +
                mat_A[197][3] * mat_B[185][3] +
                mat_A[198][0] * mat_B[193][3] +
                mat_A[198][1] * mat_B[201][3] +
                mat_A[198][2] * mat_B[209][3] +
                mat_A[198][3] * mat_B[217][3] +
                mat_A[199][0] * mat_B[225][3] +
                mat_A[199][1] * mat_B[233][3] +
                mat_A[199][2] * mat_B[241][3] +
                mat_A[199][3] * mat_B[249][3];
    mat_C[194][0] <=
                mat_A[192][0] * mat_B[2][0] +
                mat_A[192][1] * mat_B[10][0] +
                mat_A[192][2] * mat_B[18][0] +
                mat_A[192][3] * mat_B[26][0] +
                mat_A[193][0] * mat_B[34][0] +
                mat_A[193][1] * mat_B[42][0] +
                mat_A[193][2] * mat_B[50][0] +
                mat_A[193][3] * mat_B[58][0] +
                mat_A[194][0] * mat_B[66][0] +
                mat_A[194][1] * mat_B[74][0] +
                mat_A[194][2] * mat_B[82][0] +
                mat_A[194][3] * mat_B[90][0] +
                mat_A[195][0] * mat_B[98][0] +
                mat_A[195][1] * mat_B[106][0] +
                mat_A[195][2] * mat_B[114][0] +
                mat_A[195][3] * mat_B[122][0] +
                mat_A[196][0] * mat_B[130][0] +
                mat_A[196][1] * mat_B[138][0] +
                mat_A[196][2] * mat_B[146][0] +
                mat_A[196][3] * mat_B[154][0] +
                mat_A[197][0] * mat_B[162][0] +
                mat_A[197][1] * mat_B[170][0] +
                mat_A[197][2] * mat_B[178][0] +
                mat_A[197][3] * mat_B[186][0] +
                mat_A[198][0] * mat_B[194][0] +
                mat_A[198][1] * mat_B[202][0] +
                mat_A[198][2] * mat_B[210][0] +
                mat_A[198][3] * mat_B[218][0] +
                mat_A[199][0] * mat_B[226][0] +
                mat_A[199][1] * mat_B[234][0] +
                mat_A[199][2] * mat_B[242][0] +
                mat_A[199][3] * mat_B[250][0];
    mat_C[194][1] <=
                mat_A[192][0] * mat_B[2][1] +
                mat_A[192][1] * mat_B[10][1] +
                mat_A[192][2] * mat_B[18][1] +
                mat_A[192][3] * mat_B[26][1] +
                mat_A[193][0] * mat_B[34][1] +
                mat_A[193][1] * mat_B[42][1] +
                mat_A[193][2] * mat_B[50][1] +
                mat_A[193][3] * mat_B[58][1] +
                mat_A[194][0] * mat_B[66][1] +
                mat_A[194][1] * mat_B[74][1] +
                mat_A[194][2] * mat_B[82][1] +
                mat_A[194][3] * mat_B[90][1] +
                mat_A[195][0] * mat_B[98][1] +
                mat_A[195][1] * mat_B[106][1] +
                mat_A[195][2] * mat_B[114][1] +
                mat_A[195][3] * mat_B[122][1] +
                mat_A[196][0] * mat_B[130][1] +
                mat_A[196][1] * mat_B[138][1] +
                mat_A[196][2] * mat_B[146][1] +
                mat_A[196][3] * mat_B[154][1] +
                mat_A[197][0] * mat_B[162][1] +
                mat_A[197][1] * mat_B[170][1] +
                mat_A[197][2] * mat_B[178][1] +
                mat_A[197][3] * mat_B[186][1] +
                mat_A[198][0] * mat_B[194][1] +
                mat_A[198][1] * mat_B[202][1] +
                mat_A[198][2] * mat_B[210][1] +
                mat_A[198][3] * mat_B[218][1] +
                mat_A[199][0] * mat_B[226][1] +
                mat_A[199][1] * mat_B[234][1] +
                mat_A[199][2] * mat_B[242][1] +
                mat_A[199][3] * mat_B[250][1];
    mat_C[194][2] <=
                mat_A[192][0] * mat_B[2][2] +
                mat_A[192][1] * mat_B[10][2] +
                mat_A[192][2] * mat_B[18][2] +
                mat_A[192][3] * mat_B[26][2] +
                mat_A[193][0] * mat_B[34][2] +
                mat_A[193][1] * mat_B[42][2] +
                mat_A[193][2] * mat_B[50][2] +
                mat_A[193][3] * mat_B[58][2] +
                mat_A[194][0] * mat_B[66][2] +
                mat_A[194][1] * mat_B[74][2] +
                mat_A[194][2] * mat_B[82][2] +
                mat_A[194][3] * mat_B[90][2] +
                mat_A[195][0] * mat_B[98][2] +
                mat_A[195][1] * mat_B[106][2] +
                mat_A[195][2] * mat_B[114][2] +
                mat_A[195][3] * mat_B[122][2] +
                mat_A[196][0] * mat_B[130][2] +
                mat_A[196][1] * mat_B[138][2] +
                mat_A[196][2] * mat_B[146][2] +
                mat_A[196][3] * mat_B[154][2] +
                mat_A[197][0] * mat_B[162][2] +
                mat_A[197][1] * mat_B[170][2] +
                mat_A[197][2] * mat_B[178][2] +
                mat_A[197][3] * mat_B[186][2] +
                mat_A[198][0] * mat_B[194][2] +
                mat_A[198][1] * mat_B[202][2] +
                mat_A[198][2] * mat_B[210][2] +
                mat_A[198][3] * mat_B[218][2] +
                mat_A[199][0] * mat_B[226][2] +
                mat_A[199][1] * mat_B[234][2] +
                mat_A[199][2] * mat_B[242][2] +
                mat_A[199][3] * mat_B[250][2];
    mat_C[194][3] <=
                mat_A[192][0] * mat_B[2][3] +
                mat_A[192][1] * mat_B[10][3] +
                mat_A[192][2] * mat_B[18][3] +
                mat_A[192][3] * mat_B[26][3] +
                mat_A[193][0] * mat_B[34][3] +
                mat_A[193][1] * mat_B[42][3] +
                mat_A[193][2] * mat_B[50][3] +
                mat_A[193][3] * mat_B[58][3] +
                mat_A[194][0] * mat_B[66][3] +
                mat_A[194][1] * mat_B[74][3] +
                mat_A[194][2] * mat_B[82][3] +
                mat_A[194][3] * mat_B[90][3] +
                mat_A[195][0] * mat_B[98][3] +
                mat_A[195][1] * mat_B[106][3] +
                mat_A[195][2] * mat_B[114][3] +
                mat_A[195][3] * mat_B[122][3] +
                mat_A[196][0] * mat_B[130][3] +
                mat_A[196][1] * mat_B[138][3] +
                mat_A[196][2] * mat_B[146][3] +
                mat_A[196][3] * mat_B[154][3] +
                mat_A[197][0] * mat_B[162][3] +
                mat_A[197][1] * mat_B[170][3] +
                mat_A[197][2] * mat_B[178][3] +
                mat_A[197][3] * mat_B[186][3] +
                mat_A[198][0] * mat_B[194][3] +
                mat_A[198][1] * mat_B[202][3] +
                mat_A[198][2] * mat_B[210][3] +
                mat_A[198][3] * mat_B[218][3] +
                mat_A[199][0] * mat_B[226][3] +
                mat_A[199][1] * mat_B[234][3] +
                mat_A[199][2] * mat_B[242][3] +
                mat_A[199][3] * mat_B[250][3];
    mat_C[195][0] <=
                mat_A[192][0] * mat_B[3][0] +
                mat_A[192][1] * mat_B[11][0] +
                mat_A[192][2] * mat_B[19][0] +
                mat_A[192][3] * mat_B[27][0] +
                mat_A[193][0] * mat_B[35][0] +
                mat_A[193][1] * mat_B[43][0] +
                mat_A[193][2] * mat_B[51][0] +
                mat_A[193][3] * mat_B[59][0] +
                mat_A[194][0] * mat_B[67][0] +
                mat_A[194][1] * mat_B[75][0] +
                mat_A[194][2] * mat_B[83][0] +
                mat_A[194][3] * mat_B[91][0] +
                mat_A[195][0] * mat_B[99][0] +
                mat_A[195][1] * mat_B[107][0] +
                mat_A[195][2] * mat_B[115][0] +
                mat_A[195][3] * mat_B[123][0] +
                mat_A[196][0] * mat_B[131][0] +
                mat_A[196][1] * mat_B[139][0] +
                mat_A[196][2] * mat_B[147][0] +
                mat_A[196][3] * mat_B[155][0] +
                mat_A[197][0] * mat_B[163][0] +
                mat_A[197][1] * mat_B[171][0] +
                mat_A[197][2] * mat_B[179][0] +
                mat_A[197][3] * mat_B[187][0] +
                mat_A[198][0] * mat_B[195][0] +
                mat_A[198][1] * mat_B[203][0] +
                mat_A[198][2] * mat_B[211][0] +
                mat_A[198][3] * mat_B[219][0] +
                mat_A[199][0] * mat_B[227][0] +
                mat_A[199][1] * mat_B[235][0] +
                mat_A[199][2] * mat_B[243][0] +
                mat_A[199][3] * mat_B[251][0];
    mat_C[195][1] <=
                mat_A[192][0] * mat_B[3][1] +
                mat_A[192][1] * mat_B[11][1] +
                mat_A[192][2] * mat_B[19][1] +
                mat_A[192][3] * mat_B[27][1] +
                mat_A[193][0] * mat_B[35][1] +
                mat_A[193][1] * mat_B[43][1] +
                mat_A[193][2] * mat_B[51][1] +
                mat_A[193][3] * mat_B[59][1] +
                mat_A[194][0] * mat_B[67][1] +
                mat_A[194][1] * mat_B[75][1] +
                mat_A[194][2] * mat_B[83][1] +
                mat_A[194][3] * mat_B[91][1] +
                mat_A[195][0] * mat_B[99][1] +
                mat_A[195][1] * mat_B[107][1] +
                mat_A[195][2] * mat_B[115][1] +
                mat_A[195][3] * mat_B[123][1] +
                mat_A[196][0] * mat_B[131][1] +
                mat_A[196][1] * mat_B[139][1] +
                mat_A[196][2] * mat_B[147][1] +
                mat_A[196][3] * mat_B[155][1] +
                mat_A[197][0] * mat_B[163][1] +
                mat_A[197][1] * mat_B[171][1] +
                mat_A[197][2] * mat_B[179][1] +
                mat_A[197][3] * mat_B[187][1] +
                mat_A[198][0] * mat_B[195][1] +
                mat_A[198][1] * mat_B[203][1] +
                mat_A[198][2] * mat_B[211][1] +
                mat_A[198][3] * mat_B[219][1] +
                mat_A[199][0] * mat_B[227][1] +
                mat_A[199][1] * mat_B[235][1] +
                mat_A[199][2] * mat_B[243][1] +
                mat_A[199][3] * mat_B[251][1];
    mat_C[195][2] <=
                mat_A[192][0] * mat_B[3][2] +
                mat_A[192][1] * mat_B[11][2] +
                mat_A[192][2] * mat_B[19][2] +
                mat_A[192][3] * mat_B[27][2] +
                mat_A[193][0] * mat_B[35][2] +
                mat_A[193][1] * mat_B[43][2] +
                mat_A[193][2] * mat_B[51][2] +
                mat_A[193][3] * mat_B[59][2] +
                mat_A[194][0] * mat_B[67][2] +
                mat_A[194][1] * mat_B[75][2] +
                mat_A[194][2] * mat_B[83][2] +
                mat_A[194][3] * mat_B[91][2] +
                mat_A[195][0] * mat_B[99][2] +
                mat_A[195][1] * mat_B[107][2] +
                mat_A[195][2] * mat_B[115][2] +
                mat_A[195][3] * mat_B[123][2] +
                mat_A[196][0] * mat_B[131][2] +
                mat_A[196][1] * mat_B[139][2] +
                mat_A[196][2] * mat_B[147][2] +
                mat_A[196][3] * mat_B[155][2] +
                mat_A[197][0] * mat_B[163][2] +
                mat_A[197][1] * mat_B[171][2] +
                mat_A[197][2] * mat_B[179][2] +
                mat_A[197][3] * mat_B[187][2] +
                mat_A[198][0] * mat_B[195][2] +
                mat_A[198][1] * mat_B[203][2] +
                mat_A[198][2] * mat_B[211][2] +
                mat_A[198][3] * mat_B[219][2] +
                mat_A[199][0] * mat_B[227][2] +
                mat_A[199][1] * mat_B[235][2] +
                mat_A[199][2] * mat_B[243][2] +
                mat_A[199][3] * mat_B[251][2];
    mat_C[195][3] <=
                mat_A[192][0] * mat_B[3][3] +
                mat_A[192][1] * mat_B[11][3] +
                mat_A[192][2] * mat_B[19][3] +
                mat_A[192][3] * mat_B[27][3] +
                mat_A[193][0] * mat_B[35][3] +
                mat_A[193][1] * mat_B[43][3] +
                mat_A[193][2] * mat_B[51][3] +
                mat_A[193][3] * mat_B[59][3] +
                mat_A[194][0] * mat_B[67][3] +
                mat_A[194][1] * mat_B[75][3] +
                mat_A[194][2] * mat_B[83][3] +
                mat_A[194][3] * mat_B[91][3] +
                mat_A[195][0] * mat_B[99][3] +
                mat_A[195][1] * mat_B[107][3] +
                mat_A[195][2] * mat_B[115][3] +
                mat_A[195][3] * mat_B[123][3] +
                mat_A[196][0] * mat_B[131][3] +
                mat_A[196][1] * mat_B[139][3] +
                mat_A[196][2] * mat_B[147][3] +
                mat_A[196][3] * mat_B[155][3] +
                mat_A[197][0] * mat_B[163][3] +
                mat_A[197][1] * mat_B[171][3] +
                mat_A[197][2] * mat_B[179][3] +
                mat_A[197][3] * mat_B[187][3] +
                mat_A[198][0] * mat_B[195][3] +
                mat_A[198][1] * mat_B[203][3] +
                mat_A[198][2] * mat_B[211][3] +
                mat_A[198][3] * mat_B[219][3] +
                mat_A[199][0] * mat_B[227][3] +
                mat_A[199][1] * mat_B[235][3] +
                mat_A[199][2] * mat_B[243][3] +
                mat_A[199][3] * mat_B[251][3];
    mat_C[196][0] <=
                mat_A[192][0] * mat_B[4][0] +
                mat_A[192][1] * mat_B[12][0] +
                mat_A[192][2] * mat_B[20][0] +
                mat_A[192][3] * mat_B[28][0] +
                mat_A[193][0] * mat_B[36][0] +
                mat_A[193][1] * mat_B[44][0] +
                mat_A[193][2] * mat_B[52][0] +
                mat_A[193][3] * mat_B[60][0] +
                mat_A[194][0] * mat_B[68][0] +
                mat_A[194][1] * mat_B[76][0] +
                mat_A[194][2] * mat_B[84][0] +
                mat_A[194][3] * mat_B[92][0] +
                mat_A[195][0] * mat_B[100][0] +
                mat_A[195][1] * mat_B[108][0] +
                mat_A[195][2] * mat_B[116][0] +
                mat_A[195][3] * mat_B[124][0] +
                mat_A[196][0] * mat_B[132][0] +
                mat_A[196][1] * mat_B[140][0] +
                mat_A[196][2] * mat_B[148][0] +
                mat_A[196][3] * mat_B[156][0] +
                mat_A[197][0] * mat_B[164][0] +
                mat_A[197][1] * mat_B[172][0] +
                mat_A[197][2] * mat_B[180][0] +
                mat_A[197][3] * mat_B[188][0] +
                mat_A[198][0] * mat_B[196][0] +
                mat_A[198][1] * mat_B[204][0] +
                mat_A[198][2] * mat_B[212][0] +
                mat_A[198][3] * mat_B[220][0] +
                mat_A[199][0] * mat_B[228][0] +
                mat_A[199][1] * mat_B[236][0] +
                mat_A[199][2] * mat_B[244][0] +
                mat_A[199][3] * mat_B[252][0];
    mat_C[196][1] <=
                mat_A[192][0] * mat_B[4][1] +
                mat_A[192][1] * mat_B[12][1] +
                mat_A[192][2] * mat_B[20][1] +
                mat_A[192][3] * mat_B[28][1] +
                mat_A[193][0] * mat_B[36][1] +
                mat_A[193][1] * mat_B[44][1] +
                mat_A[193][2] * mat_B[52][1] +
                mat_A[193][3] * mat_B[60][1] +
                mat_A[194][0] * mat_B[68][1] +
                mat_A[194][1] * mat_B[76][1] +
                mat_A[194][2] * mat_B[84][1] +
                mat_A[194][3] * mat_B[92][1] +
                mat_A[195][0] * mat_B[100][1] +
                mat_A[195][1] * mat_B[108][1] +
                mat_A[195][2] * mat_B[116][1] +
                mat_A[195][3] * mat_B[124][1] +
                mat_A[196][0] * mat_B[132][1] +
                mat_A[196][1] * mat_B[140][1] +
                mat_A[196][2] * mat_B[148][1] +
                mat_A[196][3] * mat_B[156][1] +
                mat_A[197][0] * mat_B[164][1] +
                mat_A[197][1] * mat_B[172][1] +
                mat_A[197][2] * mat_B[180][1] +
                mat_A[197][3] * mat_B[188][1] +
                mat_A[198][0] * mat_B[196][1] +
                mat_A[198][1] * mat_B[204][1] +
                mat_A[198][2] * mat_B[212][1] +
                mat_A[198][3] * mat_B[220][1] +
                mat_A[199][0] * mat_B[228][1] +
                mat_A[199][1] * mat_B[236][1] +
                mat_A[199][2] * mat_B[244][1] +
                mat_A[199][3] * mat_B[252][1];
    mat_C[196][2] <=
                mat_A[192][0] * mat_B[4][2] +
                mat_A[192][1] * mat_B[12][2] +
                mat_A[192][2] * mat_B[20][2] +
                mat_A[192][3] * mat_B[28][2] +
                mat_A[193][0] * mat_B[36][2] +
                mat_A[193][1] * mat_B[44][2] +
                mat_A[193][2] * mat_B[52][2] +
                mat_A[193][3] * mat_B[60][2] +
                mat_A[194][0] * mat_B[68][2] +
                mat_A[194][1] * mat_B[76][2] +
                mat_A[194][2] * mat_B[84][2] +
                mat_A[194][3] * mat_B[92][2] +
                mat_A[195][0] * mat_B[100][2] +
                mat_A[195][1] * mat_B[108][2] +
                mat_A[195][2] * mat_B[116][2] +
                mat_A[195][3] * mat_B[124][2] +
                mat_A[196][0] * mat_B[132][2] +
                mat_A[196][1] * mat_B[140][2] +
                mat_A[196][2] * mat_B[148][2] +
                mat_A[196][3] * mat_B[156][2] +
                mat_A[197][0] * mat_B[164][2] +
                mat_A[197][1] * mat_B[172][2] +
                mat_A[197][2] * mat_B[180][2] +
                mat_A[197][3] * mat_B[188][2] +
                mat_A[198][0] * mat_B[196][2] +
                mat_A[198][1] * mat_B[204][2] +
                mat_A[198][2] * mat_B[212][2] +
                mat_A[198][3] * mat_B[220][2] +
                mat_A[199][0] * mat_B[228][2] +
                mat_A[199][1] * mat_B[236][2] +
                mat_A[199][2] * mat_B[244][2] +
                mat_A[199][3] * mat_B[252][2];
    mat_C[196][3] <=
                mat_A[192][0] * mat_B[4][3] +
                mat_A[192][1] * mat_B[12][3] +
                mat_A[192][2] * mat_B[20][3] +
                mat_A[192][3] * mat_B[28][3] +
                mat_A[193][0] * mat_B[36][3] +
                mat_A[193][1] * mat_B[44][3] +
                mat_A[193][2] * mat_B[52][3] +
                mat_A[193][3] * mat_B[60][3] +
                mat_A[194][0] * mat_B[68][3] +
                mat_A[194][1] * mat_B[76][3] +
                mat_A[194][2] * mat_B[84][3] +
                mat_A[194][3] * mat_B[92][3] +
                mat_A[195][0] * mat_B[100][3] +
                mat_A[195][1] * mat_B[108][3] +
                mat_A[195][2] * mat_B[116][3] +
                mat_A[195][3] * mat_B[124][3] +
                mat_A[196][0] * mat_B[132][3] +
                mat_A[196][1] * mat_B[140][3] +
                mat_A[196][2] * mat_B[148][3] +
                mat_A[196][3] * mat_B[156][3] +
                mat_A[197][0] * mat_B[164][3] +
                mat_A[197][1] * mat_B[172][3] +
                mat_A[197][2] * mat_B[180][3] +
                mat_A[197][3] * mat_B[188][3] +
                mat_A[198][0] * mat_B[196][3] +
                mat_A[198][1] * mat_B[204][3] +
                mat_A[198][2] * mat_B[212][3] +
                mat_A[198][3] * mat_B[220][3] +
                mat_A[199][0] * mat_B[228][3] +
                mat_A[199][1] * mat_B[236][3] +
                mat_A[199][2] * mat_B[244][3] +
                mat_A[199][3] * mat_B[252][3];
    mat_C[197][0] <=
                mat_A[192][0] * mat_B[5][0] +
                mat_A[192][1] * mat_B[13][0] +
                mat_A[192][2] * mat_B[21][0] +
                mat_A[192][3] * mat_B[29][0] +
                mat_A[193][0] * mat_B[37][0] +
                mat_A[193][1] * mat_B[45][0] +
                mat_A[193][2] * mat_B[53][0] +
                mat_A[193][3] * mat_B[61][0] +
                mat_A[194][0] * mat_B[69][0] +
                mat_A[194][1] * mat_B[77][0] +
                mat_A[194][2] * mat_B[85][0] +
                mat_A[194][3] * mat_B[93][0] +
                mat_A[195][0] * mat_B[101][0] +
                mat_A[195][1] * mat_B[109][0] +
                mat_A[195][2] * mat_B[117][0] +
                mat_A[195][3] * mat_B[125][0] +
                mat_A[196][0] * mat_B[133][0] +
                mat_A[196][1] * mat_B[141][0] +
                mat_A[196][2] * mat_B[149][0] +
                mat_A[196][3] * mat_B[157][0] +
                mat_A[197][0] * mat_B[165][0] +
                mat_A[197][1] * mat_B[173][0] +
                mat_A[197][2] * mat_B[181][0] +
                mat_A[197][3] * mat_B[189][0] +
                mat_A[198][0] * mat_B[197][0] +
                mat_A[198][1] * mat_B[205][0] +
                mat_A[198][2] * mat_B[213][0] +
                mat_A[198][3] * mat_B[221][0] +
                mat_A[199][0] * mat_B[229][0] +
                mat_A[199][1] * mat_B[237][0] +
                mat_A[199][2] * mat_B[245][0] +
                mat_A[199][3] * mat_B[253][0];
    mat_C[197][1] <=
                mat_A[192][0] * mat_B[5][1] +
                mat_A[192][1] * mat_B[13][1] +
                mat_A[192][2] * mat_B[21][1] +
                mat_A[192][3] * mat_B[29][1] +
                mat_A[193][0] * mat_B[37][1] +
                mat_A[193][1] * mat_B[45][1] +
                mat_A[193][2] * mat_B[53][1] +
                mat_A[193][3] * mat_B[61][1] +
                mat_A[194][0] * mat_B[69][1] +
                mat_A[194][1] * mat_B[77][1] +
                mat_A[194][2] * mat_B[85][1] +
                mat_A[194][3] * mat_B[93][1] +
                mat_A[195][0] * mat_B[101][1] +
                mat_A[195][1] * mat_B[109][1] +
                mat_A[195][2] * mat_B[117][1] +
                mat_A[195][3] * mat_B[125][1] +
                mat_A[196][0] * mat_B[133][1] +
                mat_A[196][1] * mat_B[141][1] +
                mat_A[196][2] * mat_B[149][1] +
                mat_A[196][3] * mat_B[157][1] +
                mat_A[197][0] * mat_B[165][1] +
                mat_A[197][1] * mat_B[173][1] +
                mat_A[197][2] * mat_B[181][1] +
                mat_A[197][3] * mat_B[189][1] +
                mat_A[198][0] * mat_B[197][1] +
                mat_A[198][1] * mat_B[205][1] +
                mat_A[198][2] * mat_B[213][1] +
                mat_A[198][3] * mat_B[221][1] +
                mat_A[199][0] * mat_B[229][1] +
                mat_A[199][1] * mat_B[237][1] +
                mat_A[199][2] * mat_B[245][1] +
                mat_A[199][3] * mat_B[253][1];
    mat_C[197][2] <=
                mat_A[192][0] * mat_B[5][2] +
                mat_A[192][1] * mat_B[13][2] +
                mat_A[192][2] * mat_B[21][2] +
                mat_A[192][3] * mat_B[29][2] +
                mat_A[193][0] * mat_B[37][2] +
                mat_A[193][1] * mat_B[45][2] +
                mat_A[193][2] * mat_B[53][2] +
                mat_A[193][3] * mat_B[61][2] +
                mat_A[194][0] * mat_B[69][2] +
                mat_A[194][1] * mat_B[77][2] +
                mat_A[194][2] * mat_B[85][2] +
                mat_A[194][3] * mat_B[93][2] +
                mat_A[195][0] * mat_B[101][2] +
                mat_A[195][1] * mat_B[109][2] +
                mat_A[195][2] * mat_B[117][2] +
                mat_A[195][3] * mat_B[125][2] +
                mat_A[196][0] * mat_B[133][2] +
                mat_A[196][1] * mat_B[141][2] +
                mat_A[196][2] * mat_B[149][2] +
                mat_A[196][3] * mat_B[157][2] +
                mat_A[197][0] * mat_B[165][2] +
                mat_A[197][1] * mat_B[173][2] +
                mat_A[197][2] * mat_B[181][2] +
                mat_A[197][3] * mat_B[189][2] +
                mat_A[198][0] * mat_B[197][2] +
                mat_A[198][1] * mat_B[205][2] +
                mat_A[198][2] * mat_B[213][2] +
                mat_A[198][3] * mat_B[221][2] +
                mat_A[199][0] * mat_B[229][2] +
                mat_A[199][1] * mat_B[237][2] +
                mat_A[199][2] * mat_B[245][2] +
                mat_A[199][3] * mat_B[253][2];
    mat_C[197][3] <=
                mat_A[192][0] * mat_B[5][3] +
                mat_A[192][1] * mat_B[13][3] +
                mat_A[192][2] * mat_B[21][3] +
                mat_A[192][3] * mat_B[29][3] +
                mat_A[193][0] * mat_B[37][3] +
                mat_A[193][1] * mat_B[45][3] +
                mat_A[193][2] * mat_B[53][3] +
                mat_A[193][3] * mat_B[61][3] +
                mat_A[194][0] * mat_B[69][3] +
                mat_A[194][1] * mat_B[77][3] +
                mat_A[194][2] * mat_B[85][3] +
                mat_A[194][3] * mat_B[93][3] +
                mat_A[195][0] * mat_B[101][3] +
                mat_A[195][1] * mat_B[109][3] +
                mat_A[195][2] * mat_B[117][3] +
                mat_A[195][3] * mat_B[125][3] +
                mat_A[196][0] * mat_B[133][3] +
                mat_A[196][1] * mat_B[141][3] +
                mat_A[196][2] * mat_B[149][3] +
                mat_A[196][3] * mat_B[157][3] +
                mat_A[197][0] * mat_B[165][3] +
                mat_A[197][1] * mat_B[173][3] +
                mat_A[197][2] * mat_B[181][3] +
                mat_A[197][3] * mat_B[189][3] +
                mat_A[198][0] * mat_B[197][3] +
                mat_A[198][1] * mat_B[205][3] +
                mat_A[198][2] * mat_B[213][3] +
                mat_A[198][3] * mat_B[221][3] +
                mat_A[199][0] * mat_B[229][3] +
                mat_A[199][1] * mat_B[237][3] +
                mat_A[199][2] * mat_B[245][3] +
                mat_A[199][3] * mat_B[253][3];
    mat_C[198][0] <=
                mat_A[192][0] * mat_B[6][0] +
                mat_A[192][1] * mat_B[14][0] +
                mat_A[192][2] * mat_B[22][0] +
                mat_A[192][3] * mat_B[30][0] +
                mat_A[193][0] * mat_B[38][0] +
                mat_A[193][1] * mat_B[46][0] +
                mat_A[193][2] * mat_B[54][0] +
                mat_A[193][3] * mat_B[62][0] +
                mat_A[194][0] * mat_B[70][0] +
                mat_A[194][1] * mat_B[78][0] +
                mat_A[194][2] * mat_B[86][0] +
                mat_A[194][3] * mat_B[94][0] +
                mat_A[195][0] * mat_B[102][0] +
                mat_A[195][1] * mat_B[110][0] +
                mat_A[195][2] * mat_B[118][0] +
                mat_A[195][3] * mat_B[126][0] +
                mat_A[196][0] * mat_B[134][0] +
                mat_A[196][1] * mat_B[142][0] +
                mat_A[196][2] * mat_B[150][0] +
                mat_A[196][3] * mat_B[158][0] +
                mat_A[197][0] * mat_B[166][0] +
                mat_A[197][1] * mat_B[174][0] +
                mat_A[197][2] * mat_B[182][0] +
                mat_A[197][3] * mat_B[190][0] +
                mat_A[198][0] * mat_B[198][0] +
                mat_A[198][1] * mat_B[206][0] +
                mat_A[198][2] * mat_B[214][0] +
                mat_A[198][3] * mat_B[222][0] +
                mat_A[199][0] * mat_B[230][0] +
                mat_A[199][1] * mat_B[238][0] +
                mat_A[199][2] * mat_B[246][0] +
                mat_A[199][3] * mat_B[254][0];
    mat_C[198][1] <=
                mat_A[192][0] * mat_B[6][1] +
                mat_A[192][1] * mat_B[14][1] +
                mat_A[192][2] * mat_B[22][1] +
                mat_A[192][3] * mat_B[30][1] +
                mat_A[193][0] * mat_B[38][1] +
                mat_A[193][1] * mat_B[46][1] +
                mat_A[193][2] * mat_B[54][1] +
                mat_A[193][3] * mat_B[62][1] +
                mat_A[194][0] * mat_B[70][1] +
                mat_A[194][1] * mat_B[78][1] +
                mat_A[194][2] * mat_B[86][1] +
                mat_A[194][3] * mat_B[94][1] +
                mat_A[195][0] * mat_B[102][1] +
                mat_A[195][1] * mat_B[110][1] +
                mat_A[195][2] * mat_B[118][1] +
                mat_A[195][3] * mat_B[126][1] +
                mat_A[196][0] * mat_B[134][1] +
                mat_A[196][1] * mat_B[142][1] +
                mat_A[196][2] * mat_B[150][1] +
                mat_A[196][3] * mat_B[158][1] +
                mat_A[197][0] * mat_B[166][1] +
                mat_A[197][1] * mat_B[174][1] +
                mat_A[197][2] * mat_B[182][1] +
                mat_A[197][3] * mat_B[190][1] +
                mat_A[198][0] * mat_B[198][1] +
                mat_A[198][1] * mat_B[206][1] +
                mat_A[198][2] * mat_B[214][1] +
                mat_A[198][3] * mat_B[222][1] +
                mat_A[199][0] * mat_B[230][1] +
                mat_A[199][1] * mat_B[238][1] +
                mat_A[199][2] * mat_B[246][1] +
                mat_A[199][3] * mat_B[254][1];
    mat_C[198][2] <=
                mat_A[192][0] * mat_B[6][2] +
                mat_A[192][1] * mat_B[14][2] +
                mat_A[192][2] * mat_B[22][2] +
                mat_A[192][3] * mat_B[30][2] +
                mat_A[193][0] * mat_B[38][2] +
                mat_A[193][1] * mat_B[46][2] +
                mat_A[193][2] * mat_B[54][2] +
                mat_A[193][3] * mat_B[62][2] +
                mat_A[194][0] * mat_B[70][2] +
                mat_A[194][1] * mat_B[78][2] +
                mat_A[194][2] * mat_B[86][2] +
                mat_A[194][3] * mat_B[94][2] +
                mat_A[195][0] * mat_B[102][2] +
                mat_A[195][1] * mat_B[110][2] +
                mat_A[195][2] * mat_B[118][2] +
                mat_A[195][3] * mat_B[126][2] +
                mat_A[196][0] * mat_B[134][2] +
                mat_A[196][1] * mat_B[142][2] +
                mat_A[196][2] * mat_B[150][2] +
                mat_A[196][3] * mat_B[158][2] +
                mat_A[197][0] * mat_B[166][2] +
                mat_A[197][1] * mat_B[174][2] +
                mat_A[197][2] * mat_B[182][2] +
                mat_A[197][3] * mat_B[190][2] +
                mat_A[198][0] * mat_B[198][2] +
                mat_A[198][1] * mat_B[206][2] +
                mat_A[198][2] * mat_B[214][2] +
                mat_A[198][3] * mat_B[222][2] +
                mat_A[199][0] * mat_B[230][2] +
                mat_A[199][1] * mat_B[238][2] +
                mat_A[199][2] * mat_B[246][2] +
                mat_A[199][3] * mat_B[254][2];
    mat_C[198][3] <=
                mat_A[192][0] * mat_B[6][3] +
                mat_A[192][1] * mat_B[14][3] +
                mat_A[192][2] * mat_B[22][3] +
                mat_A[192][3] * mat_B[30][3] +
                mat_A[193][0] * mat_B[38][3] +
                mat_A[193][1] * mat_B[46][3] +
                mat_A[193][2] * mat_B[54][3] +
                mat_A[193][3] * mat_B[62][3] +
                mat_A[194][0] * mat_B[70][3] +
                mat_A[194][1] * mat_B[78][3] +
                mat_A[194][2] * mat_B[86][3] +
                mat_A[194][3] * mat_B[94][3] +
                mat_A[195][0] * mat_B[102][3] +
                mat_A[195][1] * mat_B[110][3] +
                mat_A[195][2] * mat_B[118][3] +
                mat_A[195][3] * mat_B[126][3] +
                mat_A[196][0] * mat_B[134][3] +
                mat_A[196][1] * mat_B[142][3] +
                mat_A[196][2] * mat_B[150][3] +
                mat_A[196][3] * mat_B[158][3] +
                mat_A[197][0] * mat_B[166][3] +
                mat_A[197][1] * mat_B[174][3] +
                mat_A[197][2] * mat_B[182][3] +
                mat_A[197][3] * mat_B[190][3] +
                mat_A[198][0] * mat_B[198][3] +
                mat_A[198][1] * mat_B[206][3] +
                mat_A[198][2] * mat_B[214][3] +
                mat_A[198][3] * mat_B[222][3] +
                mat_A[199][0] * mat_B[230][3] +
                mat_A[199][1] * mat_B[238][3] +
                mat_A[199][2] * mat_B[246][3] +
                mat_A[199][3] * mat_B[254][3];
    mat_C[199][0] <=
                mat_A[192][0] * mat_B[7][0] +
                mat_A[192][1] * mat_B[15][0] +
                mat_A[192][2] * mat_B[23][0] +
                mat_A[192][3] * mat_B[31][0] +
                mat_A[193][0] * mat_B[39][0] +
                mat_A[193][1] * mat_B[47][0] +
                mat_A[193][2] * mat_B[55][0] +
                mat_A[193][3] * mat_B[63][0] +
                mat_A[194][0] * mat_B[71][0] +
                mat_A[194][1] * mat_B[79][0] +
                mat_A[194][2] * mat_B[87][0] +
                mat_A[194][3] * mat_B[95][0] +
                mat_A[195][0] * mat_B[103][0] +
                mat_A[195][1] * mat_B[111][0] +
                mat_A[195][2] * mat_B[119][0] +
                mat_A[195][3] * mat_B[127][0] +
                mat_A[196][0] * mat_B[135][0] +
                mat_A[196][1] * mat_B[143][0] +
                mat_A[196][2] * mat_B[151][0] +
                mat_A[196][3] * mat_B[159][0] +
                mat_A[197][0] * mat_B[167][0] +
                mat_A[197][1] * mat_B[175][0] +
                mat_A[197][2] * mat_B[183][0] +
                mat_A[197][3] * mat_B[191][0] +
                mat_A[198][0] * mat_B[199][0] +
                mat_A[198][1] * mat_B[207][0] +
                mat_A[198][2] * mat_B[215][0] +
                mat_A[198][3] * mat_B[223][0] +
                mat_A[199][0] * mat_B[231][0] +
                mat_A[199][1] * mat_B[239][0] +
                mat_A[199][2] * mat_B[247][0] +
                mat_A[199][3] * mat_B[255][0];
    mat_C[199][1] <=
                mat_A[192][0] * mat_B[7][1] +
                mat_A[192][1] * mat_B[15][1] +
                mat_A[192][2] * mat_B[23][1] +
                mat_A[192][3] * mat_B[31][1] +
                mat_A[193][0] * mat_B[39][1] +
                mat_A[193][1] * mat_B[47][1] +
                mat_A[193][2] * mat_B[55][1] +
                mat_A[193][3] * mat_B[63][1] +
                mat_A[194][0] * mat_B[71][1] +
                mat_A[194][1] * mat_B[79][1] +
                mat_A[194][2] * mat_B[87][1] +
                mat_A[194][3] * mat_B[95][1] +
                mat_A[195][0] * mat_B[103][1] +
                mat_A[195][1] * mat_B[111][1] +
                mat_A[195][2] * mat_B[119][1] +
                mat_A[195][3] * mat_B[127][1] +
                mat_A[196][0] * mat_B[135][1] +
                mat_A[196][1] * mat_B[143][1] +
                mat_A[196][2] * mat_B[151][1] +
                mat_A[196][3] * mat_B[159][1] +
                mat_A[197][0] * mat_B[167][1] +
                mat_A[197][1] * mat_B[175][1] +
                mat_A[197][2] * mat_B[183][1] +
                mat_A[197][3] * mat_B[191][1] +
                mat_A[198][0] * mat_B[199][1] +
                mat_A[198][1] * mat_B[207][1] +
                mat_A[198][2] * mat_B[215][1] +
                mat_A[198][3] * mat_B[223][1] +
                mat_A[199][0] * mat_B[231][1] +
                mat_A[199][1] * mat_B[239][1] +
                mat_A[199][2] * mat_B[247][1] +
                mat_A[199][3] * mat_B[255][1];
    mat_C[199][2] <=
                mat_A[192][0] * mat_B[7][2] +
                mat_A[192][1] * mat_B[15][2] +
                mat_A[192][2] * mat_B[23][2] +
                mat_A[192][3] * mat_B[31][2] +
                mat_A[193][0] * mat_B[39][2] +
                mat_A[193][1] * mat_B[47][2] +
                mat_A[193][2] * mat_B[55][2] +
                mat_A[193][3] * mat_B[63][2] +
                mat_A[194][0] * mat_B[71][2] +
                mat_A[194][1] * mat_B[79][2] +
                mat_A[194][2] * mat_B[87][2] +
                mat_A[194][3] * mat_B[95][2] +
                mat_A[195][0] * mat_B[103][2] +
                mat_A[195][1] * mat_B[111][2] +
                mat_A[195][2] * mat_B[119][2] +
                mat_A[195][3] * mat_B[127][2] +
                mat_A[196][0] * mat_B[135][2] +
                mat_A[196][1] * mat_B[143][2] +
                mat_A[196][2] * mat_B[151][2] +
                mat_A[196][3] * mat_B[159][2] +
                mat_A[197][0] * mat_B[167][2] +
                mat_A[197][1] * mat_B[175][2] +
                mat_A[197][2] * mat_B[183][2] +
                mat_A[197][3] * mat_B[191][2] +
                mat_A[198][0] * mat_B[199][2] +
                mat_A[198][1] * mat_B[207][2] +
                mat_A[198][2] * mat_B[215][2] +
                mat_A[198][3] * mat_B[223][2] +
                mat_A[199][0] * mat_B[231][2] +
                mat_A[199][1] * mat_B[239][2] +
                mat_A[199][2] * mat_B[247][2] +
                mat_A[199][3] * mat_B[255][2];
    mat_C[199][3] <=
                mat_A[192][0] * mat_B[7][3] +
                mat_A[192][1] * mat_B[15][3] +
                mat_A[192][2] * mat_B[23][3] +
                mat_A[192][3] * mat_B[31][3] +
                mat_A[193][0] * mat_B[39][3] +
                mat_A[193][1] * mat_B[47][3] +
                mat_A[193][2] * mat_B[55][3] +
                mat_A[193][3] * mat_B[63][3] +
                mat_A[194][0] * mat_B[71][3] +
                mat_A[194][1] * mat_B[79][3] +
                mat_A[194][2] * mat_B[87][3] +
                mat_A[194][3] * mat_B[95][3] +
                mat_A[195][0] * mat_B[103][3] +
                mat_A[195][1] * mat_B[111][3] +
                mat_A[195][2] * mat_B[119][3] +
                mat_A[195][3] * mat_B[127][3] +
                mat_A[196][0] * mat_B[135][3] +
                mat_A[196][1] * mat_B[143][3] +
                mat_A[196][2] * mat_B[151][3] +
                mat_A[196][3] * mat_B[159][3] +
                mat_A[197][0] * mat_B[167][3] +
                mat_A[197][1] * mat_B[175][3] +
                mat_A[197][2] * mat_B[183][3] +
                mat_A[197][3] * mat_B[191][3] +
                mat_A[198][0] * mat_B[199][3] +
                mat_A[198][1] * mat_B[207][3] +
                mat_A[198][2] * mat_B[215][3] +
                mat_A[198][3] * mat_B[223][3] +
                mat_A[199][0] * mat_B[231][3] +
                mat_A[199][1] * mat_B[239][3] +
                mat_A[199][2] * mat_B[247][3] +
                mat_A[199][3] * mat_B[255][3];
    mat_C[200][0] <=
                mat_A[200][0] * mat_B[0][0] +
                mat_A[200][1] * mat_B[8][0] +
                mat_A[200][2] * mat_B[16][0] +
                mat_A[200][3] * mat_B[24][0] +
                mat_A[201][0] * mat_B[32][0] +
                mat_A[201][1] * mat_B[40][0] +
                mat_A[201][2] * mat_B[48][0] +
                mat_A[201][3] * mat_B[56][0] +
                mat_A[202][0] * mat_B[64][0] +
                mat_A[202][1] * mat_B[72][0] +
                mat_A[202][2] * mat_B[80][0] +
                mat_A[202][3] * mat_B[88][0] +
                mat_A[203][0] * mat_B[96][0] +
                mat_A[203][1] * mat_B[104][0] +
                mat_A[203][2] * mat_B[112][0] +
                mat_A[203][3] * mat_B[120][0] +
                mat_A[204][0] * mat_B[128][0] +
                mat_A[204][1] * mat_B[136][0] +
                mat_A[204][2] * mat_B[144][0] +
                mat_A[204][3] * mat_B[152][0] +
                mat_A[205][0] * mat_B[160][0] +
                mat_A[205][1] * mat_B[168][0] +
                mat_A[205][2] * mat_B[176][0] +
                mat_A[205][3] * mat_B[184][0] +
                mat_A[206][0] * mat_B[192][0] +
                mat_A[206][1] * mat_B[200][0] +
                mat_A[206][2] * mat_B[208][0] +
                mat_A[206][3] * mat_B[216][0] +
                mat_A[207][0] * mat_B[224][0] +
                mat_A[207][1] * mat_B[232][0] +
                mat_A[207][2] * mat_B[240][0] +
                mat_A[207][3] * mat_B[248][0];
    mat_C[200][1] <=
                mat_A[200][0] * mat_B[0][1] +
                mat_A[200][1] * mat_B[8][1] +
                mat_A[200][2] * mat_B[16][1] +
                mat_A[200][3] * mat_B[24][1] +
                mat_A[201][0] * mat_B[32][1] +
                mat_A[201][1] * mat_B[40][1] +
                mat_A[201][2] * mat_B[48][1] +
                mat_A[201][3] * mat_B[56][1] +
                mat_A[202][0] * mat_B[64][1] +
                mat_A[202][1] * mat_B[72][1] +
                mat_A[202][2] * mat_B[80][1] +
                mat_A[202][3] * mat_B[88][1] +
                mat_A[203][0] * mat_B[96][1] +
                mat_A[203][1] * mat_B[104][1] +
                mat_A[203][2] * mat_B[112][1] +
                mat_A[203][3] * mat_B[120][1] +
                mat_A[204][0] * mat_B[128][1] +
                mat_A[204][1] * mat_B[136][1] +
                mat_A[204][2] * mat_B[144][1] +
                mat_A[204][3] * mat_B[152][1] +
                mat_A[205][0] * mat_B[160][1] +
                mat_A[205][1] * mat_B[168][1] +
                mat_A[205][2] * mat_B[176][1] +
                mat_A[205][3] * mat_B[184][1] +
                mat_A[206][0] * mat_B[192][1] +
                mat_A[206][1] * mat_B[200][1] +
                mat_A[206][2] * mat_B[208][1] +
                mat_A[206][3] * mat_B[216][1] +
                mat_A[207][0] * mat_B[224][1] +
                mat_A[207][1] * mat_B[232][1] +
                mat_A[207][2] * mat_B[240][1] +
                mat_A[207][3] * mat_B[248][1];
    mat_C[200][2] <=
                mat_A[200][0] * mat_B[0][2] +
                mat_A[200][1] * mat_B[8][2] +
                mat_A[200][2] * mat_B[16][2] +
                mat_A[200][3] * mat_B[24][2] +
                mat_A[201][0] * mat_B[32][2] +
                mat_A[201][1] * mat_B[40][2] +
                mat_A[201][2] * mat_B[48][2] +
                mat_A[201][3] * mat_B[56][2] +
                mat_A[202][0] * mat_B[64][2] +
                mat_A[202][1] * mat_B[72][2] +
                mat_A[202][2] * mat_B[80][2] +
                mat_A[202][3] * mat_B[88][2] +
                mat_A[203][0] * mat_B[96][2] +
                mat_A[203][1] * mat_B[104][2] +
                mat_A[203][2] * mat_B[112][2] +
                mat_A[203][3] * mat_B[120][2] +
                mat_A[204][0] * mat_B[128][2] +
                mat_A[204][1] * mat_B[136][2] +
                mat_A[204][2] * mat_B[144][2] +
                mat_A[204][3] * mat_B[152][2] +
                mat_A[205][0] * mat_B[160][2] +
                mat_A[205][1] * mat_B[168][2] +
                mat_A[205][2] * mat_B[176][2] +
                mat_A[205][3] * mat_B[184][2] +
                mat_A[206][0] * mat_B[192][2] +
                mat_A[206][1] * mat_B[200][2] +
                mat_A[206][2] * mat_B[208][2] +
                mat_A[206][3] * mat_B[216][2] +
                mat_A[207][0] * mat_B[224][2] +
                mat_A[207][1] * mat_B[232][2] +
                mat_A[207][2] * mat_B[240][2] +
                mat_A[207][3] * mat_B[248][2];
    mat_C[200][3] <=
                mat_A[200][0] * mat_B[0][3] +
                mat_A[200][1] * mat_B[8][3] +
                mat_A[200][2] * mat_B[16][3] +
                mat_A[200][3] * mat_B[24][3] +
                mat_A[201][0] * mat_B[32][3] +
                mat_A[201][1] * mat_B[40][3] +
                mat_A[201][2] * mat_B[48][3] +
                mat_A[201][3] * mat_B[56][3] +
                mat_A[202][0] * mat_B[64][3] +
                mat_A[202][1] * mat_B[72][3] +
                mat_A[202][2] * mat_B[80][3] +
                mat_A[202][3] * mat_B[88][3] +
                mat_A[203][0] * mat_B[96][3] +
                mat_A[203][1] * mat_B[104][3] +
                mat_A[203][2] * mat_B[112][3] +
                mat_A[203][3] * mat_B[120][3] +
                mat_A[204][0] * mat_B[128][3] +
                mat_A[204][1] * mat_B[136][3] +
                mat_A[204][2] * mat_B[144][3] +
                mat_A[204][3] * mat_B[152][3] +
                mat_A[205][0] * mat_B[160][3] +
                mat_A[205][1] * mat_B[168][3] +
                mat_A[205][2] * mat_B[176][3] +
                mat_A[205][3] * mat_B[184][3] +
                mat_A[206][0] * mat_B[192][3] +
                mat_A[206][1] * mat_B[200][3] +
                mat_A[206][2] * mat_B[208][3] +
                mat_A[206][3] * mat_B[216][3] +
                mat_A[207][0] * mat_B[224][3] +
                mat_A[207][1] * mat_B[232][3] +
                mat_A[207][2] * mat_B[240][3] +
                mat_A[207][3] * mat_B[248][3];
    mat_C[201][0] <=
                mat_A[200][0] * mat_B[1][0] +
                mat_A[200][1] * mat_B[9][0] +
                mat_A[200][2] * mat_B[17][0] +
                mat_A[200][3] * mat_B[25][0] +
                mat_A[201][0] * mat_B[33][0] +
                mat_A[201][1] * mat_B[41][0] +
                mat_A[201][2] * mat_B[49][0] +
                mat_A[201][3] * mat_B[57][0] +
                mat_A[202][0] * mat_B[65][0] +
                mat_A[202][1] * mat_B[73][0] +
                mat_A[202][2] * mat_B[81][0] +
                mat_A[202][3] * mat_B[89][0] +
                mat_A[203][0] * mat_B[97][0] +
                mat_A[203][1] * mat_B[105][0] +
                mat_A[203][2] * mat_B[113][0] +
                mat_A[203][3] * mat_B[121][0] +
                mat_A[204][0] * mat_B[129][0] +
                mat_A[204][1] * mat_B[137][0] +
                mat_A[204][2] * mat_B[145][0] +
                mat_A[204][3] * mat_B[153][0] +
                mat_A[205][0] * mat_B[161][0] +
                mat_A[205][1] * mat_B[169][0] +
                mat_A[205][2] * mat_B[177][0] +
                mat_A[205][3] * mat_B[185][0] +
                mat_A[206][0] * mat_B[193][0] +
                mat_A[206][1] * mat_B[201][0] +
                mat_A[206][2] * mat_B[209][0] +
                mat_A[206][3] * mat_B[217][0] +
                mat_A[207][0] * mat_B[225][0] +
                mat_A[207][1] * mat_B[233][0] +
                mat_A[207][2] * mat_B[241][0] +
                mat_A[207][3] * mat_B[249][0];
    mat_C[201][1] <=
                mat_A[200][0] * mat_B[1][1] +
                mat_A[200][1] * mat_B[9][1] +
                mat_A[200][2] * mat_B[17][1] +
                mat_A[200][3] * mat_B[25][1] +
                mat_A[201][0] * mat_B[33][1] +
                mat_A[201][1] * mat_B[41][1] +
                mat_A[201][2] * mat_B[49][1] +
                mat_A[201][3] * mat_B[57][1] +
                mat_A[202][0] * mat_B[65][1] +
                mat_A[202][1] * mat_B[73][1] +
                mat_A[202][2] * mat_B[81][1] +
                mat_A[202][3] * mat_B[89][1] +
                mat_A[203][0] * mat_B[97][1] +
                mat_A[203][1] * mat_B[105][1] +
                mat_A[203][2] * mat_B[113][1] +
                mat_A[203][3] * mat_B[121][1] +
                mat_A[204][0] * mat_B[129][1] +
                mat_A[204][1] * mat_B[137][1] +
                mat_A[204][2] * mat_B[145][1] +
                mat_A[204][3] * mat_B[153][1] +
                mat_A[205][0] * mat_B[161][1] +
                mat_A[205][1] * mat_B[169][1] +
                mat_A[205][2] * mat_B[177][1] +
                mat_A[205][3] * mat_B[185][1] +
                mat_A[206][0] * mat_B[193][1] +
                mat_A[206][1] * mat_B[201][1] +
                mat_A[206][2] * mat_B[209][1] +
                mat_A[206][3] * mat_B[217][1] +
                mat_A[207][0] * mat_B[225][1] +
                mat_A[207][1] * mat_B[233][1] +
                mat_A[207][2] * mat_B[241][1] +
                mat_A[207][3] * mat_B[249][1];
    mat_C[201][2] <=
                mat_A[200][0] * mat_B[1][2] +
                mat_A[200][1] * mat_B[9][2] +
                mat_A[200][2] * mat_B[17][2] +
                mat_A[200][3] * mat_B[25][2] +
                mat_A[201][0] * mat_B[33][2] +
                mat_A[201][1] * mat_B[41][2] +
                mat_A[201][2] * mat_B[49][2] +
                mat_A[201][3] * mat_B[57][2] +
                mat_A[202][0] * mat_B[65][2] +
                mat_A[202][1] * mat_B[73][2] +
                mat_A[202][2] * mat_B[81][2] +
                mat_A[202][3] * mat_B[89][2] +
                mat_A[203][0] * mat_B[97][2] +
                mat_A[203][1] * mat_B[105][2] +
                mat_A[203][2] * mat_B[113][2] +
                mat_A[203][3] * mat_B[121][2] +
                mat_A[204][0] * mat_B[129][2] +
                mat_A[204][1] * mat_B[137][2] +
                mat_A[204][2] * mat_B[145][2] +
                mat_A[204][3] * mat_B[153][2] +
                mat_A[205][0] * mat_B[161][2] +
                mat_A[205][1] * mat_B[169][2] +
                mat_A[205][2] * mat_B[177][2] +
                mat_A[205][3] * mat_B[185][2] +
                mat_A[206][0] * mat_B[193][2] +
                mat_A[206][1] * mat_B[201][2] +
                mat_A[206][2] * mat_B[209][2] +
                mat_A[206][3] * mat_B[217][2] +
                mat_A[207][0] * mat_B[225][2] +
                mat_A[207][1] * mat_B[233][2] +
                mat_A[207][2] * mat_B[241][2] +
                mat_A[207][3] * mat_B[249][2];
    mat_C[201][3] <=
                mat_A[200][0] * mat_B[1][3] +
                mat_A[200][1] * mat_B[9][3] +
                mat_A[200][2] * mat_B[17][3] +
                mat_A[200][3] * mat_B[25][3] +
                mat_A[201][0] * mat_B[33][3] +
                mat_A[201][1] * mat_B[41][3] +
                mat_A[201][2] * mat_B[49][3] +
                mat_A[201][3] * mat_B[57][3] +
                mat_A[202][0] * mat_B[65][3] +
                mat_A[202][1] * mat_B[73][3] +
                mat_A[202][2] * mat_B[81][3] +
                mat_A[202][3] * mat_B[89][3] +
                mat_A[203][0] * mat_B[97][3] +
                mat_A[203][1] * mat_B[105][3] +
                mat_A[203][2] * mat_B[113][3] +
                mat_A[203][3] * mat_B[121][3] +
                mat_A[204][0] * mat_B[129][3] +
                mat_A[204][1] * mat_B[137][3] +
                mat_A[204][2] * mat_B[145][3] +
                mat_A[204][3] * mat_B[153][3] +
                mat_A[205][0] * mat_B[161][3] +
                mat_A[205][1] * mat_B[169][3] +
                mat_A[205][2] * mat_B[177][3] +
                mat_A[205][3] * mat_B[185][3] +
                mat_A[206][0] * mat_B[193][3] +
                mat_A[206][1] * mat_B[201][3] +
                mat_A[206][2] * mat_B[209][3] +
                mat_A[206][3] * mat_B[217][3] +
                mat_A[207][0] * mat_B[225][3] +
                mat_A[207][1] * mat_B[233][3] +
                mat_A[207][2] * mat_B[241][3] +
                mat_A[207][3] * mat_B[249][3];
    mat_C[202][0] <=
                mat_A[200][0] * mat_B[2][0] +
                mat_A[200][1] * mat_B[10][0] +
                mat_A[200][2] * mat_B[18][0] +
                mat_A[200][3] * mat_B[26][0] +
                mat_A[201][0] * mat_B[34][0] +
                mat_A[201][1] * mat_B[42][0] +
                mat_A[201][2] * mat_B[50][0] +
                mat_A[201][3] * mat_B[58][0] +
                mat_A[202][0] * mat_B[66][0] +
                mat_A[202][1] * mat_B[74][0] +
                mat_A[202][2] * mat_B[82][0] +
                mat_A[202][3] * mat_B[90][0] +
                mat_A[203][0] * mat_B[98][0] +
                mat_A[203][1] * mat_B[106][0] +
                mat_A[203][2] * mat_B[114][0] +
                mat_A[203][3] * mat_B[122][0] +
                mat_A[204][0] * mat_B[130][0] +
                mat_A[204][1] * mat_B[138][0] +
                mat_A[204][2] * mat_B[146][0] +
                mat_A[204][3] * mat_B[154][0] +
                mat_A[205][0] * mat_B[162][0] +
                mat_A[205][1] * mat_B[170][0] +
                mat_A[205][2] * mat_B[178][0] +
                mat_A[205][3] * mat_B[186][0] +
                mat_A[206][0] * mat_B[194][0] +
                mat_A[206][1] * mat_B[202][0] +
                mat_A[206][2] * mat_B[210][0] +
                mat_A[206][3] * mat_B[218][0] +
                mat_A[207][0] * mat_B[226][0] +
                mat_A[207][1] * mat_B[234][0] +
                mat_A[207][2] * mat_B[242][0] +
                mat_A[207][3] * mat_B[250][0];
    mat_C[202][1] <=
                mat_A[200][0] * mat_B[2][1] +
                mat_A[200][1] * mat_B[10][1] +
                mat_A[200][2] * mat_B[18][1] +
                mat_A[200][3] * mat_B[26][1] +
                mat_A[201][0] * mat_B[34][1] +
                mat_A[201][1] * mat_B[42][1] +
                mat_A[201][2] * mat_B[50][1] +
                mat_A[201][3] * mat_B[58][1] +
                mat_A[202][0] * mat_B[66][1] +
                mat_A[202][1] * mat_B[74][1] +
                mat_A[202][2] * mat_B[82][1] +
                mat_A[202][3] * mat_B[90][1] +
                mat_A[203][0] * mat_B[98][1] +
                mat_A[203][1] * mat_B[106][1] +
                mat_A[203][2] * mat_B[114][1] +
                mat_A[203][3] * mat_B[122][1] +
                mat_A[204][0] * mat_B[130][1] +
                mat_A[204][1] * mat_B[138][1] +
                mat_A[204][2] * mat_B[146][1] +
                mat_A[204][3] * mat_B[154][1] +
                mat_A[205][0] * mat_B[162][1] +
                mat_A[205][1] * mat_B[170][1] +
                mat_A[205][2] * mat_B[178][1] +
                mat_A[205][3] * mat_B[186][1] +
                mat_A[206][0] * mat_B[194][1] +
                mat_A[206][1] * mat_B[202][1] +
                mat_A[206][2] * mat_B[210][1] +
                mat_A[206][3] * mat_B[218][1] +
                mat_A[207][0] * mat_B[226][1] +
                mat_A[207][1] * mat_B[234][1] +
                mat_A[207][2] * mat_B[242][1] +
                mat_A[207][3] * mat_B[250][1];
    mat_C[202][2] <=
                mat_A[200][0] * mat_B[2][2] +
                mat_A[200][1] * mat_B[10][2] +
                mat_A[200][2] * mat_B[18][2] +
                mat_A[200][3] * mat_B[26][2] +
                mat_A[201][0] * mat_B[34][2] +
                mat_A[201][1] * mat_B[42][2] +
                mat_A[201][2] * mat_B[50][2] +
                mat_A[201][3] * mat_B[58][2] +
                mat_A[202][0] * mat_B[66][2] +
                mat_A[202][1] * mat_B[74][2] +
                mat_A[202][2] * mat_B[82][2] +
                mat_A[202][3] * mat_B[90][2] +
                mat_A[203][0] * mat_B[98][2] +
                mat_A[203][1] * mat_B[106][2] +
                mat_A[203][2] * mat_B[114][2] +
                mat_A[203][3] * mat_B[122][2] +
                mat_A[204][0] * mat_B[130][2] +
                mat_A[204][1] * mat_B[138][2] +
                mat_A[204][2] * mat_B[146][2] +
                mat_A[204][3] * mat_B[154][2] +
                mat_A[205][0] * mat_B[162][2] +
                mat_A[205][1] * mat_B[170][2] +
                mat_A[205][2] * mat_B[178][2] +
                mat_A[205][3] * mat_B[186][2] +
                mat_A[206][0] * mat_B[194][2] +
                mat_A[206][1] * mat_B[202][2] +
                mat_A[206][2] * mat_B[210][2] +
                mat_A[206][3] * mat_B[218][2] +
                mat_A[207][0] * mat_B[226][2] +
                mat_A[207][1] * mat_B[234][2] +
                mat_A[207][2] * mat_B[242][2] +
                mat_A[207][3] * mat_B[250][2];
    mat_C[202][3] <=
                mat_A[200][0] * mat_B[2][3] +
                mat_A[200][1] * mat_B[10][3] +
                mat_A[200][2] * mat_B[18][3] +
                mat_A[200][3] * mat_B[26][3] +
                mat_A[201][0] * mat_B[34][3] +
                mat_A[201][1] * mat_B[42][3] +
                mat_A[201][2] * mat_B[50][3] +
                mat_A[201][3] * mat_B[58][3] +
                mat_A[202][0] * mat_B[66][3] +
                mat_A[202][1] * mat_B[74][3] +
                mat_A[202][2] * mat_B[82][3] +
                mat_A[202][3] * mat_B[90][3] +
                mat_A[203][0] * mat_B[98][3] +
                mat_A[203][1] * mat_B[106][3] +
                mat_A[203][2] * mat_B[114][3] +
                mat_A[203][3] * mat_B[122][3] +
                mat_A[204][0] * mat_B[130][3] +
                mat_A[204][1] * mat_B[138][3] +
                mat_A[204][2] * mat_B[146][3] +
                mat_A[204][3] * mat_B[154][3] +
                mat_A[205][0] * mat_B[162][3] +
                mat_A[205][1] * mat_B[170][3] +
                mat_A[205][2] * mat_B[178][3] +
                mat_A[205][3] * mat_B[186][3] +
                mat_A[206][0] * mat_B[194][3] +
                mat_A[206][1] * mat_B[202][3] +
                mat_A[206][2] * mat_B[210][3] +
                mat_A[206][3] * mat_B[218][3] +
                mat_A[207][0] * mat_B[226][3] +
                mat_A[207][1] * mat_B[234][3] +
                mat_A[207][2] * mat_B[242][3] +
                mat_A[207][3] * mat_B[250][3];
    mat_C[203][0] <=
                mat_A[200][0] * mat_B[3][0] +
                mat_A[200][1] * mat_B[11][0] +
                mat_A[200][2] * mat_B[19][0] +
                mat_A[200][3] * mat_B[27][0] +
                mat_A[201][0] * mat_B[35][0] +
                mat_A[201][1] * mat_B[43][0] +
                mat_A[201][2] * mat_B[51][0] +
                mat_A[201][3] * mat_B[59][0] +
                mat_A[202][0] * mat_B[67][0] +
                mat_A[202][1] * mat_B[75][0] +
                mat_A[202][2] * mat_B[83][0] +
                mat_A[202][3] * mat_B[91][0] +
                mat_A[203][0] * mat_B[99][0] +
                mat_A[203][1] * mat_B[107][0] +
                mat_A[203][2] * mat_B[115][0] +
                mat_A[203][3] * mat_B[123][0] +
                mat_A[204][0] * mat_B[131][0] +
                mat_A[204][1] * mat_B[139][0] +
                mat_A[204][2] * mat_B[147][0] +
                mat_A[204][3] * mat_B[155][0] +
                mat_A[205][0] * mat_B[163][0] +
                mat_A[205][1] * mat_B[171][0] +
                mat_A[205][2] * mat_B[179][0] +
                mat_A[205][3] * mat_B[187][0] +
                mat_A[206][0] * mat_B[195][0] +
                mat_A[206][1] * mat_B[203][0] +
                mat_A[206][2] * mat_B[211][0] +
                mat_A[206][3] * mat_B[219][0] +
                mat_A[207][0] * mat_B[227][0] +
                mat_A[207][1] * mat_B[235][0] +
                mat_A[207][2] * mat_B[243][0] +
                mat_A[207][3] * mat_B[251][0];
    mat_C[203][1] <=
                mat_A[200][0] * mat_B[3][1] +
                mat_A[200][1] * mat_B[11][1] +
                mat_A[200][2] * mat_B[19][1] +
                mat_A[200][3] * mat_B[27][1] +
                mat_A[201][0] * mat_B[35][1] +
                mat_A[201][1] * mat_B[43][1] +
                mat_A[201][2] * mat_B[51][1] +
                mat_A[201][3] * mat_B[59][1] +
                mat_A[202][0] * mat_B[67][1] +
                mat_A[202][1] * mat_B[75][1] +
                mat_A[202][2] * mat_B[83][1] +
                mat_A[202][3] * mat_B[91][1] +
                mat_A[203][0] * mat_B[99][1] +
                mat_A[203][1] * mat_B[107][1] +
                mat_A[203][2] * mat_B[115][1] +
                mat_A[203][3] * mat_B[123][1] +
                mat_A[204][0] * mat_B[131][1] +
                mat_A[204][1] * mat_B[139][1] +
                mat_A[204][2] * mat_B[147][1] +
                mat_A[204][3] * mat_B[155][1] +
                mat_A[205][0] * mat_B[163][1] +
                mat_A[205][1] * mat_B[171][1] +
                mat_A[205][2] * mat_B[179][1] +
                mat_A[205][3] * mat_B[187][1] +
                mat_A[206][0] * mat_B[195][1] +
                mat_A[206][1] * mat_B[203][1] +
                mat_A[206][2] * mat_B[211][1] +
                mat_A[206][3] * mat_B[219][1] +
                mat_A[207][0] * mat_B[227][1] +
                mat_A[207][1] * mat_B[235][1] +
                mat_A[207][2] * mat_B[243][1] +
                mat_A[207][3] * mat_B[251][1];
    mat_C[203][2] <=
                mat_A[200][0] * mat_B[3][2] +
                mat_A[200][1] * mat_B[11][2] +
                mat_A[200][2] * mat_B[19][2] +
                mat_A[200][3] * mat_B[27][2] +
                mat_A[201][0] * mat_B[35][2] +
                mat_A[201][1] * mat_B[43][2] +
                mat_A[201][2] * mat_B[51][2] +
                mat_A[201][3] * mat_B[59][2] +
                mat_A[202][0] * mat_B[67][2] +
                mat_A[202][1] * mat_B[75][2] +
                mat_A[202][2] * mat_B[83][2] +
                mat_A[202][3] * mat_B[91][2] +
                mat_A[203][0] * mat_B[99][2] +
                mat_A[203][1] * mat_B[107][2] +
                mat_A[203][2] * mat_B[115][2] +
                mat_A[203][3] * mat_B[123][2] +
                mat_A[204][0] * mat_B[131][2] +
                mat_A[204][1] * mat_B[139][2] +
                mat_A[204][2] * mat_B[147][2] +
                mat_A[204][3] * mat_B[155][2] +
                mat_A[205][0] * mat_B[163][2] +
                mat_A[205][1] * mat_B[171][2] +
                mat_A[205][2] * mat_B[179][2] +
                mat_A[205][3] * mat_B[187][2] +
                mat_A[206][0] * mat_B[195][2] +
                mat_A[206][1] * mat_B[203][2] +
                mat_A[206][2] * mat_B[211][2] +
                mat_A[206][3] * mat_B[219][2] +
                mat_A[207][0] * mat_B[227][2] +
                mat_A[207][1] * mat_B[235][2] +
                mat_A[207][2] * mat_B[243][2] +
                mat_A[207][3] * mat_B[251][2];
    mat_C[203][3] <=
                mat_A[200][0] * mat_B[3][3] +
                mat_A[200][1] * mat_B[11][3] +
                mat_A[200][2] * mat_B[19][3] +
                mat_A[200][3] * mat_B[27][3] +
                mat_A[201][0] * mat_B[35][3] +
                mat_A[201][1] * mat_B[43][3] +
                mat_A[201][2] * mat_B[51][3] +
                mat_A[201][3] * mat_B[59][3] +
                mat_A[202][0] * mat_B[67][3] +
                mat_A[202][1] * mat_B[75][3] +
                mat_A[202][2] * mat_B[83][3] +
                mat_A[202][3] * mat_B[91][3] +
                mat_A[203][0] * mat_B[99][3] +
                mat_A[203][1] * mat_B[107][3] +
                mat_A[203][2] * mat_B[115][3] +
                mat_A[203][3] * mat_B[123][3] +
                mat_A[204][0] * mat_B[131][3] +
                mat_A[204][1] * mat_B[139][3] +
                mat_A[204][2] * mat_B[147][3] +
                mat_A[204][3] * mat_B[155][3] +
                mat_A[205][0] * mat_B[163][3] +
                mat_A[205][1] * mat_B[171][3] +
                mat_A[205][2] * mat_B[179][3] +
                mat_A[205][3] * mat_B[187][3] +
                mat_A[206][0] * mat_B[195][3] +
                mat_A[206][1] * mat_B[203][3] +
                mat_A[206][2] * mat_B[211][3] +
                mat_A[206][3] * mat_B[219][3] +
                mat_A[207][0] * mat_B[227][3] +
                mat_A[207][1] * mat_B[235][3] +
                mat_A[207][2] * mat_B[243][3] +
                mat_A[207][3] * mat_B[251][3];
    mat_C[204][0] <=
                mat_A[200][0] * mat_B[4][0] +
                mat_A[200][1] * mat_B[12][0] +
                mat_A[200][2] * mat_B[20][0] +
                mat_A[200][3] * mat_B[28][0] +
                mat_A[201][0] * mat_B[36][0] +
                mat_A[201][1] * mat_B[44][0] +
                mat_A[201][2] * mat_B[52][0] +
                mat_A[201][3] * mat_B[60][0] +
                mat_A[202][0] * mat_B[68][0] +
                mat_A[202][1] * mat_B[76][0] +
                mat_A[202][2] * mat_B[84][0] +
                mat_A[202][3] * mat_B[92][0] +
                mat_A[203][0] * mat_B[100][0] +
                mat_A[203][1] * mat_B[108][0] +
                mat_A[203][2] * mat_B[116][0] +
                mat_A[203][3] * mat_B[124][0] +
                mat_A[204][0] * mat_B[132][0] +
                mat_A[204][1] * mat_B[140][0] +
                mat_A[204][2] * mat_B[148][0] +
                mat_A[204][3] * mat_B[156][0] +
                mat_A[205][0] * mat_B[164][0] +
                mat_A[205][1] * mat_B[172][0] +
                mat_A[205][2] * mat_B[180][0] +
                mat_A[205][3] * mat_B[188][0] +
                mat_A[206][0] * mat_B[196][0] +
                mat_A[206][1] * mat_B[204][0] +
                mat_A[206][2] * mat_B[212][0] +
                mat_A[206][3] * mat_B[220][0] +
                mat_A[207][0] * mat_B[228][0] +
                mat_A[207][1] * mat_B[236][0] +
                mat_A[207][2] * mat_B[244][0] +
                mat_A[207][3] * mat_B[252][0];
    mat_C[204][1] <=
                mat_A[200][0] * mat_B[4][1] +
                mat_A[200][1] * mat_B[12][1] +
                mat_A[200][2] * mat_B[20][1] +
                mat_A[200][3] * mat_B[28][1] +
                mat_A[201][0] * mat_B[36][1] +
                mat_A[201][1] * mat_B[44][1] +
                mat_A[201][2] * mat_B[52][1] +
                mat_A[201][3] * mat_B[60][1] +
                mat_A[202][0] * mat_B[68][1] +
                mat_A[202][1] * mat_B[76][1] +
                mat_A[202][2] * mat_B[84][1] +
                mat_A[202][3] * mat_B[92][1] +
                mat_A[203][0] * mat_B[100][1] +
                mat_A[203][1] * mat_B[108][1] +
                mat_A[203][2] * mat_B[116][1] +
                mat_A[203][3] * mat_B[124][1] +
                mat_A[204][0] * mat_B[132][1] +
                mat_A[204][1] * mat_B[140][1] +
                mat_A[204][2] * mat_B[148][1] +
                mat_A[204][3] * mat_B[156][1] +
                mat_A[205][0] * mat_B[164][1] +
                mat_A[205][1] * mat_B[172][1] +
                mat_A[205][2] * mat_B[180][1] +
                mat_A[205][3] * mat_B[188][1] +
                mat_A[206][0] * mat_B[196][1] +
                mat_A[206][1] * mat_B[204][1] +
                mat_A[206][2] * mat_B[212][1] +
                mat_A[206][3] * mat_B[220][1] +
                mat_A[207][0] * mat_B[228][1] +
                mat_A[207][1] * mat_B[236][1] +
                mat_A[207][2] * mat_B[244][1] +
                mat_A[207][3] * mat_B[252][1];
    mat_C[204][2] <=
                mat_A[200][0] * mat_B[4][2] +
                mat_A[200][1] * mat_B[12][2] +
                mat_A[200][2] * mat_B[20][2] +
                mat_A[200][3] * mat_B[28][2] +
                mat_A[201][0] * mat_B[36][2] +
                mat_A[201][1] * mat_B[44][2] +
                mat_A[201][2] * mat_B[52][2] +
                mat_A[201][3] * mat_B[60][2] +
                mat_A[202][0] * mat_B[68][2] +
                mat_A[202][1] * mat_B[76][2] +
                mat_A[202][2] * mat_B[84][2] +
                mat_A[202][3] * mat_B[92][2] +
                mat_A[203][0] * mat_B[100][2] +
                mat_A[203][1] * mat_B[108][2] +
                mat_A[203][2] * mat_B[116][2] +
                mat_A[203][3] * mat_B[124][2] +
                mat_A[204][0] * mat_B[132][2] +
                mat_A[204][1] * mat_B[140][2] +
                mat_A[204][2] * mat_B[148][2] +
                mat_A[204][3] * mat_B[156][2] +
                mat_A[205][0] * mat_B[164][2] +
                mat_A[205][1] * mat_B[172][2] +
                mat_A[205][2] * mat_B[180][2] +
                mat_A[205][3] * mat_B[188][2] +
                mat_A[206][0] * mat_B[196][2] +
                mat_A[206][1] * mat_B[204][2] +
                mat_A[206][2] * mat_B[212][2] +
                mat_A[206][3] * mat_B[220][2] +
                mat_A[207][0] * mat_B[228][2] +
                mat_A[207][1] * mat_B[236][2] +
                mat_A[207][2] * mat_B[244][2] +
                mat_A[207][3] * mat_B[252][2];
    mat_C[204][3] <=
                mat_A[200][0] * mat_B[4][3] +
                mat_A[200][1] * mat_B[12][3] +
                mat_A[200][2] * mat_B[20][3] +
                mat_A[200][3] * mat_B[28][3] +
                mat_A[201][0] * mat_B[36][3] +
                mat_A[201][1] * mat_B[44][3] +
                mat_A[201][2] * mat_B[52][3] +
                mat_A[201][3] * mat_B[60][3] +
                mat_A[202][0] * mat_B[68][3] +
                mat_A[202][1] * mat_B[76][3] +
                mat_A[202][2] * mat_B[84][3] +
                mat_A[202][3] * mat_B[92][3] +
                mat_A[203][0] * mat_B[100][3] +
                mat_A[203][1] * mat_B[108][3] +
                mat_A[203][2] * mat_B[116][3] +
                mat_A[203][3] * mat_B[124][3] +
                mat_A[204][0] * mat_B[132][3] +
                mat_A[204][1] * mat_B[140][3] +
                mat_A[204][2] * mat_B[148][3] +
                mat_A[204][3] * mat_B[156][3] +
                mat_A[205][0] * mat_B[164][3] +
                mat_A[205][1] * mat_B[172][3] +
                mat_A[205][2] * mat_B[180][3] +
                mat_A[205][3] * mat_B[188][3] +
                mat_A[206][0] * mat_B[196][3] +
                mat_A[206][1] * mat_B[204][3] +
                mat_A[206][2] * mat_B[212][3] +
                mat_A[206][3] * mat_B[220][3] +
                mat_A[207][0] * mat_B[228][3] +
                mat_A[207][1] * mat_B[236][3] +
                mat_A[207][2] * mat_B[244][3] +
                mat_A[207][3] * mat_B[252][3];
    mat_C[205][0] <=
                mat_A[200][0] * mat_B[5][0] +
                mat_A[200][1] * mat_B[13][0] +
                mat_A[200][2] * mat_B[21][0] +
                mat_A[200][3] * mat_B[29][0] +
                mat_A[201][0] * mat_B[37][0] +
                mat_A[201][1] * mat_B[45][0] +
                mat_A[201][2] * mat_B[53][0] +
                mat_A[201][3] * mat_B[61][0] +
                mat_A[202][0] * mat_B[69][0] +
                mat_A[202][1] * mat_B[77][0] +
                mat_A[202][2] * mat_B[85][0] +
                mat_A[202][3] * mat_B[93][0] +
                mat_A[203][0] * mat_B[101][0] +
                mat_A[203][1] * mat_B[109][0] +
                mat_A[203][2] * mat_B[117][0] +
                mat_A[203][3] * mat_B[125][0] +
                mat_A[204][0] * mat_B[133][0] +
                mat_A[204][1] * mat_B[141][0] +
                mat_A[204][2] * mat_B[149][0] +
                mat_A[204][3] * mat_B[157][0] +
                mat_A[205][0] * mat_B[165][0] +
                mat_A[205][1] * mat_B[173][0] +
                mat_A[205][2] * mat_B[181][0] +
                mat_A[205][3] * mat_B[189][0] +
                mat_A[206][0] * mat_B[197][0] +
                mat_A[206][1] * mat_B[205][0] +
                mat_A[206][2] * mat_B[213][0] +
                mat_A[206][3] * mat_B[221][0] +
                mat_A[207][0] * mat_B[229][0] +
                mat_A[207][1] * mat_B[237][0] +
                mat_A[207][2] * mat_B[245][0] +
                mat_A[207][3] * mat_B[253][0];
    mat_C[205][1] <=
                mat_A[200][0] * mat_B[5][1] +
                mat_A[200][1] * mat_B[13][1] +
                mat_A[200][2] * mat_B[21][1] +
                mat_A[200][3] * mat_B[29][1] +
                mat_A[201][0] * mat_B[37][1] +
                mat_A[201][1] * mat_B[45][1] +
                mat_A[201][2] * mat_B[53][1] +
                mat_A[201][3] * mat_B[61][1] +
                mat_A[202][0] * mat_B[69][1] +
                mat_A[202][1] * mat_B[77][1] +
                mat_A[202][2] * mat_B[85][1] +
                mat_A[202][3] * mat_B[93][1] +
                mat_A[203][0] * mat_B[101][1] +
                mat_A[203][1] * mat_B[109][1] +
                mat_A[203][2] * mat_B[117][1] +
                mat_A[203][3] * mat_B[125][1] +
                mat_A[204][0] * mat_B[133][1] +
                mat_A[204][1] * mat_B[141][1] +
                mat_A[204][2] * mat_B[149][1] +
                mat_A[204][3] * mat_B[157][1] +
                mat_A[205][0] * mat_B[165][1] +
                mat_A[205][1] * mat_B[173][1] +
                mat_A[205][2] * mat_B[181][1] +
                mat_A[205][3] * mat_B[189][1] +
                mat_A[206][0] * mat_B[197][1] +
                mat_A[206][1] * mat_B[205][1] +
                mat_A[206][2] * mat_B[213][1] +
                mat_A[206][3] * mat_B[221][1] +
                mat_A[207][0] * mat_B[229][1] +
                mat_A[207][1] * mat_B[237][1] +
                mat_A[207][2] * mat_B[245][1] +
                mat_A[207][3] * mat_B[253][1];
    mat_C[205][2] <=
                mat_A[200][0] * mat_B[5][2] +
                mat_A[200][1] * mat_B[13][2] +
                mat_A[200][2] * mat_B[21][2] +
                mat_A[200][3] * mat_B[29][2] +
                mat_A[201][0] * mat_B[37][2] +
                mat_A[201][1] * mat_B[45][2] +
                mat_A[201][2] * mat_B[53][2] +
                mat_A[201][3] * mat_B[61][2] +
                mat_A[202][0] * mat_B[69][2] +
                mat_A[202][1] * mat_B[77][2] +
                mat_A[202][2] * mat_B[85][2] +
                mat_A[202][3] * mat_B[93][2] +
                mat_A[203][0] * mat_B[101][2] +
                mat_A[203][1] * mat_B[109][2] +
                mat_A[203][2] * mat_B[117][2] +
                mat_A[203][3] * mat_B[125][2] +
                mat_A[204][0] * mat_B[133][2] +
                mat_A[204][1] * mat_B[141][2] +
                mat_A[204][2] * mat_B[149][2] +
                mat_A[204][3] * mat_B[157][2] +
                mat_A[205][0] * mat_B[165][2] +
                mat_A[205][1] * mat_B[173][2] +
                mat_A[205][2] * mat_B[181][2] +
                mat_A[205][3] * mat_B[189][2] +
                mat_A[206][0] * mat_B[197][2] +
                mat_A[206][1] * mat_B[205][2] +
                mat_A[206][2] * mat_B[213][2] +
                mat_A[206][3] * mat_B[221][2] +
                mat_A[207][0] * mat_B[229][2] +
                mat_A[207][1] * mat_B[237][2] +
                mat_A[207][2] * mat_B[245][2] +
                mat_A[207][3] * mat_B[253][2];
    mat_C[205][3] <=
                mat_A[200][0] * mat_B[5][3] +
                mat_A[200][1] * mat_B[13][3] +
                mat_A[200][2] * mat_B[21][3] +
                mat_A[200][3] * mat_B[29][3] +
                mat_A[201][0] * mat_B[37][3] +
                mat_A[201][1] * mat_B[45][3] +
                mat_A[201][2] * mat_B[53][3] +
                mat_A[201][3] * mat_B[61][3] +
                mat_A[202][0] * mat_B[69][3] +
                mat_A[202][1] * mat_B[77][3] +
                mat_A[202][2] * mat_B[85][3] +
                mat_A[202][3] * mat_B[93][3] +
                mat_A[203][0] * mat_B[101][3] +
                mat_A[203][1] * mat_B[109][3] +
                mat_A[203][2] * mat_B[117][3] +
                mat_A[203][3] * mat_B[125][3] +
                mat_A[204][0] * mat_B[133][3] +
                mat_A[204][1] * mat_B[141][3] +
                mat_A[204][2] * mat_B[149][3] +
                mat_A[204][3] * mat_B[157][3] +
                mat_A[205][0] * mat_B[165][3] +
                mat_A[205][1] * mat_B[173][3] +
                mat_A[205][2] * mat_B[181][3] +
                mat_A[205][3] * mat_B[189][3] +
                mat_A[206][0] * mat_B[197][3] +
                mat_A[206][1] * mat_B[205][3] +
                mat_A[206][2] * mat_B[213][3] +
                mat_A[206][3] * mat_B[221][3] +
                mat_A[207][0] * mat_B[229][3] +
                mat_A[207][1] * mat_B[237][3] +
                mat_A[207][2] * mat_B[245][3] +
                mat_A[207][3] * mat_B[253][3];
    mat_C[206][0] <=
                mat_A[200][0] * mat_B[6][0] +
                mat_A[200][1] * mat_B[14][0] +
                mat_A[200][2] * mat_B[22][0] +
                mat_A[200][3] * mat_B[30][0] +
                mat_A[201][0] * mat_B[38][0] +
                mat_A[201][1] * mat_B[46][0] +
                mat_A[201][2] * mat_B[54][0] +
                mat_A[201][3] * mat_B[62][0] +
                mat_A[202][0] * mat_B[70][0] +
                mat_A[202][1] * mat_B[78][0] +
                mat_A[202][2] * mat_B[86][0] +
                mat_A[202][3] * mat_B[94][0] +
                mat_A[203][0] * mat_B[102][0] +
                mat_A[203][1] * mat_B[110][0] +
                mat_A[203][2] * mat_B[118][0] +
                mat_A[203][3] * mat_B[126][0] +
                mat_A[204][0] * mat_B[134][0] +
                mat_A[204][1] * mat_B[142][0] +
                mat_A[204][2] * mat_B[150][0] +
                mat_A[204][3] * mat_B[158][0] +
                mat_A[205][0] * mat_B[166][0] +
                mat_A[205][1] * mat_B[174][0] +
                mat_A[205][2] * mat_B[182][0] +
                mat_A[205][3] * mat_B[190][0] +
                mat_A[206][0] * mat_B[198][0] +
                mat_A[206][1] * mat_B[206][0] +
                mat_A[206][2] * mat_B[214][0] +
                mat_A[206][3] * mat_B[222][0] +
                mat_A[207][0] * mat_B[230][0] +
                mat_A[207][1] * mat_B[238][0] +
                mat_A[207][2] * mat_B[246][0] +
                mat_A[207][3] * mat_B[254][0];
    mat_C[206][1] <=
                mat_A[200][0] * mat_B[6][1] +
                mat_A[200][1] * mat_B[14][1] +
                mat_A[200][2] * mat_B[22][1] +
                mat_A[200][3] * mat_B[30][1] +
                mat_A[201][0] * mat_B[38][1] +
                mat_A[201][1] * mat_B[46][1] +
                mat_A[201][2] * mat_B[54][1] +
                mat_A[201][3] * mat_B[62][1] +
                mat_A[202][0] * mat_B[70][1] +
                mat_A[202][1] * mat_B[78][1] +
                mat_A[202][2] * mat_B[86][1] +
                mat_A[202][3] * mat_B[94][1] +
                mat_A[203][0] * mat_B[102][1] +
                mat_A[203][1] * mat_B[110][1] +
                mat_A[203][2] * mat_B[118][1] +
                mat_A[203][3] * mat_B[126][1] +
                mat_A[204][0] * mat_B[134][1] +
                mat_A[204][1] * mat_B[142][1] +
                mat_A[204][2] * mat_B[150][1] +
                mat_A[204][3] * mat_B[158][1] +
                mat_A[205][0] * mat_B[166][1] +
                mat_A[205][1] * mat_B[174][1] +
                mat_A[205][2] * mat_B[182][1] +
                mat_A[205][3] * mat_B[190][1] +
                mat_A[206][0] * mat_B[198][1] +
                mat_A[206][1] * mat_B[206][1] +
                mat_A[206][2] * mat_B[214][1] +
                mat_A[206][3] * mat_B[222][1] +
                mat_A[207][0] * mat_B[230][1] +
                mat_A[207][1] * mat_B[238][1] +
                mat_A[207][2] * mat_B[246][1] +
                mat_A[207][3] * mat_B[254][1];
    mat_C[206][2] <=
                mat_A[200][0] * mat_B[6][2] +
                mat_A[200][1] * mat_B[14][2] +
                mat_A[200][2] * mat_B[22][2] +
                mat_A[200][3] * mat_B[30][2] +
                mat_A[201][0] * mat_B[38][2] +
                mat_A[201][1] * mat_B[46][2] +
                mat_A[201][2] * mat_B[54][2] +
                mat_A[201][3] * mat_B[62][2] +
                mat_A[202][0] * mat_B[70][2] +
                mat_A[202][1] * mat_B[78][2] +
                mat_A[202][2] * mat_B[86][2] +
                mat_A[202][3] * mat_B[94][2] +
                mat_A[203][0] * mat_B[102][2] +
                mat_A[203][1] * mat_B[110][2] +
                mat_A[203][2] * mat_B[118][2] +
                mat_A[203][3] * mat_B[126][2] +
                mat_A[204][0] * mat_B[134][2] +
                mat_A[204][1] * mat_B[142][2] +
                mat_A[204][2] * mat_B[150][2] +
                mat_A[204][3] * mat_B[158][2] +
                mat_A[205][0] * mat_B[166][2] +
                mat_A[205][1] * mat_B[174][2] +
                mat_A[205][2] * mat_B[182][2] +
                mat_A[205][3] * mat_B[190][2] +
                mat_A[206][0] * mat_B[198][2] +
                mat_A[206][1] * mat_B[206][2] +
                mat_A[206][2] * mat_B[214][2] +
                mat_A[206][3] * mat_B[222][2] +
                mat_A[207][0] * mat_B[230][2] +
                mat_A[207][1] * mat_B[238][2] +
                mat_A[207][2] * mat_B[246][2] +
                mat_A[207][3] * mat_B[254][2];
    mat_C[206][3] <=
                mat_A[200][0] * mat_B[6][3] +
                mat_A[200][1] * mat_B[14][3] +
                mat_A[200][2] * mat_B[22][3] +
                mat_A[200][3] * mat_B[30][3] +
                mat_A[201][0] * mat_B[38][3] +
                mat_A[201][1] * mat_B[46][3] +
                mat_A[201][2] * mat_B[54][3] +
                mat_A[201][3] * mat_B[62][3] +
                mat_A[202][0] * mat_B[70][3] +
                mat_A[202][1] * mat_B[78][3] +
                mat_A[202][2] * mat_B[86][3] +
                mat_A[202][3] * mat_B[94][3] +
                mat_A[203][0] * mat_B[102][3] +
                mat_A[203][1] * mat_B[110][3] +
                mat_A[203][2] * mat_B[118][3] +
                mat_A[203][3] * mat_B[126][3] +
                mat_A[204][0] * mat_B[134][3] +
                mat_A[204][1] * mat_B[142][3] +
                mat_A[204][2] * mat_B[150][3] +
                mat_A[204][3] * mat_B[158][3] +
                mat_A[205][0] * mat_B[166][3] +
                mat_A[205][1] * mat_B[174][3] +
                mat_A[205][2] * mat_B[182][3] +
                mat_A[205][3] * mat_B[190][3] +
                mat_A[206][0] * mat_B[198][3] +
                mat_A[206][1] * mat_B[206][3] +
                mat_A[206][2] * mat_B[214][3] +
                mat_A[206][3] * mat_B[222][3] +
                mat_A[207][0] * mat_B[230][3] +
                mat_A[207][1] * mat_B[238][3] +
                mat_A[207][2] * mat_B[246][3] +
                mat_A[207][3] * mat_B[254][3];
    mat_C[207][0] <=
                mat_A[200][0] * mat_B[7][0] +
                mat_A[200][1] * mat_B[15][0] +
                mat_A[200][2] * mat_B[23][0] +
                mat_A[200][3] * mat_B[31][0] +
                mat_A[201][0] * mat_B[39][0] +
                mat_A[201][1] * mat_B[47][0] +
                mat_A[201][2] * mat_B[55][0] +
                mat_A[201][3] * mat_B[63][0] +
                mat_A[202][0] * mat_B[71][0] +
                mat_A[202][1] * mat_B[79][0] +
                mat_A[202][2] * mat_B[87][0] +
                mat_A[202][3] * mat_B[95][0] +
                mat_A[203][0] * mat_B[103][0] +
                mat_A[203][1] * mat_B[111][0] +
                mat_A[203][2] * mat_B[119][0] +
                mat_A[203][3] * mat_B[127][0] +
                mat_A[204][0] * mat_B[135][0] +
                mat_A[204][1] * mat_B[143][0] +
                mat_A[204][2] * mat_B[151][0] +
                mat_A[204][3] * mat_B[159][0] +
                mat_A[205][0] * mat_B[167][0] +
                mat_A[205][1] * mat_B[175][0] +
                mat_A[205][2] * mat_B[183][0] +
                mat_A[205][3] * mat_B[191][0] +
                mat_A[206][0] * mat_B[199][0] +
                mat_A[206][1] * mat_B[207][0] +
                mat_A[206][2] * mat_B[215][0] +
                mat_A[206][3] * mat_B[223][0] +
                mat_A[207][0] * mat_B[231][0] +
                mat_A[207][1] * mat_B[239][0] +
                mat_A[207][2] * mat_B[247][0] +
                mat_A[207][3] * mat_B[255][0];
    mat_C[207][1] <=
                mat_A[200][0] * mat_B[7][1] +
                mat_A[200][1] * mat_B[15][1] +
                mat_A[200][2] * mat_B[23][1] +
                mat_A[200][3] * mat_B[31][1] +
                mat_A[201][0] * mat_B[39][1] +
                mat_A[201][1] * mat_B[47][1] +
                mat_A[201][2] * mat_B[55][1] +
                mat_A[201][3] * mat_B[63][1] +
                mat_A[202][0] * mat_B[71][1] +
                mat_A[202][1] * mat_B[79][1] +
                mat_A[202][2] * mat_B[87][1] +
                mat_A[202][3] * mat_B[95][1] +
                mat_A[203][0] * mat_B[103][1] +
                mat_A[203][1] * mat_B[111][1] +
                mat_A[203][2] * mat_B[119][1] +
                mat_A[203][3] * mat_B[127][1] +
                mat_A[204][0] * mat_B[135][1] +
                mat_A[204][1] * mat_B[143][1] +
                mat_A[204][2] * mat_B[151][1] +
                mat_A[204][3] * mat_B[159][1] +
                mat_A[205][0] * mat_B[167][1] +
                mat_A[205][1] * mat_B[175][1] +
                mat_A[205][2] * mat_B[183][1] +
                mat_A[205][3] * mat_B[191][1] +
                mat_A[206][0] * mat_B[199][1] +
                mat_A[206][1] * mat_B[207][1] +
                mat_A[206][2] * mat_B[215][1] +
                mat_A[206][3] * mat_B[223][1] +
                mat_A[207][0] * mat_B[231][1] +
                mat_A[207][1] * mat_B[239][1] +
                mat_A[207][2] * mat_B[247][1] +
                mat_A[207][3] * mat_B[255][1];
    mat_C[207][2] <=
                mat_A[200][0] * mat_B[7][2] +
                mat_A[200][1] * mat_B[15][2] +
                mat_A[200][2] * mat_B[23][2] +
                mat_A[200][3] * mat_B[31][2] +
                mat_A[201][0] * mat_B[39][2] +
                mat_A[201][1] * mat_B[47][2] +
                mat_A[201][2] * mat_B[55][2] +
                mat_A[201][3] * mat_B[63][2] +
                mat_A[202][0] * mat_B[71][2] +
                mat_A[202][1] * mat_B[79][2] +
                mat_A[202][2] * mat_B[87][2] +
                mat_A[202][3] * mat_B[95][2] +
                mat_A[203][0] * mat_B[103][2] +
                mat_A[203][1] * mat_B[111][2] +
                mat_A[203][2] * mat_B[119][2] +
                mat_A[203][3] * mat_B[127][2] +
                mat_A[204][0] * mat_B[135][2] +
                mat_A[204][1] * mat_B[143][2] +
                mat_A[204][2] * mat_B[151][2] +
                mat_A[204][3] * mat_B[159][2] +
                mat_A[205][0] * mat_B[167][2] +
                mat_A[205][1] * mat_B[175][2] +
                mat_A[205][2] * mat_B[183][2] +
                mat_A[205][3] * mat_B[191][2] +
                mat_A[206][0] * mat_B[199][2] +
                mat_A[206][1] * mat_B[207][2] +
                mat_A[206][2] * mat_B[215][2] +
                mat_A[206][3] * mat_B[223][2] +
                mat_A[207][0] * mat_B[231][2] +
                mat_A[207][1] * mat_B[239][2] +
                mat_A[207][2] * mat_B[247][2] +
                mat_A[207][3] * mat_B[255][2];
    mat_C[207][3] <=
                mat_A[200][0] * mat_B[7][3] +
                mat_A[200][1] * mat_B[15][3] +
                mat_A[200][2] * mat_B[23][3] +
                mat_A[200][3] * mat_B[31][3] +
                mat_A[201][0] * mat_B[39][3] +
                mat_A[201][1] * mat_B[47][3] +
                mat_A[201][2] * mat_B[55][3] +
                mat_A[201][3] * mat_B[63][3] +
                mat_A[202][0] * mat_B[71][3] +
                mat_A[202][1] * mat_B[79][3] +
                mat_A[202][2] * mat_B[87][3] +
                mat_A[202][3] * mat_B[95][3] +
                mat_A[203][0] * mat_B[103][3] +
                mat_A[203][1] * mat_B[111][3] +
                mat_A[203][2] * mat_B[119][3] +
                mat_A[203][3] * mat_B[127][3] +
                mat_A[204][0] * mat_B[135][3] +
                mat_A[204][1] * mat_B[143][3] +
                mat_A[204][2] * mat_B[151][3] +
                mat_A[204][3] * mat_B[159][3] +
                mat_A[205][0] * mat_B[167][3] +
                mat_A[205][1] * mat_B[175][3] +
                mat_A[205][2] * mat_B[183][3] +
                mat_A[205][3] * mat_B[191][3] +
                mat_A[206][0] * mat_B[199][3] +
                mat_A[206][1] * mat_B[207][3] +
                mat_A[206][2] * mat_B[215][3] +
                mat_A[206][3] * mat_B[223][3] +
                mat_A[207][0] * mat_B[231][3] +
                mat_A[207][1] * mat_B[239][3] +
                mat_A[207][2] * mat_B[247][3] +
                mat_A[207][3] * mat_B[255][3];
    mat_C[208][0] <=
                mat_A[208][0] * mat_B[0][0] +
                mat_A[208][1] * mat_B[8][0] +
                mat_A[208][2] * mat_B[16][0] +
                mat_A[208][3] * mat_B[24][0] +
                mat_A[209][0] * mat_B[32][0] +
                mat_A[209][1] * mat_B[40][0] +
                mat_A[209][2] * mat_B[48][0] +
                mat_A[209][3] * mat_B[56][0] +
                mat_A[210][0] * mat_B[64][0] +
                mat_A[210][1] * mat_B[72][0] +
                mat_A[210][2] * mat_B[80][0] +
                mat_A[210][3] * mat_B[88][0] +
                mat_A[211][0] * mat_B[96][0] +
                mat_A[211][1] * mat_B[104][0] +
                mat_A[211][2] * mat_B[112][0] +
                mat_A[211][3] * mat_B[120][0] +
                mat_A[212][0] * mat_B[128][0] +
                mat_A[212][1] * mat_B[136][0] +
                mat_A[212][2] * mat_B[144][0] +
                mat_A[212][3] * mat_B[152][0] +
                mat_A[213][0] * mat_B[160][0] +
                mat_A[213][1] * mat_B[168][0] +
                mat_A[213][2] * mat_B[176][0] +
                mat_A[213][3] * mat_B[184][0] +
                mat_A[214][0] * mat_B[192][0] +
                mat_A[214][1] * mat_B[200][0] +
                mat_A[214][2] * mat_B[208][0] +
                mat_A[214][3] * mat_B[216][0] +
                mat_A[215][0] * mat_B[224][0] +
                mat_A[215][1] * mat_B[232][0] +
                mat_A[215][2] * mat_B[240][0] +
                mat_A[215][3] * mat_B[248][0];
    mat_C[208][1] <=
                mat_A[208][0] * mat_B[0][1] +
                mat_A[208][1] * mat_B[8][1] +
                mat_A[208][2] * mat_B[16][1] +
                mat_A[208][3] * mat_B[24][1] +
                mat_A[209][0] * mat_B[32][1] +
                mat_A[209][1] * mat_B[40][1] +
                mat_A[209][2] * mat_B[48][1] +
                mat_A[209][3] * mat_B[56][1] +
                mat_A[210][0] * mat_B[64][1] +
                mat_A[210][1] * mat_B[72][1] +
                mat_A[210][2] * mat_B[80][1] +
                mat_A[210][3] * mat_B[88][1] +
                mat_A[211][0] * mat_B[96][1] +
                mat_A[211][1] * mat_B[104][1] +
                mat_A[211][2] * mat_B[112][1] +
                mat_A[211][3] * mat_B[120][1] +
                mat_A[212][0] * mat_B[128][1] +
                mat_A[212][1] * mat_B[136][1] +
                mat_A[212][2] * mat_B[144][1] +
                mat_A[212][3] * mat_B[152][1] +
                mat_A[213][0] * mat_B[160][1] +
                mat_A[213][1] * mat_B[168][1] +
                mat_A[213][2] * mat_B[176][1] +
                mat_A[213][3] * mat_B[184][1] +
                mat_A[214][0] * mat_B[192][1] +
                mat_A[214][1] * mat_B[200][1] +
                mat_A[214][2] * mat_B[208][1] +
                mat_A[214][3] * mat_B[216][1] +
                mat_A[215][0] * mat_B[224][1] +
                mat_A[215][1] * mat_B[232][1] +
                mat_A[215][2] * mat_B[240][1] +
                mat_A[215][3] * mat_B[248][1];
    mat_C[208][2] <=
                mat_A[208][0] * mat_B[0][2] +
                mat_A[208][1] * mat_B[8][2] +
                mat_A[208][2] * mat_B[16][2] +
                mat_A[208][3] * mat_B[24][2] +
                mat_A[209][0] * mat_B[32][2] +
                mat_A[209][1] * mat_B[40][2] +
                mat_A[209][2] * mat_B[48][2] +
                mat_A[209][3] * mat_B[56][2] +
                mat_A[210][0] * mat_B[64][2] +
                mat_A[210][1] * mat_B[72][2] +
                mat_A[210][2] * mat_B[80][2] +
                mat_A[210][3] * mat_B[88][2] +
                mat_A[211][0] * mat_B[96][2] +
                mat_A[211][1] * mat_B[104][2] +
                mat_A[211][2] * mat_B[112][2] +
                mat_A[211][3] * mat_B[120][2] +
                mat_A[212][0] * mat_B[128][2] +
                mat_A[212][1] * mat_B[136][2] +
                mat_A[212][2] * mat_B[144][2] +
                mat_A[212][3] * mat_B[152][2] +
                mat_A[213][0] * mat_B[160][2] +
                mat_A[213][1] * mat_B[168][2] +
                mat_A[213][2] * mat_B[176][2] +
                mat_A[213][3] * mat_B[184][2] +
                mat_A[214][0] * mat_B[192][2] +
                mat_A[214][1] * mat_B[200][2] +
                mat_A[214][2] * mat_B[208][2] +
                mat_A[214][3] * mat_B[216][2] +
                mat_A[215][0] * mat_B[224][2] +
                mat_A[215][1] * mat_B[232][2] +
                mat_A[215][2] * mat_B[240][2] +
                mat_A[215][3] * mat_B[248][2];
    mat_C[208][3] <=
                mat_A[208][0] * mat_B[0][3] +
                mat_A[208][1] * mat_B[8][3] +
                mat_A[208][2] * mat_B[16][3] +
                mat_A[208][3] * mat_B[24][3] +
                mat_A[209][0] * mat_B[32][3] +
                mat_A[209][1] * mat_B[40][3] +
                mat_A[209][2] * mat_B[48][3] +
                mat_A[209][3] * mat_B[56][3] +
                mat_A[210][0] * mat_B[64][3] +
                mat_A[210][1] * mat_B[72][3] +
                mat_A[210][2] * mat_B[80][3] +
                mat_A[210][3] * mat_B[88][3] +
                mat_A[211][0] * mat_B[96][3] +
                mat_A[211][1] * mat_B[104][3] +
                mat_A[211][2] * mat_B[112][3] +
                mat_A[211][3] * mat_B[120][3] +
                mat_A[212][0] * mat_B[128][3] +
                mat_A[212][1] * mat_B[136][3] +
                mat_A[212][2] * mat_B[144][3] +
                mat_A[212][3] * mat_B[152][3] +
                mat_A[213][0] * mat_B[160][3] +
                mat_A[213][1] * mat_B[168][3] +
                mat_A[213][2] * mat_B[176][3] +
                mat_A[213][3] * mat_B[184][3] +
                mat_A[214][0] * mat_B[192][3] +
                mat_A[214][1] * mat_B[200][3] +
                mat_A[214][2] * mat_B[208][3] +
                mat_A[214][3] * mat_B[216][3] +
                mat_A[215][0] * mat_B[224][3] +
                mat_A[215][1] * mat_B[232][3] +
                mat_A[215][2] * mat_B[240][3] +
                mat_A[215][3] * mat_B[248][3];
    mat_C[209][0] <=
                mat_A[208][0] * mat_B[1][0] +
                mat_A[208][1] * mat_B[9][0] +
                mat_A[208][2] * mat_B[17][0] +
                mat_A[208][3] * mat_B[25][0] +
                mat_A[209][0] * mat_B[33][0] +
                mat_A[209][1] * mat_B[41][0] +
                mat_A[209][2] * mat_B[49][0] +
                mat_A[209][3] * mat_B[57][0] +
                mat_A[210][0] * mat_B[65][0] +
                mat_A[210][1] * mat_B[73][0] +
                mat_A[210][2] * mat_B[81][0] +
                mat_A[210][3] * mat_B[89][0] +
                mat_A[211][0] * mat_B[97][0] +
                mat_A[211][1] * mat_B[105][0] +
                mat_A[211][2] * mat_B[113][0] +
                mat_A[211][3] * mat_B[121][0] +
                mat_A[212][0] * mat_B[129][0] +
                mat_A[212][1] * mat_B[137][0] +
                mat_A[212][2] * mat_B[145][0] +
                mat_A[212][3] * mat_B[153][0] +
                mat_A[213][0] * mat_B[161][0] +
                mat_A[213][1] * mat_B[169][0] +
                mat_A[213][2] * mat_B[177][0] +
                mat_A[213][3] * mat_B[185][0] +
                mat_A[214][0] * mat_B[193][0] +
                mat_A[214][1] * mat_B[201][0] +
                mat_A[214][2] * mat_B[209][0] +
                mat_A[214][3] * mat_B[217][0] +
                mat_A[215][0] * mat_B[225][0] +
                mat_A[215][1] * mat_B[233][0] +
                mat_A[215][2] * mat_B[241][0] +
                mat_A[215][3] * mat_B[249][0];
    mat_C[209][1] <=
                mat_A[208][0] * mat_B[1][1] +
                mat_A[208][1] * mat_B[9][1] +
                mat_A[208][2] * mat_B[17][1] +
                mat_A[208][3] * mat_B[25][1] +
                mat_A[209][0] * mat_B[33][1] +
                mat_A[209][1] * mat_B[41][1] +
                mat_A[209][2] * mat_B[49][1] +
                mat_A[209][3] * mat_B[57][1] +
                mat_A[210][0] * mat_B[65][1] +
                mat_A[210][1] * mat_B[73][1] +
                mat_A[210][2] * mat_B[81][1] +
                mat_A[210][3] * mat_B[89][1] +
                mat_A[211][0] * mat_B[97][1] +
                mat_A[211][1] * mat_B[105][1] +
                mat_A[211][2] * mat_B[113][1] +
                mat_A[211][3] * mat_B[121][1] +
                mat_A[212][0] * mat_B[129][1] +
                mat_A[212][1] * mat_B[137][1] +
                mat_A[212][2] * mat_B[145][1] +
                mat_A[212][3] * mat_B[153][1] +
                mat_A[213][0] * mat_B[161][1] +
                mat_A[213][1] * mat_B[169][1] +
                mat_A[213][2] * mat_B[177][1] +
                mat_A[213][3] * mat_B[185][1] +
                mat_A[214][0] * mat_B[193][1] +
                mat_A[214][1] * mat_B[201][1] +
                mat_A[214][2] * mat_B[209][1] +
                mat_A[214][3] * mat_B[217][1] +
                mat_A[215][0] * mat_B[225][1] +
                mat_A[215][1] * mat_B[233][1] +
                mat_A[215][2] * mat_B[241][1] +
                mat_A[215][3] * mat_B[249][1];
    mat_C[209][2] <=
                mat_A[208][0] * mat_B[1][2] +
                mat_A[208][1] * mat_B[9][2] +
                mat_A[208][2] * mat_B[17][2] +
                mat_A[208][3] * mat_B[25][2] +
                mat_A[209][0] * mat_B[33][2] +
                mat_A[209][1] * mat_B[41][2] +
                mat_A[209][2] * mat_B[49][2] +
                mat_A[209][3] * mat_B[57][2] +
                mat_A[210][0] * mat_B[65][2] +
                mat_A[210][1] * mat_B[73][2] +
                mat_A[210][2] * mat_B[81][2] +
                mat_A[210][3] * mat_B[89][2] +
                mat_A[211][0] * mat_B[97][2] +
                mat_A[211][1] * mat_B[105][2] +
                mat_A[211][2] * mat_B[113][2] +
                mat_A[211][3] * mat_B[121][2] +
                mat_A[212][0] * mat_B[129][2] +
                mat_A[212][1] * mat_B[137][2] +
                mat_A[212][2] * mat_B[145][2] +
                mat_A[212][3] * mat_B[153][2] +
                mat_A[213][0] * mat_B[161][2] +
                mat_A[213][1] * mat_B[169][2] +
                mat_A[213][2] * mat_B[177][2] +
                mat_A[213][3] * mat_B[185][2] +
                mat_A[214][0] * mat_B[193][2] +
                mat_A[214][1] * mat_B[201][2] +
                mat_A[214][2] * mat_B[209][2] +
                mat_A[214][3] * mat_B[217][2] +
                mat_A[215][0] * mat_B[225][2] +
                mat_A[215][1] * mat_B[233][2] +
                mat_A[215][2] * mat_B[241][2] +
                mat_A[215][3] * mat_B[249][2];
    mat_C[209][3] <=
                mat_A[208][0] * mat_B[1][3] +
                mat_A[208][1] * mat_B[9][3] +
                mat_A[208][2] * mat_B[17][3] +
                mat_A[208][3] * mat_B[25][3] +
                mat_A[209][0] * mat_B[33][3] +
                mat_A[209][1] * mat_B[41][3] +
                mat_A[209][2] * mat_B[49][3] +
                mat_A[209][3] * mat_B[57][3] +
                mat_A[210][0] * mat_B[65][3] +
                mat_A[210][1] * mat_B[73][3] +
                mat_A[210][2] * mat_B[81][3] +
                mat_A[210][3] * mat_B[89][3] +
                mat_A[211][0] * mat_B[97][3] +
                mat_A[211][1] * mat_B[105][3] +
                mat_A[211][2] * mat_B[113][3] +
                mat_A[211][3] * mat_B[121][3] +
                mat_A[212][0] * mat_B[129][3] +
                mat_A[212][1] * mat_B[137][3] +
                mat_A[212][2] * mat_B[145][3] +
                mat_A[212][3] * mat_B[153][3] +
                mat_A[213][0] * mat_B[161][3] +
                mat_A[213][1] * mat_B[169][3] +
                mat_A[213][2] * mat_B[177][3] +
                mat_A[213][3] * mat_B[185][3] +
                mat_A[214][0] * mat_B[193][3] +
                mat_A[214][1] * mat_B[201][3] +
                mat_A[214][2] * mat_B[209][3] +
                mat_A[214][3] * mat_B[217][3] +
                mat_A[215][0] * mat_B[225][3] +
                mat_A[215][1] * mat_B[233][3] +
                mat_A[215][2] * mat_B[241][3] +
                mat_A[215][3] * mat_B[249][3];
    mat_C[210][0] <=
                mat_A[208][0] * mat_B[2][0] +
                mat_A[208][1] * mat_B[10][0] +
                mat_A[208][2] * mat_B[18][0] +
                mat_A[208][3] * mat_B[26][0] +
                mat_A[209][0] * mat_B[34][0] +
                mat_A[209][1] * mat_B[42][0] +
                mat_A[209][2] * mat_B[50][0] +
                mat_A[209][3] * mat_B[58][0] +
                mat_A[210][0] * mat_B[66][0] +
                mat_A[210][1] * mat_B[74][0] +
                mat_A[210][2] * mat_B[82][0] +
                mat_A[210][3] * mat_B[90][0] +
                mat_A[211][0] * mat_B[98][0] +
                mat_A[211][1] * mat_B[106][0] +
                mat_A[211][2] * mat_B[114][0] +
                mat_A[211][3] * mat_B[122][0] +
                mat_A[212][0] * mat_B[130][0] +
                mat_A[212][1] * mat_B[138][0] +
                mat_A[212][2] * mat_B[146][0] +
                mat_A[212][3] * mat_B[154][0] +
                mat_A[213][0] * mat_B[162][0] +
                mat_A[213][1] * mat_B[170][0] +
                mat_A[213][2] * mat_B[178][0] +
                mat_A[213][3] * mat_B[186][0] +
                mat_A[214][0] * mat_B[194][0] +
                mat_A[214][1] * mat_B[202][0] +
                mat_A[214][2] * mat_B[210][0] +
                mat_A[214][3] * mat_B[218][0] +
                mat_A[215][0] * mat_B[226][0] +
                mat_A[215][1] * mat_B[234][0] +
                mat_A[215][2] * mat_B[242][0] +
                mat_A[215][3] * mat_B[250][0];
    mat_C[210][1] <=
                mat_A[208][0] * mat_B[2][1] +
                mat_A[208][1] * mat_B[10][1] +
                mat_A[208][2] * mat_B[18][1] +
                mat_A[208][3] * mat_B[26][1] +
                mat_A[209][0] * mat_B[34][1] +
                mat_A[209][1] * mat_B[42][1] +
                mat_A[209][2] * mat_B[50][1] +
                mat_A[209][3] * mat_B[58][1] +
                mat_A[210][0] * mat_B[66][1] +
                mat_A[210][1] * mat_B[74][1] +
                mat_A[210][2] * mat_B[82][1] +
                mat_A[210][3] * mat_B[90][1] +
                mat_A[211][0] * mat_B[98][1] +
                mat_A[211][1] * mat_B[106][1] +
                mat_A[211][2] * mat_B[114][1] +
                mat_A[211][3] * mat_B[122][1] +
                mat_A[212][0] * mat_B[130][1] +
                mat_A[212][1] * mat_B[138][1] +
                mat_A[212][2] * mat_B[146][1] +
                mat_A[212][3] * mat_B[154][1] +
                mat_A[213][0] * mat_B[162][1] +
                mat_A[213][1] * mat_B[170][1] +
                mat_A[213][2] * mat_B[178][1] +
                mat_A[213][3] * mat_B[186][1] +
                mat_A[214][0] * mat_B[194][1] +
                mat_A[214][1] * mat_B[202][1] +
                mat_A[214][2] * mat_B[210][1] +
                mat_A[214][3] * mat_B[218][1] +
                mat_A[215][0] * mat_B[226][1] +
                mat_A[215][1] * mat_B[234][1] +
                mat_A[215][2] * mat_B[242][1] +
                mat_A[215][3] * mat_B[250][1];
    mat_C[210][2] <=
                mat_A[208][0] * mat_B[2][2] +
                mat_A[208][1] * mat_B[10][2] +
                mat_A[208][2] * mat_B[18][2] +
                mat_A[208][3] * mat_B[26][2] +
                mat_A[209][0] * mat_B[34][2] +
                mat_A[209][1] * mat_B[42][2] +
                mat_A[209][2] * mat_B[50][2] +
                mat_A[209][3] * mat_B[58][2] +
                mat_A[210][0] * mat_B[66][2] +
                mat_A[210][1] * mat_B[74][2] +
                mat_A[210][2] * mat_B[82][2] +
                mat_A[210][3] * mat_B[90][2] +
                mat_A[211][0] * mat_B[98][2] +
                mat_A[211][1] * mat_B[106][2] +
                mat_A[211][2] * mat_B[114][2] +
                mat_A[211][3] * mat_B[122][2] +
                mat_A[212][0] * mat_B[130][2] +
                mat_A[212][1] * mat_B[138][2] +
                mat_A[212][2] * mat_B[146][2] +
                mat_A[212][3] * mat_B[154][2] +
                mat_A[213][0] * mat_B[162][2] +
                mat_A[213][1] * mat_B[170][2] +
                mat_A[213][2] * mat_B[178][2] +
                mat_A[213][3] * mat_B[186][2] +
                mat_A[214][0] * mat_B[194][2] +
                mat_A[214][1] * mat_B[202][2] +
                mat_A[214][2] * mat_B[210][2] +
                mat_A[214][3] * mat_B[218][2] +
                mat_A[215][0] * mat_B[226][2] +
                mat_A[215][1] * mat_B[234][2] +
                mat_A[215][2] * mat_B[242][2] +
                mat_A[215][3] * mat_B[250][2];
    mat_C[210][3] <=
                mat_A[208][0] * mat_B[2][3] +
                mat_A[208][1] * mat_B[10][3] +
                mat_A[208][2] * mat_B[18][3] +
                mat_A[208][3] * mat_B[26][3] +
                mat_A[209][0] * mat_B[34][3] +
                mat_A[209][1] * mat_B[42][3] +
                mat_A[209][2] * mat_B[50][3] +
                mat_A[209][3] * mat_B[58][3] +
                mat_A[210][0] * mat_B[66][3] +
                mat_A[210][1] * mat_B[74][3] +
                mat_A[210][2] * mat_B[82][3] +
                mat_A[210][3] * mat_B[90][3] +
                mat_A[211][0] * mat_B[98][3] +
                mat_A[211][1] * mat_B[106][3] +
                mat_A[211][2] * mat_B[114][3] +
                mat_A[211][3] * mat_B[122][3] +
                mat_A[212][0] * mat_B[130][3] +
                mat_A[212][1] * mat_B[138][3] +
                mat_A[212][2] * mat_B[146][3] +
                mat_A[212][3] * mat_B[154][3] +
                mat_A[213][0] * mat_B[162][3] +
                mat_A[213][1] * mat_B[170][3] +
                mat_A[213][2] * mat_B[178][3] +
                mat_A[213][3] * mat_B[186][3] +
                mat_A[214][0] * mat_B[194][3] +
                mat_A[214][1] * mat_B[202][3] +
                mat_A[214][2] * mat_B[210][3] +
                mat_A[214][3] * mat_B[218][3] +
                mat_A[215][0] * mat_B[226][3] +
                mat_A[215][1] * mat_B[234][3] +
                mat_A[215][2] * mat_B[242][3] +
                mat_A[215][3] * mat_B[250][3];
    mat_C[211][0] <=
                mat_A[208][0] * mat_B[3][0] +
                mat_A[208][1] * mat_B[11][0] +
                mat_A[208][2] * mat_B[19][0] +
                mat_A[208][3] * mat_B[27][0] +
                mat_A[209][0] * mat_B[35][0] +
                mat_A[209][1] * mat_B[43][0] +
                mat_A[209][2] * mat_B[51][0] +
                mat_A[209][3] * mat_B[59][0] +
                mat_A[210][0] * mat_B[67][0] +
                mat_A[210][1] * mat_B[75][0] +
                mat_A[210][2] * mat_B[83][0] +
                mat_A[210][3] * mat_B[91][0] +
                mat_A[211][0] * mat_B[99][0] +
                mat_A[211][1] * mat_B[107][0] +
                mat_A[211][2] * mat_B[115][0] +
                mat_A[211][3] * mat_B[123][0] +
                mat_A[212][0] * mat_B[131][0] +
                mat_A[212][1] * mat_B[139][0] +
                mat_A[212][2] * mat_B[147][0] +
                mat_A[212][3] * mat_B[155][0] +
                mat_A[213][0] * mat_B[163][0] +
                mat_A[213][1] * mat_B[171][0] +
                mat_A[213][2] * mat_B[179][0] +
                mat_A[213][3] * mat_B[187][0] +
                mat_A[214][0] * mat_B[195][0] +
                mat_A[214][1] * mat_B[203][0] +
                mat_A[214][2] * mat_B[211][0] +
                mat_A[214][3] * mat_B[219][0] +
                mat_A[215][0] * mat_B[227][0] +
                mat_A[215][1] * mat_B[235][0] +
                mat_A[215][2] * mat_B[243][0] +
                mat_A[215][3] * mat_B[251][0];
    mat_C[211][1] <=
                mat_A[208][0] * mat_B[3][1] +
                mat_A[208][1] * mat_B[11][1] +
                mat_A[208][2] * mat_B[19][1] +
                mat_A[208][3] * mat_B[27][1] +
                mat_A[209][0] * mat_B[35][1] +
                mat_A[209][1] * mat_B[43][1] +
                mat_A[209][2] * mat_B[51][1] +
                mat_A[209][3] * mat_B[59][1] +
                mat_A[210][0] * mat_B[67][1] +
                mat_A[210][1] * mat_B[75][1] +
                mat_A[210][2] * mat_B[83][1] +
                mat_A[210][3] * mat_B[91][1] +
                mat_A[211][0] * mat_B[99][1] +
                mat_A[211][1] * mat_B[107][1] +
                mat_A[211][2] * mat_B[115][1] +
                mat_A[211][3] * mat_B[123][1] +
                mat_A[212][0] * mat_B[131][1] +
                mat_A[212][1] * mat_B[139][1] +
                mat_A[212][2] * mat_B[147][1] +
                mat_A[212][3] * mat_B[155][1] +
                mat_A[213][0] * mat_B[163][1] +
                mat_A[213][1] * mat_B[171][1] +
                mat_A[213][2] * mat_B[179][1] +
                mat_A[213][3] * mat_B[187][1] +
                mat_A[214][0] * mat_B[195][1] +
                mat_A[214][1] * mat_B[203][1] +
                mat_A[214][2] * mat_B[211][1] +
                mat_A[214][3] * mat_B[219][1] +
                mat_A[215][0] * mat_B[227][1] +
                mat_A[215][1] * mat_B[235][1] +
                mat_A[215][2] * mat_B[243][1] +
                mat_A[215][3] * mat_B[251][1];
    mat_C[211][2] <=
                mat_A[208][0] * mat_B[3][2] +
                mat_A[208][1] * mat_B[11][2] +
                mat_A[208][2] * mat_B[19][2] +
                mat_A[208][3] * mat_B[27][2] +
                mat_A[209][0] * mat_B[35][2] +
                mat_A[209][1] * mat_B[43][2] +
                mat_A[209][2] * mat_B[51][2] +
                mat_A[209][3] * mat_B[59][2] +
                mat_A[210][0] * mat_B[67][2] +
                mat_A[210][1] * mat_B[75][2] +
                mat_A[210][2] * mat_B[83][2] +
                mat_A[210][3] * mat_B[91][2] +
                mat_A[211][0] * mat_B[99][2] +
                mat_A[211][1] * mat_B[107][2] +
                mat_A[211][2] * mat_B[115][2] +
                mat_A[211][3] * mat_B[123][2] +
                mat_A[212][0] * mat_B[131][2] +
                mat_A[212][1] * mat_B[139][2] +
                mat_A[212][2] * mat_B[147][2] +
                mat_A[212][3] * mat_B[155][2] +
                mat_A[213][0] * mat_B[163][2] +
                mat_A[213][1] * mat_B[171][2] +
                mat_A[213][2] * mat_B[179][2] +
                mat_A[213][3] * mat_B[187][2] +
                mat_A[214][0] * mat_B[195][2] +
                mat_A[214][1] * mat_B[203][2] +
                mat_A[214][2] * mat_B[211][2] +
                mat_A[214][3] * mat_B[219][2] +
                mat_A[215][0] * mat_B[227][2] +
                mat_A[215][1] * mat_B[235][2] +
                mat_A[215][2] * mat_B[243][2] +
                mat_A[215][3] * mat_B[251][2];
    mat_C[211][3] <=
                mat_A[208][0] * mat_B[3][3] +
                mat_A[208][1] * mat_B[11][3] +
                mat_A[208][2] * mat_B[19][3] +
                mat_A[208][3] * mat_B[27][3] +
                mat_A[209][0] * mat_B[35][3] +
                mat_A[209][1] * mat_B[43][3] +
                mat_A[209][2] * mat_B[51][3] +
                mat_A[209][3] * mat_B[59][3] +
                mat_A[210][0] * mat_B[67][3] +
                mat_A[210][1] * mat_B[75][3] +
                mat_A[210][2] * mat_B[83][3] +
                mat_A[210][3] * mat_B[91][3] +
                mat_A[211][0] * mat_B[99][3] +
                mat_A[211][1] * mat_B[107][3] +
                mat_A[211][2] * mat_B[115][3] +
                mat_A[211][3] * mat_B[123][3] +
                mat_A[212][0] * mat_B[131][3] +
                mat_A[212][1] * mat_B[139][3] +
                mat_A[212][2] * mat_B[147][3] +
                mat_A[212][3] * mat_B[155][3] +
                mat_A[213][0] * mat_B[163][3] +
                mat_A[213][1] * mat_B[171][3] +
                mat_A[213][2] * mat_B[179][3] +
                mat_A[213][3] * mat_B[187][3] +
                mat_A[214][0] * mat_B[195][3] +
                mat_A[214][1] * mat_B[203][3] +
                mat_A[214][2] * mat_B[211][3] +
                mat_A[214][3] * mat_B[219][3] +
                mat_A[215][0] * mat_B[227][3] +
                mat_A[215][1] * mat_B[235][3] +
                mat_A[215][2] * mat_B[243][3] +
                mat_A[215][3] * mat_B[251][3];
    mat_C[212][0] <=
                mat_A[208][0] * mat_B[4][0] +
                mat_A[208][1] * mat_B[12][0] +
                mat_A[208][2] * mat_B[20][0] +
                mat_A[208][3] * mat_B[28][0] +
                mat_A[209][0] * mat_B[36][0] +
                mat_A[209][1] * mat_B[44][0] +
                mat_A[209][2] * mat_B[52][0] +
                mat_A[209][3] * mat_B[60][0] +
                mat_A[210][0] * mat_B[68][0] +
                mat_A[210][1] * mat_B[76][0] +
                mat_A[210][2] * mat_B[84][0] +
                mat_A[210][3] * mat_B[92][0] +
                mat_A[211][0] * mat_B[100][0] +
                mat_A[211][1] * mat_B[108][0] +
                mat_A[211][2] * mat_B[116][0] +
                mat_A[211][3] * mat_B[124][0] +
                mat_A[212][0] * mat_B[132][0] +
                mat_A[212][1] * mat_B[140][0] +
                mat_A[212][2] * mat_B[148][0] +
                mat_A[212][3] * mat_B[156][0] +
                mat_A[213][0] * mat_B[164][0] +
                mat_A[213][1] * mat_B[172][0] +
                mat_A[213][2] * mat_B[180][0] +
                mat_A[213][3] * mat_B[188][0] +
                mat_A[214][0] * mat_B[196][0] +
                mat_A[214][1] * mat_B[204][0] +
                mat_A[214][2] * mat_B[212][0] +
                mat_A[214][3] * mat_B[220][0] +
                mat_A[215][0] * mat_B[228][0] +
                mat_A[215][1] * mat_B[236][0] +
                mat_A[215][2] * mat_B[244][0] +
                mat_A[215][3] * mat_B[252][0];
    mat_C[212][1] <=
                mat_A[208][0] * mat_B[4][1] +
                mat_A[208][1] * mat_B[12][1] +
                mat_A[208][2] * mat_B[20][1] +
                mat_A[208][3] * mat_B[28][1] +
                mat_A[209][0] * mat_B[36][1] +
                mat_A[209][1] * mat_B[44][1] +
                mat_A[209][2] * mat_B[52][1] +
                mat_A[209][3] * mat_B[60][1] +
                mat_A[210][0] * mat_B[68][1] +
                mat_A[210][1] * mat_B[76][1] +
                mat_A[210][2] * mat_B[84][1] +
                mat_A[210][3] * mat_B[92][1] +
                mat_A[211][0] * mat_B[100][1] +
                mat_A[211][1] * mat_B[108][1] +
                mat_A[211][2] * mat_B[116][1] +
                mat_A[211][3] * mat_B[124][1] +
                mat_A[212][0] * mat_B[132][1] +
                mat_A[212][1] * mat_B[140][1] +
                mat_A[212][2] * mat_B[148][1] +
                mat_A[212][3] * mat_B[156][1] +
                mat_A[213][0] * mat_B[164][1] +
                mat_A[213][1] * mat_B[172][1] +
                mat_A[213][2] * mat_B[180][1] +
                mat_A[213][3] * mat_B[188][1] +
                mat_A[214][0] * mat_B[196][1] +
                mat_A[214][1] * mat_B[204][1] +
                mat_A[214][2] * mat_B[212][1] +
                mat_A[214][3] * mat_B[220][1] +
                mat_A[215][0] * mat_B[228][1] +
                mat_A[215][1] * mat_B[236][1] +
                mat_A[215][2] * mat_B[244][1] +
                mat_A[215][3] * mat_B[252][1];
    mat_C[212][2] <=
                mat_A[208][0] * mat_B[4][2] +
                mat_A[208][1] * mat_B[12][2] +
                mat_A[208][2] * mat_B[20][2] +
                mat_A[208][3] * mat_B[28][2] +
                mat_A[209][0] * mat_B[36][2] +
                mat_A[209][1] * mat_B[44][2] +
                mat_A[209][2] * mat_B[52][2] +
                mat_A[209][3] * mat_B[60][2] +
                mat_A[210][0] * mat_B[68][2] +
                mat_A[210][1] * mat_B[76][2] +
                mat_A[210][2] * mat_B[84][2] +
                mat_A[210][3] * mat_B[92][2] +
                mat_A[211][0] * mat_B[100][2] +
                mat_A[211][1] * mat_B[108][2] +
                mat_A[211][2] * mat_B[116][2] +
                mat_A[211][3] * mat_B[124][2] +
                mat_A[212][0] * mat_B[132][2] +
                mat_A[212][1] * mat_B[140][2] +
                mat_A[212][2] * mat_B[148][2] +
                mat_A[212][3] * mat_B[156][2] +
                mat_A[213][0] * mat_B[164][2] +
                mat_A[213][1] * mat_B[172][2] +
                mat_A[213][2] * mat_B[180][2] +
                mat_A[213][3] * mat_B[188][2] +
                mat_A[214][0] * mat_B[196][2] +
                mat_A[214][1] * mat_B[204][2] +
                mat_A[214][2] * mat_B[212][2] +
                mat_A[214][3] * mat_B[220][2] +
                mat_A[215][0] * mat_B[228][2] +
                mat_A[215][1] * mat_B[236][2] +
                mat_A[215][2] * mat_B[244][2] +
                mat_A[215][3] * mat_B[252][2];
    mat_C[212][3] <=
                mat_A[208][0] * mat_B[4][3] +
                mat_A[208][1] * mat_B[12][3] +
                mat_A[208][2] * mat_B[20][3] +
                mat_A[208][3] * mat_B[28][3] +
                mat_A[209][0] * mat_B[36][3] +
                mat_A[209][1] * mat_B[44][3] +
                mat_A[209][2] * mat_B[52][3] +
                mat_A[209][3] * mat_B[60][3] +
                mat_A[210][0] * mat_B[68][3] +
                mat_A[210][1] * mat_B[76][3] +
                mat_A[210][2] * mat_B[84][3] +
                mat_A[210][3] * mat_B[92][3] +
                mat_A[211][0] * mat_B[100][3] +
                mat_A[211][1] * mat_B[108][3] +
                mat_A[211][2] * mat_B[116][3] +
                mat_A[211][3] * mat_B[124][3] +
                mat_A[212][0] * mat_B[132][3] +
                mat_A[212][1] * mat_B[140][3] +
                mat_A[212][2] * mat_B[148][3] +
                mat_A[212][3] * mat_B[156][3] +
                mat_A[213][0] * mat_B[164][3] +
                mat_A[213][1] * mat_B[172][3] +
                mat_A[213][2] * mat_B[180][3] +
                mat_A[213][3] * mat_B[188][3] +
                mat_A[214][0] * mat_B[196][3] +
                mat_A[214][1] * mat_B[204][3] +
                mat_A[214][2] * mat_B[212][3] +
                mat_A[214][3] * mat_B[220][3] +
                mat_A[215][0] * mat_B[228][3] +
                mat_A[215][1] * mat_B[236][3] +
                mat_A[215][2] * mat_B[244][3] +
                mat_A[215][3] * mat_B[252][3];
    mat_C[213][0] <=
                mat_A[208][0] * mat_B[5][0] +
                mat_A[208][1] * mat_B[13][0] +
                mat_A[208][2] * mat_B[21][0] +
                mat_A[208][3] * mat_B[29][0] +
                mat_A[209][0] * mat_B[37][0] +
                mat_A[209][1] * mat_B[45][0] +
                mat_A[209][2] * mat_B[53][0] +
                mat_A[209][3] * mat_B[61][0] +
                mat_A[210][0] * mat_B[69][0] +
                mat_A[210][1] * mat_B[77][0] +
                mat_A[210][2] * mat_B[85][0] +
                mat_A[210][3] * mat_B[93][0] +
                mat_A[211][0] * mat_B[101][0] +
                mat_A[211][1] * mat_B[109][0] +
                mat_A[211][2] * mat_B[117][0] +
                mat_A[211][3] * mat_B[125][0] +
                mat_A[212][0] * mat_B[133][0] +
                mat_A[212][1] * mat_B[141][0] +
                mat_A[212][2] * mat_B[149][0] +
                mat_A[212][3] * mat_B[157][0] +
                mat_A[213][0] * mat_B[165][0] +
                mat_A[213][1] * mat_B[173][0] +
                mat_A[213][2] * mat_B[181][0] +
                mat_A[213][3] * mat_B[189][0] +
                mat_A[214][0] * mat_B[197][0] +
                mat_A[214][1] * mat_B[205][0] +
                mat_A[214][2] * mat_B[213][0] +
                mat_A[214][3] * mat_B[221][0] +
                mat_A[215][0] * mat_B[229][0] +
                mat_A[215][1] * mat_B[237][0] +
                mat_A[215][2] * mat_B[245][0] +
                mat_A[215][3] * mat_B[253][0];
    mat_C[213][1] <=
                mat_A[208][0] * mat_B[5][1] +
                mat_A[208][1] * mat_B[13][1] +
                mat_A[208][2] * mat_B[21][1] +
                mat_A[208][3] * mat_B[29][1] +
                mat_A[209][0] * mat_B[37][1] +
                mat_A[209][1] * mat_B[45][1] +
                mat_A[209][2] * mat_B[53][1] +
                mat_A[209][3] * mat_B[61][1] +
                mat_A[210][0] * mat_B[69][1] +
                mat_A[210][1] * mat_B[77][1] +
                mat_A[210][2] * mat_B[85][1] +
                mat_A[210][3] * mat_B[93][1] +
                mat_A[211][0] * mat_B[101][1] +
                mat_A[211][1] * mat_B[109][1] +
                mat_A[211][2] * mat_B[117][1] +
                mat_A[211][3] * mat_B[125][1] +
                mat_A[212][0] * mat_B[133][1] +
                mat_A[212][1] * mat_B[141][1] +
                mat_A[212][2] * mat_B[149][1] +
                mat_A[212][3] * mat_B[157][1] +
                mat_A[213][0] * mat_B[165][1] +
                mat_A[213][1] * mat_B[173][1] +
                mat_A[213][2] * mat_B[181][1] +
                mat_A[213][3] * mat_B[189][1] +
                mat_A[214][0] * mat_B[197][1] +
                mat_A[214][1] * mat_B[205][1] +
                mat_A[214][2] * mat_B[213][1] +
                mat_A[214][3] * mat_B[221][1] +
                mat_A[215][0] * mat_B[229][1] +
                mat_A[215][1] * mat_B[237][1] +
                mat_A[215][2] * mat_B[245][1] +
                mat_A[215][3] * mat_B[253][1];
    mat_C[213][2] <=
                mat_A[208][0] * mat_B[5][2] +
                mat_A[208][1] * mat_B[13][2] +
                mat_A[208][2] * mat_B[21][2] +
                mat_A[208][3] * mat_B[29][2] +
                mat_A[209][0] * mat_B[37][2] +
                mat_A[209][1] * mat_B[45][2] +
                mat_A[209][2] * mat_B[53][2] +
                mat_A[209][3] * mat_B[61][2] +
                mat_A[210][0] * mat_B[69][2] +
                mat_A[210][1] * mat_B[77][2] +
                mat_A[210][2] * mat_B[85][2] +
                mat_A[210][3] * mat_B[93][2] +
                mat_A[211][0] * mat_B[101][2] +
                mat_A[211][1] * mat_B[109][2] +
                mat_A[211][2] * mat_B[117][2] +
                mat_A[211][3] * mat_B[125][2] +
                mat_A[212][0] * mat_B[133][2] +
                mat_A[212][1] * mat_B[141][2] +
                mat_A[212][2] * mat_B[149][2] +
                mat_A[212][3] * mat_B[157][2] +
                mat_A[213][0] * mat_B[165][2] +
                mat_A[213][1] * mat_B[173][2] +
                mat_A[213][2] * mat_B[181][2] +
                mat_A[213][3] * mat_B[189][2] +
                mat_A[214][0] * mat_B[197][2] +
                mat_A[214][1] * mat_B[205][2] +
                mat_A[214][2] * mat_B[213][2] +
                mat_A[214][3] * mat_B[221][2] +
                mat_A[215][0] * mat_B[229][2] +
                mat_A[215][1] * mat_B[237][2] +
                mat_A[215][2] * mat_B[245][2] +
                mat_A[215][3] * mat_B[253][2];
    mat_C[213][3] <=
                mat_A[208][0] * mat_B[5][3] +
                mat_A[208][1] * mat_B[13][3] +
                mat_A[208][2] * mat_B[21][3] +
                mat_A[208][3] * mat_B[29][3] +
                mat_A[209][0] * mat_B[37][3] +
                mat_A[209][1] * mat_B[45][3] +
                mat_A[209][2] * mat_B[53][3] +
                mat_A[209][3] * mat_B[61][3] +
                mat_A[210][0] * mat_B[69][3] +
                mat_A[210][1] * mat_B[77][3] +
                mat_A[210][2] * mat_B[85][3] +
                mat_A[210][3] * mat_B[93][3] +
                mat_A[211][0] * mat_B[101][3] +
                mat_A[211][1] * mat_B[109][3] +
                mat_A[211][2] * mat_B[117][3] +
                mat_A[211][3] * mat_B[125][3] +
                mat_A[212][0] * mat_B[133][3] +
                mat_A[212][1] * mat_B[141][3] +
                mat_A[212][2] * mat_B[149][3] +
                mat_A[212][3] * mat_B[157][3] +
                mat_A[213][0] * mat_B[165][3] +
                mat_A[213][1] * mat_B[173][3] +
                mat_A[213][2] * mat_B[181][3] +
                mat_A[213][3] * mat_B[189][3] +
                mat_A[214][0] * mat_B[197][3] +
                mat_A[214][1] * mat_B[205][3] +
                mat_A[214][2] * mat_B[213][3] +
                mat_A[214][3] * mat_B[221][3] +
                mat_A[215][0] * mat_B[229][3] +
                mat_A[215][1] * mat_B[237][3] +
                mat_A[215][2] * mat_B[245][3] +
                mat_A[215][3] * mat_B[253][3];
    mat_C[214][0] <=
                mat_A[208][0] * mat_B[6][0] +
                mat_A[208][1] * mat_B[14][0] +
                mat_A[208][2] * mat_B[22][0] +
                mat_A[208][3] * mat_B[30][0] +
                mat_A[209][0] * mat_B[38][0] +
                mat_A[209][1] * mat_B[46][0] +
                mat_A[209][2] * mat_B[54][0] +
                mat_A[209][3] * mat_B[62][0] +
                mat_A[210][0] * mat_B[70][0] +
                mat_A[210][1] * mat_B[78][0] +
                mat_A[210][2] * mat_B[86][0] +
                mat_A[210][3] * mat_B[94][0] +
                mat_A[211][0] * mat_B[102][0] +
                mat_A[211][1] * mat_B[110][0] +
                mat_A[211][2] * mat_B[118][0] +
                mat_A[211][3] * mat_B[126][0] +
                mat_A[212][0] * mat_B[134][0] +
                mat_A[212][1] * mat_B[142][0] +
                mat_A[212][2] * mat_B[150][0] +
                mat_A[212][3] * mat_B[158][0] +
                mat_A[213][0] * mat_B[166][0] +
                mat_A[213][1] * mat_B[174][0] +
                mat_A[213][2] * mat_B[182][0] +
                mat_A[213][3] * mat_B[190][0] +
                mat_A[214][0] * mat_B[198][0] +
                mat_A[214][1] * mat_B[206][0] +
                mat_A[214][2] * mat_B[214][0] +
                mat_A[214][3] * mat_B[222][0] +
                mat_A[215][0] * mat_B[230][0] +
                mat_A[215][1] * mat_B[238][0] +
                mat_A[215][2] * mat_B[246][0] +
                mat_A[215][3] * mat_B[254][0];
    mat_C[214][1] <=
                mat_A[208][0] * mat_B[6][1] +
                mat_A[208][1] * mat_B[14][1] +
                mat_A[208][2] * mat_B[22][1] +
                mat_A[208][3] * mat_B[30][1] +
                mat_A[209][0] * mat_B[38][1] +
                mat_A[209][1] * mat_B[46][1] +
                mat_A[209][2] * mat_B[54][1] +
                mat_A[209][3] * mat_B[62][1] +
                mat_A[210][0] * mat_B[70][1] +
                mat_A[210][1] * mat_B[78][1] +
                mat_A[210][2] * mat_B[86][1] +
                mat_A[210][3] * mat_B[94][1] +
                mat_A[211][0] * mat_B[102][1] +
                mat_A[211][1] * mat_B[110][1] +
                mat_A[211][2] * mat_B[118][1] +
                mat_A[211][3] * mat_B[126][1] +
                mat_A[212][0] * mat_B[134][1] +
                mat_A[212][1] * mat_B[142][1] +
                mat_A[212][2] * mat_B[150][1] +
                mat_A[212][3] * mat_B[158][1] +
                mat_A[213][0] * mat_B[166][1] +
                mat_A[213][1] * mat_B[174][1] +
                mat_A[213][2] * mat_B[182][1] +
                mat_A[213][3] * mat_B[190][1] +
                mat_A[214][0] * mat_B[198][1] +
                mat_A[214][1] * mat_B[206][1] +
                mat_A[214][2] * mat_B[214][1] +
                mat_A[214][3] * mat_B[222][1] +
                mat_A[215][0] * mat_B[230][1] +
                mat_A[215][1] * mat_B[238][1] +
                mat_A[215][2] * mat_B[246][1] +
                mat_A[215][3] * mat_B[254][1];
    mat_C[214][2] <=
                mat_A[208][0] * mat_B[6][2] +
                mat_A[208][1] * mat_B[14][2] +
                mat_A[208][2] * mat_B[22][2] +
                mat_A[208][3] * mat_B[30][2] +
                mat_A[209][0] * mat_B[38][2] +
                mat_A[209][1] * mat_B[46][2] +
                mat_A[209][2] * mat_B[54][2] +
                mat_A[209][3] * mat_B[62][2] +
                mat_A[210][0] * mat_B[70][2] +
                mat_A[210][1] * mat_B[78][2] +
                mat_A[210][2] * mat_B[86][2] +
                mat_A[210][3] * mat_B[94][2] +
                mat_A[211][0] * mat_B[102][2] +
                mat_A[211][1] * mat_B[110][2] +
                mat_A[211][2] * mat_B[118][2] +
                mat_A[211][3] * mat_B[126][2] +
                mat_A[212][0] * mat_B[134][2] +
                mat_A[212][1] * mat_B[142][2] +
                mat_A[212][2] * mat_B[150][2] +
                mat_A[212][3] * mat_B[158][2] +
                mat_A[213][0] * mat_B[166][2] +
                mat_A[213][1] * mat_B[174][2] +
                mat_A[213][2] * mat_B[182][2] +
                mat_A[213][3] * mat_B[190][2] +
                mat_A[214][0] * mat_B[198][2] +
                mat_A[214][1] * mat_B[206][2] +
                mat_A[214][2] * mat_B[214][2] +
                mat_A[214][3] * mat_B[222][2] +
                mat_A[215][0] * mat_B[230][2] +
                mat_A[215][1] * mat_B[238][2] +
                mat_A[215][2] * mat_B[246][2] +
                mat_A[215][3] * mat_B[254][2];
    mat_C[214][3] <=
                mat_A[208][0] * mat_B[6][3] +
                mat_A[208][1] * mat_B[14][3] +
                mat_A[208][2] * mat_B[22][3] +
                mat_A[208][3] * mat_B[30][3] +
                mat_A[209][0] * mat_B[38][3] +
                mat_A[209][1] * mat_B[46][3] +
                mat_A[209][2] * mat_B[54][3] +
                mat_A[209][3] * mat_B[62][3] +
                mat_A[210][0] * mat_B[70][3] +
                mat_A[210][1] * mat_B[78][3] +
                mat_A[210][2] * mat_B[86][3] +
                mat_A[210][3] * mat_B[94][3] +
                mat_A[211][0] * mat_B[102][3] +
                mat_A[211][1] * mat_B[110][3] +
                mat_A[211][2] * mat_B[118][3] +
                mat_A[211][3] * mat_B[126][3] +
                mat_A[212][0] * mat_B[134][3] +
                mat_A[212][1] * mat_B[142][3] +
                mat_A[212][2] * mat_B[150][3] +
                mat_A[212][3] * mat_B[158][3] +
                mat_A[213][0] * mat_B[166][3] +
                mat_A[213][1] * mat_B[174][3] +
                mat_A[213][2] * mat_B[182][3] +
                mat_A[213][3] * mat_B[190][3] +
                mat_A[214][0] * mat_B[198][3] +
                mat_A[214][1] * mat_B[206][3] +
                mat_A[214][2] * mat_B[214][3] +
                mat_A[214][3] * mat_B[222][3] +
                mat_A[215][0] * mat_B[230][3] +
                mat_A[215][1] * mat_B[238][3] +
                mat_A[215][2] * mat_B[246][3] +
                mat_A[215][3] * mat_B[254][3];
    mat_C[215][0] <=
                mat_A[208][0] * mat_B[7][0] +
                mat_A[208][1] * mat_B[15][0] +
                mat_A[208][2] * mat_B[23][0] +
                mat_A[208][3] * mat_B[31][0] +
                mat_A[209][0] * mat_B[39][0] +
                mat_A[209][1] * mat_B[47][0] +
                mat_A[209][2] * mat_B[55][0] +
                mat_A[209][3] * mat_B[63][0] +
                mat_A[210][0] * mat_B[71][0] +
                mat_A[210][1] * mat_B[79][0] +
                mat_A[210][2] * mat_B[87][0] +
                mat_A[210][3] * mat_B[95][0] +
                mat_A[211][0] * mat_B[103][0] +
                mat_A[211][1] * mat_B[111][0] +
                mat_A[211][2] * mat_B[119][0] +
                mat_A[211][3] * mat_B[127][0] +
                mat_A[212][0] * mat_B[135][0] +
                mat_A[212][1] * mat_B[143][0] +
                mat_A[212][2] * mat_B[151][0] +
                mat_A[212][3] * mat_B[159][0] +
                mat_A[213][0] * mat_B[167][0] +
                mat_A[213][1] * mat_B[175][0] +
                mat_A[213][2] * mat_B[183][0] +
                mat_A[213][3] * mat_B[191][0] +
                mat_A[214][0] * mat_B[199][0] +
                mat_A[214][1] * mat_B[207][0] +
                mat_A[214][2] * mat_B[215][0] +
                mat_A[214][3] * mat_B[223][0] +
                mat_A[215][0] * mat_B[231][0] +
                mat_A[215][1] * mat_B[239][0] +
                mat_A[215][2] * mat_B[247][0] +
                mat_A[215][3] * mat_B[255][0];
    mat_C[215][1] <=
                mat_A[208][0] * mat_B[7][1] +
                mat_A[208][1] * mat_B[15][1] +
                mat_A[208][2] * mat_B[23][1] +
                mat_A[208][3] * mat_B[31][1] +
                mat_A[209][0] * mat_B[39][1] +
                mat_A[209][1] * mat_B[47][1] +
                mat_A[209][2] * mat_B[55][1] +
                mat_A[209][3] * mat_B[63][1] +
                mat_A[210][0] * mat_B[71][1] +
                mat_A[210][1] * mat_B[79][1] +
                mat_A[210][2] * mat_B[87][1] +
                mat_A[210][3] * mat_B[95][1] +
                mat_A[211][0] * mat_B[103][1] +
                mat_A[211][1] * mat_B[111][1] +
                mat_A[211][2] * mat_B[119][1] +
                mat_A[211][3] * mat_B[127][1] +
                mat_A[212][0] * mat_B[135][1] +
                mat_A[212][1] * mat_B[143][1] +
                mat_A[212][2] * mat_B[151][1] +
                mat_A[212][3] * mat_B[159][1] +
                mat_A[213][0] * mat_B[167][1] +
                mat_A[213][1] * mat_B[175][1] +
                mat_A[213][2] * mat_B[183][1] +
                mat_A[213][3] * mat_B[191][1] +
                mat_A[214][0] * mat_B[199][1] +
                mat_A[214][1] * mat_B[207][1] +
                mat_A[214][2] * mat_B[215][1] +
                mat_A[214][3] * mat_B[223][1] +
                mat_A[215][0] * mat_B[231][1] +
                mat_A[215][1] * mat_B[239][1] +
                mat_A[215][2] * mat_B[247][1] +
                mat_A[215][3] * mat_B[255][1];
    mat_C[215][2] <=
                mat_A[208][0] * mat_B[7][2] +
                mat_A[208][1] * mat_B[15][2] +
                mat_A[208][2] * mat_B[23][2] +
                mat_A[208][3] * mat_B[31][2] +
                mat_A[209][0] * mat_B[39][2] +
                mat_A[209][1] * mat_B[47][2] +
                mat_A[209][2] * mat_B[55][2] +
                mat_A[209][3] * mat_B[63][2] +
                mat_A[210][0] * mat_B[71][2] +
                mat_A[210][1] * mat_B[79][2] +
                mat_A[210][2] * mat_B[87][2] +
                mat_A[210][3] * mat_B[95][2] +
                mat_A[211][0] * mat_B[103][2] +
                mat_A[211][1] * mat_B[111][2] +
                mat_A[211][2] * mat_B[119][2] +
                mat_A[211][3] * mat_B[127][2] +
                mat_A[212][0] * mat_B[135][2] +
                mat_A[212][1] * mat_B[143][2] +
                mat_A[212][2] * mat_B[151][2] +
                mat_A[212][3] * mat_B[159][2] +
                mat_A[213][0] * mat_B[167][2] +
                mat_A[213][1] * mat_B[175][2] +
                mat_A[213][2] * mat_B[183][2] +
                mat_A[213][3] * mat_B[191][2] +
                mat_A[214][0] * mat_B[199][2] +
                mat_A[214][1] * mat_B[207][2] +
                mat_A[214][2] * mat_B[215][2] +
                mat_A[214][3] * mat_B[223][2] +
                mat_A[215][0] * mat_B[231][2] +
                mat_A[215][1] * mat_B[239][2] +
                mat_A[215][2] * mat_B[247][2] +
                mat_A[215][3] * mat_B[255][2];
    mat_C[215][3] <=
                mat_A[208][0] * mat_B[7][3] +
                mat_A[208][1] * mat_B[15][3] +
                mat_A[208][2] * mat_B[23][3] +
                mat_A[208][3] * mat_B[31][3] +
                mat_A[209][0] * mat_B[39][3] +
                mat_A[209][1] * mat_B[47][3] +
                mat_A[209][2] * mat_B[55][3] +
                mat_A[209][3] * mat_B[63][3] +
                mat_A[210][0] * mat_B[71][3] +
                mat_A[210][1] * mat_B[79][3] +
                mat_A[210][2] * mat_B[87][3] +
                mat_A[210][3] * mat_B[95][3] +
                mat_A[211][0] * mat_B[103][3] +
                mat_A[211][1] * mat_B[111][3] +
                mat_A[211][2] * mat_B[119][3] +
                mat_A[211][3] * mat_B[127][3] +
                mat_A[212][0] * mat_B[135][3] +
                mat_A[212][1] * mat_B[143][3] +
                mat_A[212][2] * mat_B[151][3] +
                mat_A[212][3] * mat_B[159][3] +
                mat_A[213][0] * mat_B[167][3] +
                mat_A[213][1] * mat_B[175][3] +
                mat_A[213][2] * mat_B[183][3] +
                mat_A[213][3] * mat_B[191][3] +
                mat_A[214][0] * mat_B[199][3] +
                mat_A[214][1] * mat_B[207][3] +
                mat_A[214][2] * mat_B[215][3] +
                mat_A[214][3] * mat_B[223][3] +
                mat_A[215][0] * mat_B[231][3] +
                mat_A[215][1] * mat_B[239][3] +
                mat_A[215][2] * mat_B[247][3] +
                mat_A[215][3] * mat_B[255][3];
    mat_C[216][0] <=
                mat_A[216][0] * mat_B[0][0] +
                mat_A[216][1] * mat_B[8][0] +
                mat_A[216][2] * mat_B[16][0] +
                mat_A[216][3] * mat_B[24][0] +
                mat_A[217][0] * mat_B[32][0] +
                mat_A[217][1] * mat_B[40][0] +
                mat_A[217][2] * mat_B[48][0] +
                mat_A[217][3] * mat_B[56][0] +
                mat_A[218][0] * mat_B[64][0] +
                mat_A[218][1] * mat_B[72][0] +
                mat_A[218][2] * mat_B[80][0] +
                mat_A[218][3] * mat_B[88][0] +
                mat_A[219][0] * mat_B[96][0] +
                mat_A[219][1] * mat_B[104][0] +
                mat_A[219][2] * mat_B[112][0] +
                mat_A[219][3] * mat_B[120][0] +
                mat_A[220][0] * mat_B[128][0] +
                mat_A[220][1] * mat_B[136][0] +
                mat_A[220][2] * mat_B[144][0] +
                mat_A[220][3] * mat_B[152][0] +
                mat_A[221][0] * mat_B[160][0] +
                mat_A[221][1] * mat_B[168][0] +
                mat_A[221][2] * mat_B[176][0] +
                mat_A[221][3] * mat_B[184][0] +
                mat_A[222][0] * mat_B[192][0] +
                mat_A[222][1] * mat_B[200][0] +
                mat_A[222][2] * mat_B[208][0] +
                mat_A[222][3] * mat_B[216][0] +
                mat_A[223][0] * mat_B[224][0] +
                mat_A[223][1] * mat_B[232][0] +
                mat_A[223][2] * mat_B[240][0] +
                mat_A[223][3] * mat_B[248][0];
    mat_C[216][1] <=
                mat_A[216][0] * mat_B[0][1] +
                mat_A[216][1] * mat_B[8][1] +
                mat_A[216][2] * mat_B[16][1] +
                mat_A[216][3] * mat_B[24][1] +
                mat_A[217][0] * mat_B[32][1] +
                mat_A[217][1] * mat_B[40][1] +
                mat_A[217][2] * mat_B[48][1] +
                mat_A[217][3] * mat_B[56][1] +
                mat_A[218][0] * mat_B[64][1] +
                mat_A[218][1] * mat_B[72][1] +
                mat_A[218][2] * mat_B[80][1] +
                mat_A[218][3] * mat_B[88][1] +
                mat_A[219][0] * mat_B[96][1] +
                mat_A[219][1] * mat_B[104][1] +
                mat_A[219][2] * mat_B[112][1] +
                mat_A[219][3] * mat_B[120][1] +
                mat_A[220][0] * mat_B[128][1] +
                mat_A[220][1] * mat_B[136][1] +
                mat_A[220][2] * mat_B[144][1] +
                mat_A[220][3] * mat_B[152][1] +
                mat_A[221][0] * mat_B[160][1] +
                mat_A[221][1] * mat_B[168][1] +
                mat_A[221][2] * mat_B[176][1] +
                mat_A[221][3] * mat_B[184][1] +
                mat_A[222][0] * mat_B[192][1] +
                mat_A[222][1] * mat_B[200][1] +
                mat_A[222][2] * mat_B[208][1] +
                mat_A[222][3] * mat_B[216][1] +
                mat_A[223][0] * mat_B[224][1] +
                mat_A[223][1] * mat_B[232][1] +
                mat_A[223][2] * mat_B[240][1] +
                mat_A[223][3] * mat_B[248][1];
    mat_C[216][2] <=
                mat_A[216][0] * mat_B[0][2] +
                mat_A[216][1] * mat_B[8][2] +
                mat_A[216][2] * mat_B[16][2] +
                mat_A[216][3] * mat_B[24][2] +
                mat_A[217][0] * mat_B[32][2] +
                mat_A[217][1] * mat_B[40][2] +
                mat_A[217][2] * mat_B[48][2] +
                mat_A[217][3] * mat_B[56][2] +
                mat_A[218][0] * mat_B[64][2] +
                mat_A[218][1] * mat_B[72][2] +
                mat_A[218][2] * mat_B[80][2] +
                mat_A[218][3] * mat_B[88][2] +
                mat_A[219][0] * mat_B[96][2] +
                mat_A[219][1] * mat_B[104][2] +
                mat_A[219][2] * mat_B[112][2] +
                mat_A[219][3] * mat_B[120][2] +
                mat_A[220][0] * mat_B[128][2] +
                mat_A[220][1] * mat_B[136][2] +
                mat_A[220][2] * mat_B[144][2] +
                mat_A[220][3] * mat_B[152][2] +
                mat_A[221][0] * mat_B[160][2] +
                mat_A[221][1] * mat_B[168][2] +
                mat_A[221][2] * mat_B[176][2] +
                mat_A[221][3] * mat_B[184][2] +
                mat_A[222][0] * mat_B[192][2] +
                mat_A[222][1] * mat_B[200][2] +
                mat_A[222][2] * mat_B[208][2] +
                mat_A[222][3] * mat_B[216][2] +
                mat_A[223][0] * mat_B[224][2] +
                mat_A[223][1] * mat_B[232][2] +
                mat_A[223][2] * mat_B[240][2] +
                mat_A[223][3] * mat_B[248][2];
    mat_C[216][3] <=
                mat_A[216][0] * mat_B[0][3] +
                mat_A[216][1] * mat_B[8][3] +
                mat_A[216][2] * mat_B[16][3] +
                mat_A[216][3] * mat_B[24][3] +
                mat_A[217][0] * mat_B[32][3] +
                mat_A[217][1] * mat_B[40][3] +
                mat_A[217][2] * mat_B[48][3] +
                mat_A[217][3] * mat_B[56][3] +
                mat_A[218][0] * mat_B[64][3] +
                mat_A[218][1] * mat_B[72][3] +
                mat_A[218][2] * mat_B[80][3] +
                mat_A[218][3] * mat_B[88][3] +
                mat_A[219][0] * mat_B[96][3] +
                mat_A[219][1] * mat_B[104][3] +
                mat_A[219][2] * mat_B[112][3] +
                mat_A[219][3] * mat_B[120][3] +
                mat_A[220][0] * mat_B[128][3] +
                mat_A[220][1] * mat_B[136][3] +
                mat_A[220][2] * mat_B[144][3] +
                mat_A[220][3] * mat_B[152][3] +
                mat_A[221][0] * mat_B[160][3] +
                mat_A[221][1] * mat_B[168][3] +
                mat_A[221][2] * mat_B[176][3] +
                mat_A[221][3] * mat_B[184][3] +
                mat_A[222][0] * mat_B[192][3] +
                mat_A[222][1] * mat_B[200][3] +
                mat_A[222][2] * mat_B[208][3] +
                mat_A[222][3] * mat_B[216][3] +
                mat_A[223][0] * mat_B[224][3] +
                mat_A[223][1] * mat_B[232][3] +
                mat_A[223][2] * mat_B[240][3] +
                mat_A[223][3] * mat_B[248][3];
    mat_C[217][0] <=
                mat_A[216][0] * mat_B[1][0] +
                mat_A[216][1] * mat_B[9][0] +
                mat_A[216][2] * mat_B[17][0] +
                mat_A[216][3] * mat_B[25][0] +
                mat_A[217][0] * mat_B[33][0] +
                mat_A[217][1] * mat_B[41][0] +
                mat_A[217][2] * mat_B[49][0] +
                mat_A[217][3] * mat_B[57][0] +
                mat_A[218][0] * mat_B[65][0] +
                mat_A[218][1] * mat_B[73][0] +
                mat_A[218][2] * mat_B[81][0] +
                mat_A[218][3] * mat_B[89][0] +
                mat_A[219][0] * mat_B[97][0] +
                mat_A[219][1] * mat_B[105][0] +
                mat_A[219][2] * mat_B[113][0] +
                mat_A[219][3] * mat_B[121][0] +
                mat_A[220][0] * mat_B[129][0] +
                mat_A[220][1] * mat_B[137][0] +
                mat_A[220][2] * mat_B[145][0] +
                mat_A[220][3] * mat_B[153][0] +
                mat_A[221][0] * mat_B[161][0] +
                mat_A[221][1] * mat_B[169][0] +
                mat_A[221][2] * mat_B[177][0] +
                mat_A[221][3] * mat_B[185][0] +
                mat_A[222][0] * mat_B[193][0] +
                mat_A[222][1] * mat_B[201][0] +
                mat_A[222][2] * mat_B[209][0] +
                mat_A[222][3] * mat_B[217][0] +
                mat_A[223][0] * mat_B[225][0] +
                mat_A[223][1] * mat_B[233][0] +
                mat_A[223][2] * mat_B[241][0] +
                mat_A[223][3] * mat_B[249][0];
    mat_C[217][1] <=
                mat_A[216][0] * mat_B[1][1] +
                mat_A[216][1] * mat_B[9][1] +
                mat_A[216][2] * mat_B[17][1] +
                mat_A[216][3] * mat_B[25][1] +
                mat_A[217][0] * mat_B[33][1] +
                mat_A[217][1] * mat_B[41][1] +
                mat_A[217][2] * mat_B[49][1] +
                mat_A[217][3] * mat_B[57][1] +
                mat_A[218][0] * mat_B[65][1] +
                mat_A[218][1] * mat_B[73][1] +
                mat_A[218][2] * mat_B[81][1] +
                mat_A[218][3] * mat_B[89][1] +
                mat_A[219][0] * mat_B[97][1] +
                mat_A[219][1] * mat_B[105][1] +
                mat_A[219][2] * mat_B[113][1] +
                mat_A[219][3] * mat_B[121][1] +
                mat_A[220][0] * mat_B[129][1] +
                mat_A[220][1] * mat_B[137][1] +
                mat_A[220][2] * mat_B[145][1] +
                mat_A[220][3] * mat_B[153][1] +
                mat_A[221][0] * mat_B[161][1] +
                mat_A[221][1] * mat_B[169][1] +
                mat_A[221][2] * mat_B[177][1] +
                mat_A[221][3] * mat_B[185][1] +
                mat_A[222][0] * mat_B[193][1] +
                mat_A[222][1] * mat_B[201][1] +
                mat_A[222][2] * mat_B[209][1] +
                mat_A[222][3] * mat_B[217][1] +
                mat_A[223][0] * mat_B[225][1] +
                mat_A[223][1] * mat_B[233][1] +
                mat_A[223][2] * mat_B[241][1] +
                mat_A[223][3] * mat_B[249][1];
    mat_C[217][2] <=
                mat_A[216][0] * mat_B[1][2] +
                mat_A[216][1] * mat_B[9][2] +
                mat_A[216][2] * mat_B[17][2] +
                mat_A[216][3] * mat_B[25][2] +
                mat_A[217][0] * mat_B[33][2] +
                mat_A[217][1] * mat_B[41][2] +
                mat_A[217][2] * mat_B[49][2] +
                mat_A[217][3] * mat_B[57][2] +
                mat_A[218][0] * mat_B[65][2] +
                mat_A[218][1] * mat_B[73][2] +
                mat_A[218][2] * mat_B[81][2] +
                mat_A[218][3] * mat_B[89][2] +
                mat_A[219][0] * mat_B[97][2] +
                mat_A[219][1] * mat_B[105][2] +
                mat_A[219][2] * mat_B[113][2] +
                mat_A[219][3] * mat_B[121][2] +
                mat_A[220][0] * mat_B[129][2] +
                mat_A[220][1] * mat_B[137][2] +
                mat_A[220][2] * mat_B[145][2] +
                mat_A[220][3] * mat_B[153][2] +
                mat_A[221][0] * mat_B[161][2] +
                mat_A[221][1] * mat_B[169][2] +
                mat_A[221][2] * mat_B[177][2] +
                mat_A[221][3] * mat_B[185][2] +
                mat_A[222][0] * mat_B[193][2] +
                mat_A[222][1] * mat_B[201][2] +
                mat_A[222][2] * mat_B[209][2] +
                mat_A[222][3] * mat_B[217][2] +
                mat_A[223][0] * mat_B[225][2] +
                mat_A[223][1] * mat_B[233][2] +
                mat_A[223][2] * mat_B[241][2] +
                mat_A[223][3] * mat_B[249][2];
    mat_C[217][3] <=
                mat_A[216][0] * mat_B[1][3] +
                mat_A[216][1] * mat_B[9][3] +
                mat_A[216][2] * mat_B[17][3] +
                mat_A[216][3] * mat_B[25][3] +
                mat_A[217][0] * mat_B[33][3] +
                mat_A[217][1] * mat_B[41][3] +
                mat_A[217][2] * mat_B[49][3] +
                mat_A[217][3] * mat_B[57][3] +
                mat_A[218][0] * mat_B[65][3] +
                mat_A[218][1] * mat_B[73][3] +
                mat_A[218][2] * mat_B[81][3] +
                mat_A[218][3] * mat_B[89][3] +
                mat_A[219][0] * mat_B[97][3] +
                mat_A[219][1] * mat_B[105][3] +
                mat_A[219][2] * mat_B[113][3] +
                mat_A[219][3] * mat_B[121][3] +
                mat_A[220][0] * mat_B[129][3] +
                mat_A[220][1] * mat_B[137][3] +
                mat_A[220][2] * mat_B[145][3] +
                mat_A[220][3] * mat_B[153][3] +
                mat_A[221][0] * mat_B[161][3] +
                mat_A[221][1] * mat_B[169][3] +
                mat_A[221][2] * mat_B[177][3] +
                mat_A[221][3] * mat_B[185][3] +
                mat_A[222][0] * mat_B[193][3] +
                mat_A[222][1] * mat_B[201][3] +
                mat_A[222][2] * mat_B[209][3] +
                mat_A[222][3] * mat_B[217][3] +
                mat_A[223][0] * mat_B[225][3] +
                mat_A[223][1] * mat_B[233][3] +
                mat_A[223][2] * mat_B[241][3] +
                mat_A[223][3] * mat_B[249][3];
    mat_C[218][0] <=
                mat_A[216][0] * mat_B[2][0] +
                mat_A[216][1] * mat_B[10][0] +
                mat_A[216][2] * mat_B[18][0] +
                mat_A[216][3] * mat_B[26][0] +
                mat_A[217][0] * mat_B[34][0] +
                mat_A[217][1] * mat_B[42][0] +
                mat_A[217][2] * mat_B[50][0] +
                mat_A[217][3] * mat_B[58][0] +
                mat_A[218][0] * mat_B[66][0] +
                mat_A[218][1] * mat_B[74][0] +
                mat_A[218][2] * mat_B[82][0] +
                mat_A[218][3] * mat_B[90][0] +
                mat_A[219][0] * mat_B[98][0] +
                mat_A[219][1] * mat_B[106][0] +
                mat_A[219][2] * mat_B[114][0] +
                mat_A[219][3] * mat_B[122][0] +
                mat_A[220][0] * mat_B[130][0] +
                mat_A[220][1] * mat_B[138][0] +
                mat_A[220][2] * mat_B[146][0] +
                mat_A[220][3] * mat_B[154][0] +
                mat_A[221][0] * mat_B[162][0] +
                mat_A[221][1] * mat_B[170][0] +
                mat_A[221][2] * mat_B[178][0] +
                mat_A[221][3] * mat_B[186][0] +
                mat_A[222][0] * mat_B[194][0] +
                mat_A[222][1] * mat_B[202][0] +
                mat_A[222][2] * mat_B[210][0] +
                mat_A[222][3] * mat_B[218][0] +
                mat_A[223][0] * mat_B[226][0] +
                mat_A[223][1] * mat_B[234][0] +
                mat_A[223][2] * mat_B[242][0] +
                mat_A[223][3] * mat_B[250][0];
    mat_C[218][1] <=
                mat_A[216][0] * mat_B[2][1] +
                mat_A[216][1] * mat_B[10][1] +
                mat_A[216][2] * mat_B[18][1] +
                mat_A[216][3] * mat_B[26][1] +
                mat_A[217][0] * mat_B[34][1] +
                mat_A[217][1] * mat_B[42][1] +
                mat_A[217][2] * mat_B[50][1] +
                mat_A[217][3] * mat_B[58][1] +
                mat_A[218][0] * mat_B[66][1] +
                mat_A[218][1] * mat_B[74][1] +
                mat_A[218][2] * mat_B[82][1] +
                mat_A[218][3] * mat_B[90][1] +
                mat_A[219][0] * mat_B[98][1] +
                mat_A[219][1] * mat_B[106][1] +
                mat_A[219][2] * mat_B[114][1] +
                mat_A[219][3] * mat_B[122][1] +
                mat_A[220][0] * mat_B[130][1] +
                mat_A[220][1] * mat_B[138][1] +
                mat_A[220][2] * mat_B[146][1] +
                mat_A[220][3] * mat_B[154][1] +
                mat_A[221][0] * mat_B[162][1] +
                mat_A[221][1] * mat_B[170][1] +
                mat_A[221][2] * mat_B[178][1] +
                mat_A[221][3] * mat_B[186][1] +
                mat_A[222][0] * mat_B[194][1] +
                mat_A[222][1] * mat_B[202][1] +
                mat_A[222][2] * mat_B[210][1] +
                mat_A[222][3] * mat_B[218][1] +
                mat_A[223][0] * mat_B[226][1] +
                mat_A[223][1] * mat_B[234][1] +
                mat_A[223][2] * mat_B[242][1] +
                mat_A[223][3] * mat_B[250][1];
    mat_C[218][2] <=
                mat_A[216][0] * mat_B[2][2] +
                mat_A[216][1] * mat_B[10][2] +
                mat_A[216][2] * mat_B[18][2] +
                mat_A[216][3] * mat_B[26][2] +
                mat_A[217][0] * mat_B[34][2] +
                mat_A[217][1] * mat_B[42][2] +
                mat_A[217][2] * mat_B[50][2] +
                mat_A[217][3] * mat_B[58][2] +
                mat_A[218][0] * mat_B[66][2] +
                mat_A[218][1] * mat_B[74][2] +
                mat_A[218][2] * mat_B[82][2] +
                mat_A[218][3] * mat_B[90][2] +
                mat_A[219][0] * mat_B[98][2] +
                mat_A[219][1] * mat_B[106][2] +
                mat_A[219][2] * mat_B[114][2] +
                mat_A[219][3] * mat_B[122][2] +
                mat_A[220][0] * mat_B[130][2] +
                mat_A[220][1] * mat_B[138][2] +
                mat_A[220][2] * mat_B[146][2] +
                mat_A[220][3] * mat_B[154][2] +
                mat_A[221][0] * mat_B[162][2] +
                mat_A[221][1] * mat_B[170][2] +
                mat_A[221][2] * mat_B[178][2] +
                mat_A[221][3] * mat_B[186][2] +
                mat_A[222][0] * mat_B[194][2] +
                mat_A[222][1] * mat_B[202][2] +
                mat_A[222][2] * mat_B[210][2] +
                mat_A[222][3] * mat_B[218][2] +
                mat_A[223][0] * mat_B[226][2] +
                mat_A[223][1] * mat_B[234][2] +
                mat_A[223][2] * mat_B[242][2] +
                mat_A[223][3] * mat_B[250][2];
    mat_C[218][3] <=
                mat_A[216][0] * mat_B[2][3] +
                mat_A[216][1] * mat_B[10][3] +
                mat_A[216][2] * mat_B[18][3] +
                mat_A[216][3] * mat_B[26][3] +
                mat_A[217][0] * mat_B[34][3] +
                mat_A[217][1] * mat_B[42][3] +
                mat_A[217][2] * mat_B[50][3] +
                mat_A[217][3] * mat_B[58][3] +
                mat_A[218][0] * mat_B[66][3] +
                mat_A[218][1] * mat_B[74][3] +
                mat_A[218][2] * mat_B[82][3] +
                mat_A[218][3] * mat_B[90][3] +
                mat_A[219][0] * mat_B[98][3] +
                mat_A[219][1] * mat_B[106][3] +
                mat_A[219][2] * mat_B[114][3] +
                mat_A[219][3] * mat_B[122][3] +
                mat_A[220][0] * mat_B[130][3] +
                mat_A[220][1] * mat_B[138][3] +
                mat_A[220][2] * mat_B[146][3] +
                mat_A[220][3] * mat_B[154][3] +
                mat_A[221][0] * mat_B[162][3] +
                mat_A[221][1] * mat_B[170][3] +
                mat_A[221][2] * mat_B[178][3] +
                mat_A[221][3] * mat_B[186][3] +
                mat_A[222][0] * mat_B[194][3] +
                mat_A[222][1] * mat_B[202][3] +
                mat_A[222][2] * mat_B[210][3] +
                mat_A[222][3] * mat_B[218][3] +
                mat_A[223][0] * mat_B[226][3] +
                mat_A[223][1] * mat_B[234][3] +
                mat_A[223][2] * mat_B[242][3] +
                mat_A[223][3] * mat_B[250][3];
    mat_C[219][0] <=
                mat_A[216][0] * mat_B[3][0] +
                mat_A[216][1] * mat_B[11][0] +
                mat_A[216][2] * mat_B[19][0] +
                mat_A[216][3] * mat_B[27][0] +
                mat_A[217][0] * mat_B[35][0] +
                mat_A[217][1] * mat_B[43][0] +
                mat_A[217][2] * mat_B[51][0] +
                mat_A[217][3] * mat_B[59][0] +
                mat_A[218][0] * mat_B[67][0] +
                mat_A[218][1] * mat_B[75][0] +
                mat_A[218][2] * mat_B[83][0] +
                mat_A[218][3] * mat_B[91][0] +
                mat_A[219][0] * mat_B[99][0] +
                mat_A[219][1] * mat_B[107][0] +
                mat_A[219][2] * mat_B[115][0] +
                mat_A[219][3] * mat_B[123][0] +
                mat_A[220][0] * mat_B[131][0] +
                mat_A[220][1] * mat_B[139][0] +
                mat_A[220][2] * mat_B[147][0] +
                mat_A[220][3] * mat_B[155][0] +
                mat_A[221][0] * mat_B[163][0] +
                mat_A[221][1] * mat_B[171][0] +
                mat_A[221][2] * mat_B[179][0] +
                mat_A[221][3] * mat_B[187][0] +
                mat_A[222][0] * mat_B[195][0] +
                mat_A[222][1] * mat_B[203][0] +
                mat_A[222][2] * mat_B[211][0] +
                mat_A[222][3] * mat_B[219][0] +
                mat_A[223][0] * mat_B[227][0] +
                mat_A[223][1] * mat_B[235][0] +
                mat_A[223][2] * mat_B[243][0] +
                mat_A[223][3] * mat_B[251][0];
    mat_C[219][1] <=
                mat_A[216][0] * mat_B[3][1] +
                mat_A[216][1] * mat_B[11][1] +
                mat_A[216][2] * mat_B[19][1] +
                mat_A[216][3] * mat_B[27][1] +
                mat_A[217][0] * mat_B[35][1] +
                mat_A[217][1] * mat_B[43][1] +
                mat_A[217][2] * mat_B[51][1] +
                mat_A[217][3] * mat_B[59][1] +
                mat_A[218][0] * mat_B[67][1] +
                mat_A[218][1] * mat_B[75][1] +
                mat_A[218][2] * mat_B[83][1] +
                mat_A[218][3] * mat_B[91][1] +
                mat_A[219][0] * mat_B[99][1] +
                mat_A[219][1] * mat_B[107][1] +
                mat_A[219][2] * mat_B[115][1] +
                mat_A[219][3] * mat_B[123][1] +
                mat_A[220][0] * mat_B[131][1] +
                mat_A[220][1] * mat_B[139][1] +
                mat_A[220][2] * mat_B[147][1] +
                mat_A[220][3] * mat_B[155][1] +
                mat_A[221][0] * mat_B[163][1] +
                mat_A[221][1] * mat_B[171][1] +
                mat_A[221][2] * mat_B[179][1] +
                mat_A[221][3] * mat_B[187][1] +
                mat_A[222][0] * mat_B[195][1] +
                mat_A[222][1] * mat_B[203][1] +
                mat_A[222][2] * mat_B[211][1] +
                mat_A[222][3] * mat_B[219][1] +
                mat_A[223][0] * mat_B[227][1] +
                mat_A[223][1] * mat_B[235][1] +
                mat_A[223][2] * mat_B[243][1] +
                mat_A[223][3] * mat_B[251][1];
    mat_C[219][2] <=
                mat_A[216][0] * mat_B[3][2] +
                mat_A[216][1] * mat_B[11][2] +
                mat_A[216][2] * mat_B[19][2] +
                mat_A[216][3] * mat_B[27][2] +
                mat_A[217][0] * mat_B[35][2] +
                mat_A[217][1] * mat_B[43][2] +
                mat_A[217][2] * mat_B[51][2] +
                mat_A[217][3] * mat_B[59][2] +
                mat_A[218][0] * mat_B[67][2] +
                mat_A[218][1] * mat_B[75][2] +
                mat_A[218][2] * mat_B[83][2] +
                mat_A[218][3] * mat_B[91][2] +
                mat_A[219][0] * mat_B[99][2] +
                mat_A[219][1] * mat_B[107][2] +
                mat_A[219][2] * mat_B[115][2] +
                mat_A[219][3] * mat_B[123][2] +
                mat_A[220][0] * mat_B[131][2] +
                mat_A[220][1] * mat_B[139][2] +
                mat_A[220][2] * mat_B[147][2] +
                mat_A[220][3] * mat_B[155][2] +
                mat_A[221][0] * mat_B[163][2] +
                mat_A[221][1] * mat_B[171][2] +
                mat_A[221][2] * mat_B[179][2] +
                mat_A[221][3] * mat_B[187][2] +
                mat_A[222][0] * mat_B[195][2] +
                mat_A[222][1] * mat_B[203][2] +
                mat_A[222][2] * mat_B[211][2] +
                mat_A[222][3] * mat_B[219][2] +
                mat_A[223][0] * mat_B[227][2] +
                mat_A[223][1] * mat_B[235][2] +
                mat_A[223][2] * mat_B[243][2] +
                mat_A[223][3] * mat_B[251][2];
    mat_C[219][3] <=
                mat_A[216][0] * mat_B[3][3] +
                mat_A[216][1] * mat_B[11][3] +
                mat_A[216][2] * mat_B[19][3] +
                mat_A[216][3] * mat_B[27][3] +
                mat_A[217][0] * mat_B[35][3] +
                mat_A[217][1] * mat_B[43][3] +
                mat_A[217][2] * mat_B[51][3] +
                mat_A[217][3] * mat_B[59][3] +
                mat_A[218][0] * mat_B[67][3] +
                mat_A[218][1] * mat_B[75][3] +
                mat_A[218][2] * mat_B[83][3] +
                mat_A[218][3] * mat_B[91][3] +
                mat_A[219][0] * mat_B[99][3] +
                mat_A[219][1] * mat_B[107][3] +
                mat_A[219][2] * mat_B[115][3] +
                mat_A[219][3] * mat_B[123][3] +
                mat_A[220][0] * mat_B[131][3] +
                mat_A[220][1] * mat_B[139][3] +
                mat_A[220][2] * mat_B[147][3] +
                mat_A[220][3] * mat_B[155][3] +
                mat_A[221][0] * mat_B[163][3] +
                mat_A[221][1] * mat_B[171][3] +
                mat_A[221][2] * mat_B[179][3] +
                mat_A[221][3] * mat_B[187][3] +
                mat_A[222][0] * mat_B[195][3] +
                mat_A[222][1] * mat_B[203][3] +
                mat_A[222][2] * mat_B[211][3] +
                mat_A[222][3] * mat_B[219][3] +
                mat_A[223][0] * mat_B[227][3] +
                mat_A[223][1] * mat_B[235][3] +
                mat_A[223][2] * mat_B[243][3] +
                mat_A[223][3] * mat_B[251][3];
    mat_C[220][0] <=
                mat_A[216][0] * mat_B[4][0] +
                mat_A[216][1] * mat_B[12][0] +
                mat_A[216][2] * mat_B[20][0] +
                mat_A[216][3] * mat_B[28][0] +
                mat_A[217][0] * mat_B[36][0] +
                mat_A[217][1] * mat_B[44][0] +
                mat_A[217][2] * mat_B[52][0] +
                mat_A[217][3] * mat_B[60][0] +
                mat_A[218][0] * mat_B[68][0] +
                mat_A[218][1] * mat_B[76][0] +
                mat_A[218][2] * mat_B[84][0] +
                mat_A[218][3] * mat_B[92][0] +
                mat_A[219][0] * mat_B[100][0] +
                mat_A[219][1] * mat_B[108][0] +
                mat_A[219][2] * mat_B[116][0] +
                mat_A[219][3] * mat_B[124][0] +
                mat_A[220][0] * mat_B[132][0] +
                mat_A[220][1] * mat_B[140][0] +
                mat_A[220][2] * mat_B[148][0] +
                mat_A[220][3] * mat_B[156][0] +
                mat_A[221][0] * mat_B[164][0] +
                mat_A[221][1] * mat_B[172][0] +
                mat_A[221][2] * mat_B[180][0] +
                mat_A[221][3] * mat_B[188][0] +
                mat_A[222][0] * mat_B[196][0] +
                mat_A[222][1] * mat_B[204][0] +
                mat_A[222][2] * mat_B[212][0] +
                mat_A[222][3] * mat_B[220][0] +
                mat_A[223][0] * mat_B[228][0] +
                mat_A[223][1] * mat_B[236][0] +
                mat_A[223][2] * mat_B[244][0] +
                mat_A[223][3] * mat_B[252][0];
    mat_C[220][1] <=
                mat_A[216][0] * mat_B[4][1] +
                mat_A[216][1] * mat_B[12][1] +
                mat_A[216][2] * mat_B[20][1] +
                mat_A[216][3] * mat_B[28][1] +
                mat_A[217][0] * mat_B[36][1] +
                mat_A[217][1] * mat_B[44][1] +
                mat_A[217][2] * mat_B[52][1] +
                mat_A[217][3] * mat_B[60][1] +
                mat_A[218][0] * mat_B[68][1] +
                mat_A[218][1] * mat_B[76][1] +
                mat_A[218][2] * mat_B[84][1] +
                mat_A[218][3] * mat_B[92][1] +
                mat_A[219][0] * mat_B[100][1] +
                mat_A[219][1] * mat_B[108][1] +
                mat_A[219][2] * mat_B[116][1] +
                mat_A[219][3] * mat_B[124][1] +
                mat_A[220][0] * mat_B[132][1] +
                mat_A[220][1] * mat_B[140][1] +
                mat_A[220][2] * mat_B[148][1] +
                mat_A[220][3] * mat_B[156][1] +
                mat_A[221][0] * mat_B[164][1] +
                mat_A[221][1] * mat_B[172][1] +
                mat_A[221][2] * mat_B[180][1] +
                mat_A[221][3] * mat_B[188][1] +
                mat_A[222][0] * mat_B[196][1] +
                mat_A[222][1] * mat_B[204][1] +
                mat_A[222][2] * mat_B[212][1] +
                mat_A[222][3] * mat_B[220][1] +
                mat_A[223][0] * mat_B[228][1] +
                mat_A[223][1] * mat_B[236][1] +
                mat_A[223][2] * mat_B[244][1] +
                mat_A[223][3] * mat_B[252][1];
    mat_C[220][2] <=
                mat_A[216][0] * mat_B[4][2] +
                mat_A[216][1] * mat_B[12][2] +
                mat_A[216][2] * mat_B[20][2] +
                mat_A[216][3] * mat_B[28][2] +
                mat_A[217][0] * mat_B[36][2] +
                mat_A[217][1] * mat_B[44][2] +
                mat_A[217][2] * mat_B[52][2] +
                mat_A[217][3] * mat_B[60][2] +
                mat_A[218][0] * mat_B[68][2] +
                mat_A[218][1] * mat_B[76][2] +
                mat_A[218][2] * mat_B[84][2] +
                mat_A[218][3] * mat_B[92][2] +
                mat_A[219][0] * mat_B[100][2] +
                mat_A[219][1] * mat_B[108][2] +
                mat_A[219][2] * mat_B[116][2] +
                mat_A[219][3] * mat_B[124][2] +
                mat_A[220][0] * mat_B[132][2] +
                mat_A[220][1] * mat_B[140][2] +
                mat_A[220][2] * mat_B[148][2] +
                mat_A[220][3] * mat_B[156][2] +
                mat_A[221][0] * mat_B[164][2] +
                mat_A[221][1] * mat_B[172][2] +
                mat_A[221][2] * mat_B[180][2] +
                mat_A[221][3] * mat_B[188][2] +
                mat_A[222][0] * mat_B[196][2] +
                mat_A[222][1] * mat_B[204][2] +
                mat_A[222][2] * mat_B[212][2] +
                mat_A[222][3] * mat_B[220][2] +
                mat_A[223][0] * mat_B[228][2] +
                mat_A[223][1] * mat_B[236][2] +
                mat_A[223][2] * mat_B[244][2] +
                mat_A[223][3] * mat_B[252][2];
    mat_C[220][3] <=
                mat_A[216][0] * mat_B[4][3] +
                mat_A[216][1] * mat_B[12][3] +
                mat_A[216][2] * mat_B[20][3] +
                mat_A[216][3] * mat_B[28][3] +
                mat_A[217][0] * mat_B[36][3] +
                mat_A[217][1] * mat_B[44][3] +
                mat_A[217][2] * mat_B[52][3] +
                mat_A[217][3] * mat_B[60][3] +
                mat_A[218][0] * mat_B[68][3] +
                mat_A[218][1] * mat_B[76][3] +
                mat_A[218][2] * mat_B[84][3] +
                mat_A[218][3] * mat_B[92][3] +
                mat_A[219][0] * mat_B[100][3] +
                mat_A[219][1] * mat_B[108][3] +
                mat_A[219][2] * mat_B[116][3] +
                mat_A[219][3] * mat_B[124][3] +
                mat_A[220][0] * mat_B[132][3] +
                mat_A[220][1] * mat_B[140][3] +
                mat_A[220][2] * mat_B[148][3] +
                mat_A[220][3] * mat_B[156][3] +
                mat_A[221][0] * mat_B[164][3] +
                mat_A[221][1] * mat_B[172][3] +
                mat_A[221][2] * mat_B[180][3] +
                mat_A[221][3] * mat_B[188][3] +
                mat_A[222][0] * mat_B[196][3] +
                mat_A[222][1] * mat_B[204][3] +
                mat_A[222][2] * mat_B[212][3] +
                mat_A[222][3] * mat_B[220][3] +
                mat_A[223][0] * mat_B[228][3] +
                mat_A[223][1] * mat_B[236][3] +
                mat_A[223][2] * mat_B[244][3] +
                mat_A[223][3] * mat_B[252][3];
    mat_C[221][0] <=
                mat_A[216][0] * mat_B[5][0] +
                mat_A[216][1] * mat_B[13][0] +
                mat_A[216][2] * mat_B[21][0] +
                mat_A[216][3] * mat_B[29][0] +
                mat_A[217][0] * mat_B[37][0] +
                mat_A[217][1] * mat_B[45][0] +
                mat_A[217][2] * mat_B[53][0] +
                mat_A[217][3] * mat_B[61][0] +
                mat_A[218][0] * mat_B[69][0] +
                mat_A[218][1] * mat_B[77][0] +
                mat_A[218][2] * mat_B[85][0] +
                mat_A[218][3] * mat_B[93][0] +
                mat_A[219][0] * mat_B[101][0] +
                mat_A[219][1] * mat_B[109][0] +
                mat_A[219][2] * mat_B[117][0] +
                mat_A[219][3] * mat_B[125][0] +
                mat_A[220][0] * mat_B[133][0] +
                mat_A[220][1] * mat_B[141][0] +
                mat_A[220][2] * mat_B[149][0] +
                mat_A[220][3] * mat_B[157][0] +
                mat_A[221][0] * mat_B[165][0] +
                mat_A[221][1] * mat_B[173][0] +
                mat_A[221][2] * mat_B[181][0] +
                mat_A[221][3] * mat_B[189][0] +
                mat_A[222][0] * mat_B[197][0] +
                mat_A[222][1] * mat_B[205][0] +
                mat_A[222][2] * mat_B[213][0] +
                mat_A[222][3] * mat_B[221][0] +
                mat_A[223][0] * mat_B[229][0] +
                mat_A[223][1] * mat_B[237][0] +
                mat_A[223][2] * mat_B[245][0] +
                mat_A[223][3] * mat_B[253][0];
    mat_C[221][1] <=
                mat_A[216][0] * mat_B[5][1] +
                mat_A[216][1] * mat_B[13][1] +
                mat_A[216][2] * mat_B[21][1] +
                mat_A[216][3] * mat_B[29][1] +
                mat_A[217][0] * mat_B[37][1] +
                mat_A[217][1] * mat_B[45][1] +
                mat_A[217][2] * mat_B[53][1] +
                mat_A[217][3] * mat_B[61][1] +
                mat_A[218][0] * mat_B[69][1] +
                mat_A[218][1] * mat_B[77][1] +
                mat_A[218][2] * mat_B[85][1] +
                mat_A[218][3] * mat_B[93][1] +
                mat_A[219][0] * mat_B[101][1] +
                mat_A[219][1] * mat_B[109][1] +
                mat_A[219][2] * mat_B[117][1] +
                mat_A[219][3] * mat_B[125][1] +
                mat_A[220][0] * mat_B[133][1] +
                mat_A[220][1] * mat_B[141][1] +
                mat_A[220][2] * mat_B[149][1] +
                mat_A[220][3] * mat_B[157][1] +
                mat_A[221][0] * mat_B[165][1] +
                mat_A[221][1] * mat_B[173][1] +
                mat_A[221][2] * mat_B[181][1] +
                mat_A[221][3] * mat_B[189][1] +
                mat_A[222][0] * mat_B[197][1] +
                mat_A[222][1] * mat_B[205][1] +
                mat_A[222][2] * mat_B[213][1] +
                mat_A[222][3] * mat_B[221][1] +
                mat_A[223][0] * mat_B[229][1] +
                mat_A[223][1] * mat_B[237][1] +
                mat_A[223][2] * mat_B[245][1] +
                mat_A[223][3] * mat_B[253][1];
    mat_C[221][2] <=
                mat_A[216][0] * mat_B[5][2] +
                mat_A[216][1] * mat_B[13][2] +
                mat_A[216][2] * mat_B[21][2] +
                mat_A[216][3] * mat_B[29][2] +
                mat_A[217][0] * mat_B[37][2] +
                mat_A[217][1] * mat_B[45][2] +
                mat_A[217][2] * mat_B[53][2] +
                mat_A[217][3] * mat_B[61][2] +
                mat_A[218][0] * mat_B[69][2] +
                mat_A[218][1] * mat_B[77][2] +
                mat_A[218][2] * mat_B[85][2] +
                mat_A[218][3] * mat_B[93][2] +
                mat_A[219][0] * mat_B[101][2] +
                mat_A[219][1] * mat_B[109][2] +
                mat_A[219][2] * mat_B[117][2] +
                mat_A[219][3] * mat_B[125][2] +
                mat_A[220][0] * mat_B[133][2] +
                mat_A[220][1] * mat_B[141][2] +
                mat_A[220][2] * mat_B[149][2] +
                mat_A[220][3] * mat_B[157][2] +
                mat_A[221][0] * mat_B[165][2] +
                mat_A[221][1] * mat_B[173][2] +
                mat_A[221][2] * mat_B[181][2] +
                mat_A[221][3] * mat_B[189][2] +
                mat_A[222][0] * mat_B[197][2] +
                mat_A[222][1] * mat_B[205][2] +
                mat_A[222][2] * mat_B[213][2] +
                mat_A[222][3] * mat_B[221][2] +
                mat_A[223][0] * mat_B[229][2] +
                mat_A[223][1] * mat_B[237][2] +
                mat_A[223][2] * mat_B[245][2] +
                mat_A[223][3] * mat_B[253][2];
    mat_C[221][3] <=
                mat_A[216][0] * mat_B[5][3] +
                mat_A[216][1] * mat_B[13][3] +
                mat_A[216][2] * mat_B[21][3] +
                mat_A[216][3] * mat_B[29][3] +
                mat_A[217][0] * mat_B[37][3] +
                mat_A[217][1] * mat_B[45][3] +
                mat_A[217][2] * mat_B[53][3] +
                mat_A[217][3] * mat_B[61][3] +
                mat_A[218][0] * mat_B[69][3] +
                mat_A[218][1] * mat_B[77][3] +
                mat_A[218][2] * mat_B[85][3] +
                mat_A[218][3] * mat_B[93][3] +
                mat_A[219][0] * mat_B[101][3] +
                mat_A[219][1] * mat_B[109][3] +
                mat_A[219][2] * mat_B[117][3] +
                mat_A[219][3] * mat_B[125][3] +
                mat_A[220][0] * mat_B[133][3] +
                mat_A[220][1] * mat_B[141][3] +
                mat_A[220][2] * mat_B[149][3] +
                mat_A[220][3] * mat_B[157][3] +
                mat_A[221][0] * mat_B[165][3] +
                mat_A[221][1] * mat_B[173][3] +
                mat_A[221][2] * mat_B[181][3] +
                mat_A[221][3] * mat_B[189][3] +
                mat_A[222][0] * mat_B[197][3] +
                mat_A[222][1] * mat_B[205][3] +
                mat_A[222][2] * mat_B[213][3] +
                mat_A[222][3] * mat_B[221][3] +
                mat_A[223][0] * mat_B[229][3] +
                mat_A[223][1] * mat_B[237][3] +
                mat_A[223][2] * mat_B[245][3] +
                mat_A[223][3] * mat_B[253][3];
    mat_C[222][0] <=
                mat_A[216][0] * mat_B[6][0] +
                mat_A[216][1] * mat_B[14][0] +
                mat_A[216][2] * mat_B[22][0] +
                mat_A[216][3] * mat_B[30][0] +
                mat_A[217][0] * mat_B[38][0] +
                mat_A[217][1] * mat_B[46][0] +
                mat_A[217][2] * mat_B[54][0] +
                mat_A[217][3] * mat_B[62][0] +
                mat_A[218][0] * mat_B[70][0] +
                mat_A[218][1] * mat_B[78][0] +
                mat_A[218][2] * mat_B[86][0] +
                mat_A[218][3] * mat_B[94][0] +
                mat_A[219][0] * mat_B[102][0] +
                mat_A[219][1] * mat_B[110][0] +
                mat_A[219][2] * mat_B[118][0] +
                mat_A[219][3] * mat_B[126][0] +
                mat_A[220][0] * mat_B[134][0] +
                mat_A[220][1] * mat_B[142][0] +
                mat_A[220][2] * mat_B[150][0] +
                mat_A[220][3] * mat_B[158][0] +
                mat_A[221][0] * mat_B[166][0] +
                mat_A[221][1] * mat_B[174][0] +
                mat_A[221][2] * mat_B[182][0] +
                mat_A[221][3] * mat_B[190][0] +
                mat_A[222][0] * mat_B[198][0] +
                mat_A[222][1] * mat_B[206][0] +
                mat_A[222][2] * mat_B[214][0] +
                mat_A[222][3] * mat_B[222][0] +
                mat_A[223][0] * mat_B[230][0] +
                mat_A[223][1] * mat_B[238][0] +
                mat_A[223][2] * mat_B[246][0] +
                mat_A[223][3] * mat_B[254][0];
    mat_C[222][1] <=
                mat_A[216][0] * mat_B[6][1] +
                mat_A[216][1] * mat_B[14][1] +
                mat_A[216][2] * mat_B[22][1] +
                mat_A[216][3] * mat_B[30][1] +
                mat_A[217][0] * mat_B[38][1] +
                mat_A[217][1] * mat_B[46][1] +
                mat_A[217][2] * mat_B[54][1] +
                mat_A[217][3] * mat_B[62][1] +
                mat_A[218][0] * mat_B[70][1] +
                mat_A[218][1] * mat_B[78][1] +
                mat_A[218][2] * mat_B[86][1] +
                mat_A[218][3] * mat_B[94][1] +
                mat_A[219][0] * mat_B[102][1] +
                mat_A[219][1] * mat_B[110][1] +
                mat_A[219][2] * mat_B[118][1] +
                mat_A[219][3] * mat_B[126][1] +
                mat_A[220][0] * mat_B[134][1] +
                mat_A[220][1] * mat_B[142][1] +
                mat_A[220][2] * mat_B[150][1] +
                mat_A[220][3] * mat_B[158][1] +
                mat_A[221][0] * mat_B[166][1] +
                mat_A[221][1] * mat_B[174][1] +
                mat_A[221][2] * mat_B[182][1] +
                mat_A[221][3] * mat_B[190][1] +
                mat_A[222][0] * mat_B[198][1] +
                mat_A[222][1] * mat_B[206][1] +
                mat_A[222][2] * mat_B[214][1] +
                mat_A[222][3] * mat_B[222][1] +
                mat_A[223][0] * mat_B[230][1] +
                mat_A[223][1] * mat_B[238][1] +
                mat_A[223][2] * mat_B[246][1] +
                mat_A[223][3] * mat_B[254][1];
    mat_C[222][2] <=
                mat_A[216][0] * mat_B[6][2] +
                mat_A[216][1] * mat_B[14][2] +
                mat_A[216][2] * mat_B[22][2] +
                mat_A[216][3] * mat_B[30][2] +
                mat_A[217][0] * mat_B[38][2] +
                mat_A[217][1] * mat_B[46][2] +
                mat_A[217][2] * mat_B[54][2] +
                mat_A[217][3] * mat_B[62][2] +
                mat_A[218][0] * mat_B[70][2] +
                mat_A[218][1] * mat_B[78][2] +
                mat_A[218][2] * mat_B[86][2] +
                mat_A[218][3] * mat_B[94][2] +
                mat_A[219][0] * mat_B[102][2] +
                mat_A[219][1] * mat_B[110][2] +
                mat_A[219][2] * mat_B[118][2] +
                mat_A[219][3] * mat_B[126][2] +
                mat_A[220][0] * mat_B[134][2] +
                mat_A[220][1] * mat_B[142][2] +
                mat_A[220][2] * mat_B[150][2] +
                mat_A[220][3] * mat_B[158][2] +
                mat_A[221][0] * mat_B[166][2] +
                mat_A[221][1] * mat_B[174][2] +
                mat_A[221][2] * mat_B[182][2] +
                mat_A[221][3] * mat_B[190][2] +
                mat_A[222][0] * mat_B[198][2] +
                mat_A[222][1] * mat_B[206][2] +
                mat_A[222][2] * mat_B[214][2] +
                mat_A[222][3] * mat_B[222][2] +
                mat_A[223][0] * mat_B[230][2] +
                mat_A[223][1] * mat_B[238][2] +
                mat_A[223][2] * mat_B[246][2] +
                mat_A[223][3] * mat_B[254][2];
    mat_C[222][3] <=
                mat_A[216][0] * mat_B[6][3] +
                mat_A[216][1] * mat_B[14][3] +
                mat_A[216][2] * mat_B[22][3] +
                mat_A[216][3] * mat_B[30][3] +
                mat_A[217][0] * mat_B[38][3] +
                mat_A[217][1] * mat_B[46][3] +
                mat_A[217][2] * mat_B[54][3] +
                mat_A[217][3] * mat_B[62][3] +
                mat_A[218][0] * mat_B[70][3] +
                mat_A[218][1] * mat_B[78][3] +
                mat_A[218][2] * mat_B[86][3] +
                mat_A[218][3] * mat_B[94][3] +
                mat_A[219][0] * mat_B[102][3] +
                mat_A[219][1] * mat_B[110][3] +
                mat_A[219][2] * mat_B[118][3] +
                mat_A[219][3] * mat_B[126][3] +
                mat_A[220][0] * mat_B[134][3] +
                mat_A[220][1] * mat_B[142][3] +
                mat_A[220][2] * mat_B[150][3] +
                mat_A[220][3] * mat_B[158][3] +
                mat_A[221][0] * mat_B[166][3] +
                mat_A[221][1] * mat_B[174][3] +
                mat_A[221][2] * mat_B[182][3] +
                mat_A[221][3] * mat_B[190][3] +
                mat_A[222][0] * mat_B[198][3] +
                mat_A[222][1] * mat_B[206][3] +
                mat_A[222][2] * mat_B[214][3] +
                mat_A[222][3] * mat_B[222][3] +
                mat_A[223][0] * mat_B[230][3] +
                mat_A[223][1] * mat_B[238][3] +
                mat_A[223][2] * mat_B[246][3] +
                mat_A[223][3] * mat_B[254][3];
    mat_C[223][0] <=
                mat_A[216][0] * mat_B[7][0] +
                mat_A[216][1] * mat_B[15][0] +
                mat_A[216][2] * mat_B[23][0] +
                mat_A[216][3] * mat_B[31][0] +
                mat_A[217][0] * mat_B[39][0] +
                mat_A[217][1] * mat_B[47][0] +
                mat_A[217][2] * mat_B[55][0] +
                mat_A[217][3] * mat_B[63][0] +
                mat_A[218][0] * mat_B[71][0] +
                mat_A[218][1] * mat_B[79][0] +
                mat_A[218][2] * mat_B[87][0] +
                mat_A[218][3] * mat_B[95][0] +
                mat_A[219][0] * mat_B[103][0] +
                mat_A[219][1] * mat_B[111][0] +
                mat_A[219][2] * mat_B[119][0] +
                mat_A[219][3] * mat_B[127][0] +
                mat_A[220][0] * mat_B[135][0] +
                mat_A[220][1] * mat_B[143][0] +
                mat_A[220][2] * mat_B[151][0] +
                mat_A[220][3] * mat_B[159][0] +
                mat_A[221][0] * mat_B[167][0] +
                mat_A[221][1] * mat_B[175][0] +
                mat_A[221][2] * mat_B[183][0] +
                mat_A[221][3] * mat_B[191][0] +
                mat_A[222][0] * mat_B[199][0] +
                mat_A[222][1] * mat_B[207][0] +
                mat_A[222][2] * mat_B[215][0] +
                mat_A[222][3] * mat_B[223][0] +
                mat_A[223][0] * mat_B[231][0] +
                mat_A[223][1] * mat_B[239][0] +
                mat_A[223][2] * mat_B[247][0] +
                mat_A[223][3] * mat_B[255][0];
    mat_C[223][1] <=
                mat_A[216][0] * mat_B[7][1] +
                mat_A[216][1] * mat_B[15][1] +
                mat_A[216][2] * mat_B[23][1] +
                mat_A[216][3] * mat_B[31][1] +
                mat_A[217][0] * mat_B[39][1] +
                mat_A[217][1] * mat_B[47][1] +
                mat_A[217][2] * mat_B[55][1] +
                mat_A[217][3] * mat_B[63][1] +
                mat_A[218][0] * mat_B[71][1] +
                mat_A[218][1] * mat_B[79][1] +
                mat_A[218][2] * mat_B[87][1] +
                mat_A[218][3] * mat_B[95][1] +
                mat_A[219][0] * mat_B[103][1] +
                mat_A[219][1] * mat_B[111][1] +
                mat_A[219][2] * mat_B[119][1] +
                mat_A[219][3] * mat_B[127][1] +
                mat_A[220][0] * mat_B[135][1] +
                mat_A[220][1] * mat_B[143][1] +
                mat_A[220][2] * mat_B[151][1] +
                mat_A[220][3] * mat_B[159][1] +
                mat_A[221][0] * mat_B[167][1] +
                mat_A[221][1] * mat_B[175][1] +
                mat_A[221][2] * mat_B[183][1] +
                mat_A[221][3] * mat_B[191][1] +
                mat_A[222][0] * mat_B[199][1] +
                mat_A[222][1] * mat_B[207][1] +
                mat_A[222][2] * mat_B[215][1] +
                mat_A[222][3] * mat_B[223][1] +
                mat_A[223][0] * mat_B[231][1] +
                mat_A[223][1] * mat_B[239][1] +
                mat_A[223][2] * mat_B[247][1] +
                mat_A[223][3] * mat_B[255][1];
    mat_C[223][2] <=
                mat_A[216][0] * mat_B[7][2] +
                mat_A[216][1] * mat_B[15][2] +
                mat_A[216][2] * mat_B[23][2] +
                mat_A[216][3] * mat_B[31][2] +
                mat_A[217][0] * mat_B[39][2] +
                mat_A[217][1] * mat_B[47][2] +
                mat_A[217][2] * mat_B[55][2] +
                mat_A[217][3] * mat_B[63][2] +
                mat_A[218][0] * mat_B[71][2] +
                mat_A[218][1] * mat_B[79][2] +
                mat_A[218][2] * mat_B[87][2] +
                mat_A[218][3] * mat_B[95][2] +
                mat_A[219][0] * mat_B[103][2] +
                mat_A[219][1] * mat_B[111][2] +
                mat_A[219][2] * mat_B[119][2] +
                mat_A[219][3] * mat_B[127][2] +
                mat_A[220][0] * mat_B[135][2] +
                mat_A[220][1] * mat_B[143][2] +
                mat_A[220][2] * mat_B[151][2] +
                mat_A[220][3] * mat_B[159][2] +
                mat_A[221][0] * mat_B[167][2] +
                mat_A[221][1] * mat_B[175][2] +
                mat_A[221][2] * mat_B[183][2] +
                mat_A[221][3] * mat_B[191][2] +
                mat_A[222][0] * mat_B[199][2] +
                mat_A[222][1] * mat_B[207][2] +
                mat_A[222][2] * mat_B[215][2] +
                mat_A[222][3] * mat_B[223][2] +
                mat_A[223][0] * mat_B[231][2] +
                mat_A[223][1] * mat_B[239][2] +
                mat_A[223][2] * mat_B[247][2] +
                mat_A[223][3] * mat_B[255][2];
    mat_C[223][3] <=
                mat_A[216][0] * mat_B[7][3] +
                mat_A[216][1] * mat_B[15][3] +
                mat_A[216][2] * mat_B[23][3] +
                mat_A[216][3] * mat_B[31][3] +
                mat_A[217][0] * mat_B[39][3] +
                mat_A[217][1] * mat_B[47][3] +
                mat_A[217][2] * mat_B[55][3] +
                mat_A[217][3] * mat_B[63][3] +
                mat_A[218][0] * mat_B[71][3] +
                mat_A[218][1] * mat_B[79][3] +
                mat_A[218][2] * mat_B[87][3] +
                mat_A[218][3] * mat_B[95][3] +
                mat_A[219][0] * mat_B[103][3] +
                mat_A[219][1] * mat_B[111][3] +
                mat_A[219][2] * mat_B[119][3] +
                mat_A[219][3] * mat_B[127][3] +
                mat_A[220][0] * mat_B[135][3] +
                mat_A[220][1] * mat_B[143][3] +
                mat_A[220][2] * mat_B[151][3] +
                mat_A[220][3] * mat_B[159][3] +
                mat_A[221][0] * mat_B[167][3] +
                mat_A[221][1] * mat_B[175][3] +
                mat_A[221][2] * mat_B[183][3] +
                mat_A[221][3] * mat_B[191][3] +
                mat_A[222][0] * mat_B[199][3] +
                mat_A[222][1] * mat_B[207][3] +
                mat_A[222][2] * mat_B[215][3] +
                mat_A[222][3] * mat_B[223][3] +
                mat_A[223][0] * mat_B[231][3] +
                mat_A[223][1] * mat_B[239][3] +
                mat_A[223][2] * mat_B[247][3] +
                mat_A[223][3] * mat_B[255][3];
    mat_C[224][0] <=
                mat_A[224][0] * mat_B[0][0] +
                mat_A[224][1] * mat_B[8][0] +
                mat_A[224][2] * mat_B[16][0] +
                mat_A[224][3] * mat_B[24][0] +
                mat_A[225][0] * mat_B[32][0] +
                mat_A[225][1] * mat_B[40][0] +
                mat_A[225][2] * mat_B[48][0] +
                mat_A[225][3] * mat_B[56][0] +
                mat_A[226][0] * mat_B[64][0] +
                mat_A[226][1] * mat_B[72][0] +
                mat_A[226][2] * mat_B[80][0] +
                mat_A[226][3] * mat_B[88][0] +
                mat_A[227][0] * mat_B[96][0] +
                mat_A[227][1] * mat_B[104][0] +
                mat_A[227][2] * mat_B[112][0] +
                mat_A[227][3] * mat_B[120][0] +
                mat_A[228][0] * mat_B[128][0] +
                mat_A[228][1] * mat_B[136][0] +
                mat_A[228][2] * mat_B[144][0] +
                mat_A[228][3] * mat_B[152][0] +
                mat_A[229][0] * mat_B[160][0] +
                mat_A[229][1] * mat_B[168][0] +
                mat_A[229][2] * mat_B[176][0] +
                mat_A[229][3] * mat_B[184][0] +
                mat_A[230][0] * mat_B[192][0] +
                mat_A[230][1] * mat_B[200][0] +
                mat_A[230][2] * mat_B[208][0] +
                mat_A[230][3] * mat_B[216][0] +
                mat_A[231][0] * mat_B[224][0] +
                mat_A[231][1] * mat_B[232][0] +
                mat_A[231][2] * mat_B[240][0] +
                mat_A[231][3] * mat_B[248][0];
    mat_C[224][1] <=
                mat_A[224][0] * mat_B[0][1] +
                mat_A[224][1] * mat_B[8][1] +
                mat_A[224][2] * mat_B[16][1] +
                mat_A[224][3] * mat_B[24][1] +
                mat_A[225][0] * mat_B[32][1] +
                mat_A[225][1] * mat_B[40][1] +
                mat_A[225][2] * mat_B[48][1] +
                mat_A[225][3] * mat_B[56][1] +
                mat_A[226][0] * mat_B[64][1] +
                mat_A[226][1] * mat_B[72][1] +
                mat_A[226][2] * mat_B[80][1] +
                mat_A[226][3] * mat_B[88][1] +
                mat_A[227][0] * mat_B[96][1] +
                mat_A[227][1] * mat_B[104][1] +
                mat_A[227][2] * mat_B[112][1] +
                mat_A[227][3] * mat_B[120][1] +
                mat_A[228][0] * mat_B[128][1] +
                mat_A[228][1] * mat_B[136][1] +
                mat_A[228][2] * mat_B[144][1] +
                mat_A[228][3] * mat_B[152][1] +
                mat_A[229][0] * mat_B[160][1] +
                mat_A[229][1] * mat_B[168][1] +
                mat_A[229][2] * mat_B[176][1] +
                mat_A[229][3] * mat_B[184][1] +
                mat_A[230][0] * mat_B[192][1] +
                mat_A[230][1] * mat_B[200][1] +
                mat_A[230][2] * mat_B[208][1] +
                mat_A[230][3] * mat_B[216][1] +
                mat_A[231][0] * mat_B[224][1] +
                mat_A[231][1] * mat_B[232][1] +
                mat_A[231][2] * mat_B[240][1] +
                mat_A[231][3] * mat_B[248][1];
    mat_C[224][2] <=
                mat_A[224][0] * mat_B[0][2] +
                mat_A[224][1] * mat_B[8][2] +
                mat_A[224][2] * mat_B[16][2] +
                mat_A[224][3] * mat_B[24][2] +
                mat_A[225][0] * mat_B[32][2] +
                mat_A[225][1] * mat_B[40][2] +
                mat_A[225][2] * mat_B[48][2] +
                mat_A[225][3] * mat_B[56][2] +
                mat_A[226][0] * mat_B[64][2] +
                mat_A[226][1] * mat_B[72][2] +
                mat_A[226][2] * mat_B[80][2] +
                mat_A[226][3] * mat_B[88][2] +
                mat_A[227][0] * mat_B[96][2] +
                mat_A[227][1] * mat_B[104][2] +
                mat_A[227][2] * mat_B[112][2] +
                mat_A[227][3] * mat_B[120][2] +
                mat_A[228][0] * mat_B[128][2] +
                mat_A[228][1] * mat_B[136][2] +
                mat_A[228][2] * mat_B[144][2] +
                mat_A[228][3] * mat_B[152][2] +
                mat_A[229][0] * mat_B[160][2] +
                mat_A[229][1] * mat_B[168][2] +
                mat_A[229][2] * mat_B[176][2] +
                mat_A[229][3] * mat_B[184][2] +
                mat_A[230][0] * mat_B[192][2] +
                mat_A[230][1] * mat_B[200][2] +
                mat_A[230][2] * mat_B[208][2] +
                mat_A[230][3] * mat_B[216][2] +
                mat_A[231][0] * mat_B[224][2] +
                mat_A[231][1] * mat_B[232][2] +
                mat_A[231][2] * mat_B[240][2] +
                mat_A[231][3] * mat_B[248][2];
    mat_C[224][3] <=
                mat_A[224][0] * mat_B[0][3] +
                mat_A[224][1] * mat_B[8][3] +
                mat_A[224][2] * mat_B[16][3] +
                mat_A[224][3] * mat_B[24][3] +
                mat_A[225][0] * mat_B[32][3] +
                mat_A[225][1] * mat_B[40][3] +
                mat_A[225][2] * mat_B[48][3] +
                mat_A[225][3] * mat_B[56][3] +
                mat_A[226][0] * mat_B[64][3] +
                mat_A[226][1] * mat_B[72][3] +
                mat_A[226][2] * mat_B[80][3] +
                mat_A[226][3] * mat_B[88][3] +
                mat_A[227][0] * mat_B[96][3] +
                mat_A[227][1] * mat_B[104][3] +
                mat_A[227][2] * mat_B[112][3] +
                mat_A[227][3] * mat_B[120][3] +
                mat_A[228][0] * mat_B[128][3] +
                mat_A[228][1] * mat_B[136][3] +
                mat_A[228][2] * mat_B[144][3] +
                mat_A[228][3] * mat_B[152][3] +
                mat_A[229][0] * mat_B[160][3] +
                mat_A[229][1] * mat_B[168][3] +
                mat_A[229][2] * mat_B[176][3] +
                mat_A[229][3] * mat_B[184][3] +
                mat_A[230][0] * mat_B[192][3] +
                mat_A[230][1] * mat_B[200][3] +
                mat_A[230][2] * mat_B[208][3] +
                mat_A[230][3] * mat_B[216][3] +
                mat_A[231][0] * mat_B[224][3] +
                mat_A[231][1] * mat_B[232][3] +
                mat_A[231][2] * mat_B[240][3] +
                mat_A[231][3] * mat_B[248][3];
    mat_C[225][0] <=
                mat_A[224][0] * mat_B[1][0] +
                mat_A[224][1] * mat_B[9][0] +
                mat_A[224][2] * mat_B[17][0] +
                mat_A[224][3] * mat_B[25][0] +
                mat_A[225][0] * mat_B[33][0] +
                mat_A[225][1] * mat_B[41][0] +
                mat_A[225][2] * mat_B[49][0] +
                mat_A[225][3] * mat_B[57][0] +
                mat_A[226][0] * mat_B[65][0] +
                mat_A[226][1] * mat_B[73][0] +
                mat_A[226][2] * mat_B[81][0] +
                mat_A[226][3] * mat_B[89][0] +
                mat_A[227][0] * mat_B[97][0] +
                mat_A[227][1] * mat_B[105][0] +
                mat_A[227][2] * mat_B[113][0] +
                mat_A[227][3] * mat_B[121][0] +
                mat_A[228][0] * mat_B[129][0] +
                mat_A[228][1] * mat_B[137][0] +
                mat_A[228][2] * mat_B[145][0] +
                mat_A[228][3] * mat_B[153][0] +
                mat_A[229][0] * mat_B[161][0] +
                mat_A[229][1] * mat_B[169][0] +
                mat_A[229][2] * mat_B[177][0] +
                mat_A[229][3] * mat_B[185][0] +
                mat_A[230][0] * mat_B[193][0] +
                mat_A[230][1] * mat_B[201][0] +
                mat_A[230][2] * mat_B[209][0] +
                mat_A[230][3] * mat_B[217][0] +
                mat_A[231][0] * mat_B[225][0] +
                mat_A[231][1] * mat_B[233][0] +
                mat_A[231][2] * mat_B[241][0] +
                mat_A[231][3] * mat_B[249][0];
    mat_C[225][1] <=
                mat_A[224][0] * mat_B[1][1] +
                mat_A[224][1] * mat_B[9][1] +
                mat_A[224][2] * mat_B[17][1] +
                mat_A[224][3] * mat_B[25][1] +
                mat_A[225][0] * mat_B[33][1] +
                mat_A[225][1] * mat_B[41][1] +
                mat_A[225][2] * mat_B[49][1] +
                mat_A[225][3] * mat_B[57][1] +
                mat_A[226][0] * mat_B[65][1] +
                mat_A[226][1] * mat_B[73][1] +
                mat_A[226][2] * mat_B[81][1] +
                mat_A[226][3] * mat_B[89][1] +
                mat_A[227][0] * mat_B[97][1] +
                mat_A[227][1] * mat_B[105][1] +
                mat_A[227][2] * mat_B[113][1] +
                mat_A[227][3] * mat_B[121][1] +
                mat_A[228][0] * mat_B[129][1] +
                mat_A[228][1] * mat_B[137][1] +
                mat_A[228][2] * mat_B[145][1] +
                mat_A[228][3] * mat_B[153][1] +
                mat_A[229][0] * mat_B[161][1] +
                mat_A[229][1] * mat_B[169][1] +
                mat_A[229][2] * mat_B[177][1] +
                mat_A[229][3] * mat_B[185][1] +
                mat_A[230][0] * mat_B[193][1] +
                mat_A[230][1] * mat_B[201][1] +
                mat_A[230][2] * mat_B[209][1] +
                mat_A[230][3] * mat_B[217][1] +
                mat_A[231][0] * mat_B[225][1] +
                mat_A[231][1] * mat_B[233][1] +
                mat_A[231][2] * mat_B[241][1] +
                mat_A[231][3] * mat_B[249][1];
    mat_C[225][2] <=
                mat_A[224][0] * mat_B[1][2] +
                mat_A[224][1] * mat_B[9][2] +
                mat_A[224][2] * mat_B[17][2] +
                mat_A[224][3] * mat_B[25][2] +
                mat_A[225][0] * mat_B[33][2] +
                mat_A[225][1] * mat_B[41][2] +
                mat_A[225][2] * mat_B[49][2] +
                mat_A[225][3] * mat_B[57][2] +
                mat_A[226][0] * mat_B[65][2] +
                mat_A[226][1] * mat_B[73][2] +
                mat_A[226][2] * mat_B[81][2] +
                mat_A[226][3] * mat_B[89][2] +
                mat_A[227][0] * mat_B[97][2] +
                mat_A[227][1] * mat_B[105][2] +
                mat_A[227][2] * mat_B[113][2] +
                mat_A[227][3] * mat_B[121][2] +
                mat_A[228][0] * mat_B[129][2] +
                mat_A[228][1] * mat_B[137][2] +
                mat_A[228][2] * mat_B[145][2] +
                mat_A[228][3] * mat_B[153][2] +
                mat_A[229][0] * mat_B[161][2] +
                mat_A[229][1] * mat_B[169][2] +
                mat_A[229][2] * mat_B[177][2] +
                mat_A[229][3] * mat_B[185][2] +
                mat_A[230][0] * mat_B[193][2] +
                mat_A[230][1] * mat_B[201][2] +
                mat_A[230][2] * mat_B[209][2] +
                mat_A[230][3] * mat_B[217][2] +
                mat_A[231][0] * mat_B[225][2] +
                mat_A[231][1] * mat_B[233][2] +
                mat_A[231][2] * mat_B[241][2] +
                mat_A[231][3] * mat_B[249][2];
    mat_C[225][3] <=
                mat_A[224][0] * mat_B[1][3] +
                mat_A[224][1] * mat_B[9][3] +
                mat_A[224][2] * mat_B[17][3] +
                mat_A[224][3] * mat_B[25][3] +
                mat_A[225][0] * mat_B[33][3] +
                mat_A[225][1] * mat_B[41][3] +
                mat_A[225][2] * mat_B[49][3] +
                mat_A[225][3] * mat_B[57][3] +
                mat_A[226][0] * mat_B[65][3] +
                mat_A[226][1] * mat_B[73][3] +
                mat_A[226][2] * mat_B[81][3] +
                mat_A[226][3] * mat_B[89][3] +
                mat_A[227][0] * mat_B[97][3] +
                mat_A[227][1] * mat_B[105][3] +
                mat_A[227][2] * mat_B[113][3] +
                mat_A[227][3] * mat_B[121][3] +
                mat_A[228][0] * mat_B[129][3] +
                mat_A[228][1] * mat_B[137][3] +
                mat_A[228][2] * mat_B[145][3] +
                mat_A[228][3] * mat_B[153][3] +
                mat_A[229][0] * mat_B[161][3] +
                mat_A[229][1] * mat_B[169][3] +
                mat_A[229][2] * mat_B[177][3] +
                mat_A[229][3] * mat_B[185][3] +
                mat_A[230][0] * mat_B[193][3] +
                mat_A[230][1] * mat_B[201][3] +
                mat_A[230][2] * mat_B[209][3] +
                mat_A[230][3] * mat_B[217][3] +
                mat_A[231][0] * mat_B[225][3] +
                mat_A[231][1] * mat_B[233][3] +
                mat_A[231][2] * mat_B[241][3] +
                mat_A[231][3] * mat_B[249][3];
    mat_C[226][0] <=
                mat_A[224][0] * mat_B[2][0] +
                mat_A[224][1] * mat_B[10][0] +
                mat_A[224][2] * mat_B[18][0] +
                mat_A[224][3] * mat_B[26][0] +
                mat_A[225][0] * mat_B[34][0] +
                mat_A[225][1] * mat_B[42][0] +
                mat_A[225][2] * mat_B[50][0] +
                mat_A[225][3] * mat_B[58][0] +
                mat_A[226][0] * mat_B[66][0] +
                mat_A[226][1] * mat_B[74][0] +
                mat_A[226][2] * mat_B[82][0] +
                mat_A[226][3] * mat_B[90][0] +
                mat_A[227][0] * mat_B[98][0] +
                mat_A[227][1] * mat_B[106][0] +
                mat_A[227][2] * mat_B[114][0] +
                mat_A[227][3] * mat_B[122][0] +
                mat_A[228][0] * mat_B[130][0] +
                mat_A[228][1] * mat_B[138][0] +
                mat_A[228][2] * mat_B[146][0] +
                mat_A[228][3] * mat_B[154][0] +
                mat_A[229][0] * mat_B[162][0] +
                mat_A[229][1] * mat_B[170][0] +
                mat_A[229][2] * mat_B[178][0] +
                mat_A[229][3] * mat_B[186][0] +
                mat_A[230][0] * mat_B[194][0] +
                mat_A[230][1] * mat_B[202][0] +
                mat_A[230][2] * mat_B[210][0] +
                mat_A[230][3] * mat_B[218][0] +
                mat_A[231][0] * mat_B[226][0] +
                mat_A[231][1] * mat_B[234][0] +
                mat_A[231][2] * mat_B[242][0] +
                mat_A[231][3] * mat_B[250][0];
    mat_C[226][1] <=
                mat_A[224][0] * mat_B[2][1] +
                mat_A[224][1] * mat_B[10][1] +
                mat_A[224][2] * mat_B[18][1] +
                mat_A[224][3] * mat_B[26][1] +
                mat_A[225][0] * mat_B[34][1] +
                mat_A[225][1] * mat_B[42][1] +
                mat_A[225][2] * mat_B[50][1] +
                mat_A[225][3] * mat_B[58][1] +
                mat_A[226][0] * mat_B[66][1] +
                mat_A[226][1] * mat_B[74][1] +
                mat_A[226][2] * mat_B[82][1] +
                mat_A[226][3] * mat_B[90][1] +
                mat_A[227][0] * mat_B[98][1] +
                mat_A[227][1] * mat_B[106][1] +
                mat_A[227][2] * mat_B[114][1] +
                mat_A[227][3] * mat_B[122][1] +
                mat_A[228][0] * mat_B[130][1] +
                mat_A[228][1] * mat_B[138][1] +
                mat_A[228][2] * mat_B[146][1] +
                mat_A[228][3] * mat_B[154][1] +
                mat_A[229][0] * mat_B[162][1] +
                mat_A[229][1] * mat_B[170][1] +
                mat_A[229][2] * mat_B[178][1] +
                mat_A[229][3] * mat_B[186][1] +
                mat_A[230][0] * mat_B[194][1] +
                mat_A[230][1] * mat_B[202][1] +
                mat_A[230][2] * mat_B[210][1] +
                mat_A[230][3] * mat_B[218][1] +
                mat_A[231][0] * mat_B[226][1] +
                mat_A[231][1] * mat_B[234][1] +
                mat_A[231][2] * mat_B[242][1] +
                mat_A[231][3] * mat_B[250][1];
    mat_C[226][2] <=
                mat_A[224][0] * mat_B[2][2] +
                mat_A[224][1] * mat_B[10][2] +
                mat_A[224][2] * mat_B[18][2] +
                mat_A[224][3] * mat_B[26][2] +
                mat_A[225][0] * mat_B[34][2] +
                mat_A[225][1] * mat_B[42][2] +
                mat_A[225][2] * mat_B[50][2] +
                mat_A[225][3] * mat_B[58][2] +
                mat_A[226][0] * mat_B[66][2] +
                mat_A[226][1] * mat_B[74][2] +
                mat_A[226][2] * mat_B[82][2] +
                mat_A[226][3] * mat_B[90][2] +
                mat_A[227][0] * mat_B[98][2] +
                mat_A[227][1] * mat_B[106][2] +
                mat_A[227][2] * mat_B[114][2] +
                mat_A[227][3] * mat_B[122][2] +
                mat_A[228][0] * mat_B[130][2] +
                mat_A[228][1] * mat_B[138][2] +
                mat_A[228][2] * mat_B[146][2] +
                mat_A[228][3] * mat_B[154][2] +
                mat_A[229][0] * mat_B[162][2] +
                mat_A[229][1] * mat_B[170][2] +
                mat_A[229][2] * mat_B[178][2] +
                mat_A[229][3] * mat_B[186][2] +
                mat_A[230][0] * mat_B[194][2] +
                mat_A[230][1] * mat_B[202][2] +
                mat_A[230][2] * mat_B[210][2] +
                mat_A[230][3] * mat_B[218][2] +
                mat_A[231][0] * mat_B[226][2] +
                mat_A[231][1] * mat_B[234][2] +
                mat_A[231][2] * mat_B[242][2] +
                mat_A[231][3] * mat_B[250][2];
    mat_C[226][3] <=
                mat_A[224][0] * mat_B[2][3] +
                mat_A[224][1] * mat_B[10][3] +
                mat_A[224][2] * mat_B[18][3] +
                mat_A[224][3] * mat_B[26][3] +
                mat_A[225][0] * mat_B[34][3] +
                mat_A[225][1] * mat_B[42][3] +
                mat_A[225][2] * mat_B[50][3] +
                mat_A[225][3] * mat_B[58][3] +
                mat_A[226][0] * mat_B[66][3] +
                mat_A[226][1] * mat_B[74][3] +
                mat_A[226][2] * mat_B[82][3] +
                mat_A[226][3] * mat_B[90][3] +
                mat_A[227][0] * mat_B[98][3] +
                mat_A[227][1] * mat_B[106][3] +
                mat_A[227][2] * mat_B[114][3] +
                mat_A[227][3] * mat_B[122][3] +
                mat_A[228][0] * mat_B[130][3] +
                mat_A[228][1] * mat_B[138][3] +
                mat_A[228][2] * mat_B[146][3] +
                mat_A[228][3] * mat_B[154][3] +
                mat_A[229][0] * mat_B[162][3] +
                mat_A[229][1] * mat_B[170][3] +
                mat_A[229][2] * mat_B[178][3] +
                mat_A[229][3] * mat_B[186][3] +
                mat_A[230][0] * mat_B[194][3] +
                mat_A[230][1] * mat_B[202][3] +
                mat_A[230][2] * mat_B[210][3] +
                mat_A[230][3] * mat_B[218][3] +
                mat_A[231][0] * mat_B[226][3] +
                mat_A[231][1] * mat_B[234][3] +
                mat_A[231][2] * mat_B[242][3] +
                mat_A[231][3] * mat_B[250][3];
    mat_C[227][0] <=
                mat_A[224][0] * mat_B[3][0] +
                mat_A[224][1] * mat_B[11][0] +
                mat_A[224][2] * mat_B[19][0] +
                mat_A[224][3] * mat_B[27][0] +
                mat_A[225][0] * mat_B[35][0] +
                mat_A[225][1] * mat_B[43][0] +
                mat_A[225][2] * mat_B[51][0] +
                mat_A[225][3] * mat_B[59][0] +
                mat_A[226][0] * mat_B[67][0] +
                mat_A[226][1] * mat_B[75][0] +
                mat_A[226][2] * mat_B[83][0] +
                mat_A[226][3] * mat_B[91][0] +
                mat_A[227][0] * mat_B[99][0] +
                mat_A[227][1] * mat_B[107][0] +
                mat_A[227][2] * mat_B[115][0] +
                mat_A[227][3] * mat_B[123][0] +
                mat_A[228][0] * mat_B[131][0] +
                mat_A[228][1] * mat_B[139][0] +
                mat_A[228][2] * mat_B[147][0] +
                mat_A[228][3] * mat_B[155][0] +
                mat_A[229][0] * mat_B[163][0] +
                mat_A[229][1] * mat_B[171][0] +
                mat_A[229][2] * mat_B[179][0] +
                mat_A[229][3] * mat_B[187][0] +
                mat_A[230][0] * mat_B[195][0] +
                mat_A[230][1] * mat_B[203][0] +
                mat_A[230][2] * mat_B[211][0] +
                mat_A[230][3] * mat_B[219][0] +
                mat_A[231][0] * mat_B[227][0] +
                mat_A[231][1] * mat_B[235][0] +
                mat_A[231][2] * mat_B[243][0] +
                mat_A[231][3] * mat_B[251][0];
    mat_C[227][1] <=
                mat_A[224][0] * mat_B[3][1] +
                mat_A[224][1] * mat_B[11][1] +
                mat_A[224][2] * mat_B[19][1] +
                mat_A[224][3] * mat_B[27][1] +
                mat_A[225][0] * mat_B[35][1] +
                mat_A[225][1] * mat_B[43][1] +
                mat_A[225][2] * mat_B[51][1] +
                mat_A[225][3] * mat_B[59][1] +
                mat_A[226][0] * mat_B[67][1] +
                mat_A[226][1] * mat_B[75][1] +
                mat_A[226][2] * mat_B[83][1] +
                mat_A[226][3] * mat_B[91][1] +
                mat_A[227][0] * mat_B[99][1] +
                mat_A[227][1] * mat_B[107][1] +
                mat_A[227][2] * mat_B[115][1] +
                mat_A[227][3] * mat_B[123][1] +
                mat_A[228][0] * mat_B[131][1] +
                mat_A[228][1] * mat_B[139][1] +
                mat_A[228][2] * mat_B[147][1] +
                mat_A[228][3] * mat_B[155][1] +
                mat_A[229][0] * mat_B[163][1] +
                mat_A[229][1] * mat_B[171][1] +
                mat_A[229][2] * mat_B[179][1] +
                mat_A[229][3] * mat_B[187][1] +
                mat_A[230][0] * mat_B[195][1] +
                mat_A[230][1] * mat_B[203][1] +
                mat_A[230][2] * mat_B[211][1] +
                mat_A[230][3] * mat_B[219][1] +
                mat_A[231][0] * mat_B[227][1] +
                mat_A[231][1] * mat_B[235][1] +
                mat_A[231][2] * mat_B[243][1] +
                mat_A[231][3] * mat_B[251][1];
    mat_C[227][2] <=
                mat_A[224][0] * mat_B[3][2] +
                mat_A[224][1] * mat_B[11][2] +
                mat_A[224][2] * mat_B[19][2] +
                mat_A[224][3] * mat_B[27][2] +
                mat_A[225][0] * mat_B[35][2] +
                mat_A[225][1] * mat_B[43][2] +
                mat_A[225][2] * mat_B[51][2] +
                mat_A[225][3] * mat_B[59][2] +
                mat_A[226][0] * mat_B[67][2] +
                mat_A[226][1] * mat_B[75][2] +
                mat_A[226][2] * mat_B[83][2] +
                mat_A[226][3] * mat_B[91][2] +
                mat_A[227][0] * mat_B[99][2] +
                mat_A[227][1] * mat_B[107][2] +
                mat_A[227][2] * mat_B[115][2] +
                mat_A[227][3] * mat_B[123][2] +
                mat_A[228][0] * mat_B[131][2] +
                mat_A[228][1] * mat_B[139][2] +
                mat_A[228][2] * mat_B[147][2] +
                mat_A[228][3] * mat_B[155][2] +
                mat_A[229][0] * mat_B[163][2] +
                mat_A[229][1] * mat_B[171][2] +
                mat_A[229][2] * mat_B[179][2] +
                mat_A[229][3] * mat_B[187][2] +
                mat_A[230][0] * mat_B[195][2] +
                mat_A[230][1] * mat_B[203][2] +
                mat_A[230][2] * mat_B[211][2] +
                mat_A[230][3] * mat_B[219][2] +
                mat_A[231][0] * mat_B[227][2] +
                mat_A[231][1] * mat_B[235][2] +
                mat_A[231][2] * mat_B[243][2] +
                mat_A[231][3] * mat_B[251][2];
    mat_C[227][3] <=
                mat_A[224][0] * mat_B[3][3] +
                mat_A[224][1] * mat_B[11][3] +
                mat_A[224][2] * mat_B[19][3] +
                mat_A[224][3] * mat_B[27][3] +
                mat_A[225][0] * mat_B[35][3] +
                mat_A[225][1] * mat_B[43][3] +
                mat_A[225][2] * mat_B[51][3] +
                mat_A[225][3] * mat_B[59][3] +
                mat_A[226][0] * mat_B[67][3] +
                mat_A[226][1] * mat_B[75][3] +
                mat_A[226][2] * mat_B[83][3] +
                mat_A[226][3] * mat_B[91][3] +
                mat_A[227][0] * mat_B[99][3] +
                mat_A[227][1] * mat_B[107][3] +
                mat_A[227][2] * mat_B[115][3] +
                mat_A[227][3] * mat_B[123][3] +
                mat_A[228][0] * mat_B[131][3] +
                mat_A[228][1] * mat_B[139][3] +
                mat_A[228][2] * mat_B[147][3] +
                mat_A[228][3] * mat_B[155][3] +
                mat_A[229][0] * mat_B[163][3] +
                mat_A[229][1] * mat_B[171][3] +
                mat_A[229][2] * mat_B[179][3] +
                mat_A[229][3] * mat_B[187][3] +
                mat_A[230][0] * mat_B[195][3] +
                mat_A[230][1] * mat_B[203][3] +
                mat_A[230][2] * mat_B[211][3] +
                mat_A[230][3] * mat_B[219][3] +
                mat_A[231][0] * mat_B[227][3] +
                mat_A[231][1] * mat_B[235][3] +
                mat_A[231][2] * mat_B[243][3] +
                mat_A[231][3] * mat_B[251][3];
    mat_C[228][0] <=
                mat_A[224][0] * mat_B[4][0] +
                mat_A[224][1] * mat_B[12][0] +
                mat_A[224][2] * mat_B[20][0] +
                mat_A[224][3] * mat_B[28][0] +
                mat_A[225][0] * mat_B[36][0] +
                mat_A[225][1] * mat_B[44][0] +
                mat_A[225][2] * mat_B[52][0] +
                mat_A[225][3] * mat_B[60][0] +
                mat_A[226][0] * mat_B[68][0] +
                mat_A[226][1] * mat_B[76][0] +
                mat_A[226][2] * mat_B[84][0] +
                mat_A[226][3] * mat_B[92][0] +
                mat_A[227][0] * mat_B[100][0] +
                mat_A[227][1] * mat_B[108][0] +
                mat_A[227][2] * mat_B[116][0] +
                mat_A[227][3] * mat_B[124][0] +
                mat_A[228][0] * mat_B[132][0] +
                mat_A[228][1] * mat_B[140][0] +
                mat_A[228][2] * mat_B[148][0] +
                mat_A[228][3] * mat_B[156][0] +
                mat_A[229][0] * mat_B[164][0] +
                mat_A[229][1] * mat_B[172][0] +
                mat_A[229][2] * mat_B[180][0] +
                mat_A[229][3] * mat_B[188][0] +
                mat_A[230][0] * mat_B[196][0] +
                mat_A[230][1] * mat_B[204][0] +
                mat_A[230][2] * mat_B[212][0] +
                mat_A[230][3] * mat_B[220][0] +
                mat_A[231][0] * mat_B[228][0] +
                mat_A[231][1] * mat_B[236][0] +
                mat_A[231][2] * mat_B[244][0] +
                mat_A[231][3] * mat_B[252][0];
    mat_C[228][1] <=
                mat_A[224][0] * mat_B[4][1] +
                mat_A[224][1] * mat_B[12][1] +
                mat_A[224][2] * mat_B[20][1] +
                mat_A[224][3] * mat_B[28][1] +
                mat_A[225][0] * mat_B[36][1] +
                mat_A[225][1] * mat_B[44][1] +
                mat_A[225][2] * mat_B[52][1] +
                mat_A[225][3] * mat_B[60][1] +
                mat_A[226][0] * mat_B[68][1] +
                mat_A[226][1] * mat_B[76][1] +
                mat_A[226][2] * mat_B[84][1] +
                mat_A[226][3] * mat_B[92][1] +
                mat_A[227][0] * mat_B[100][1] +
                mat_A[227][1] * mat_B[108][1] +
                mat_A[227][2] * mat_B[116][1] +
                mat_A[227][3] * mat_B[124][1] +
                mat_A[228][0] * mat_B[132][1] +
                mat_A[228][1] * mat_B[140][1] +
                mat_A[228][2] * mat_B[148][1] +
                mat_A[228][3] * mat_B[156][1] +
                mat_A[229][0] * mat_B[164][1] +
                mat_A[229][1] * mat_B[172][1] +
                mat_A[229][2] * mat_B[180][1] +
                mat_A[229][3] * mat_B[188][1] +
                mat_A[230][0] * mat_B[196][1] +
                mat_A[230][1] * mat_B[204][1] +
                mat_A[230][2] * mat_B[212][1] +
                mat_A[230][3] * mat_B[220][1] +
                mat_A[231][0] * mat_B[228][1] +
                mat_A[231][1] * mat_B[236][1] +
                mat_A[231][2] * mat_B[244][1] +
                mat_A[231][3] * mat_B[252][1];
    mat_C[228][2] <=
                mat_A[224][0] * mat_B[4][2] +
                mat_A[224][1] * mat_B[12][2] +
                mat_A[224][2] * mat_B[20][2] +
                mat_A[224][3] * mat_B[28][2] +
                mat_A[225][0] * mat_B[36][2] +
                mat_A[225][1] * mat_B[44][2] +
                mat_A[225][2] * mat_B[52][2] +
                mat_A[225][3] * mat_B[60][2] +
                mat_A[226][0] * mat_B[68][2] +
                mat_A[226][1] * mat_B[76][2] +
                mat_A[226][2] * mat_B[84][2] +
                mat_A[226][3] * mat_B[92][2] +
                mat_A[227][0] * mat_B[100][2] +
                mat_A[227][1] * mat_B[108][2] +
                mat_A[227][2] * mat_B[116][2] +
                mat_A[227][3] * mat_B[124][2] +
                mat_A[228][0] * mat_B[132][2] +
                mat_A[228][1] * mat_B[140][2] +
                mat_A[228][2] * mat_B[148][2] +
                mat_A[228][3] * mat_B[156][2] +
                mat_A[229][0] * mat_B[164][2] +
                mat_A[229][1] * mat_B[172][2] +
                mat_A[229][2] * mat_B[180][2] +
                mat_A[229][3] * mat_B[188][2] +
                mat_A[230][0] * mat_B[196][2] +
                mat_A[230][1] * mat_B[204][2] +
                mat_A[230][2] * mat_B[212][2] +
                mat_A[230][3] * mat_B[220][2] +
                mat_A[231][0] * mat_B[228][2] +
                mat_A[231][1] * mat_B[236][2] +
                mat_A[231][2] * mat_B[244][2] +
                mat_A[231][3] * mat_B[252][2];
    mat_C[228][3] <=
                mat_A[224][0] * mat_B[4][3] +
                mat_A[224][1] * mat_B[12][3] +
                mat_A[224][2] * mat_B[20][3] +
                mat_A[224][3] * mat_B[28][3] +
                mat_A[225][0] * mat_B[36][3] +
                mat_A[225][1] * mat_B[44][3] +
                mat_A[225][2] * mat_B[52][3] +
                mat_A[225][3] * mat_B[60][3] +
                mat_A[226][0] * mat_B[68][3] +
                mat_A[226][1] * mat_B[76][3] +
                mat_A[226][2] * mat_B[84][3] +
                mat_A[226][3] * mat_B[92][3] +
                mat_A[227][0] * mat_B[100][3] +
                mat_A[227][1] * mat_B[108][3] +
                mat_A[227][2] * mat_B[116][3] +
                mat_A[227][3] * mat_B[124][3] +
                mat_A[228][0] * mat_B[132][3] +
                mat_A[228][1] * mat_B[140][3] +
                mat_A[228][2] * mat_B[148][3] +
                mat_A[228][3] * mat_B[156][3] +
                mat_A[229][0] * mat_B[164][3] +
                mat_A[229][1] * mat_B[172][3] +
                mat_A[229][2] * mat_B[180][3] +
                mat_A[229][3] * mat_B[188][3] +
                mat_A[230][0] * mat_B[196][3] +
                mat_A[230][1] * mat_B[204][3] +
                mat_A[230][2] * mat_B[212][3] +
                mat_A[230][3] * mat_B[220][3] +
                mat_A[231][0] * mat_B[228][3] +
                mat_A[231][1] * mat_B[236][3] +
                mat_A[231][2] * mat_B[244][3] +
                mat_A[231][3] * mat_B[252][3];
    mat_C[229][0] <=
                mat_A[224][0] * mat_B[5][0] +
                mat_A[224][1] * mat_B[13][0] +
                mat_A[224][2] * mat_B[21][0] +
                mat_A[224][3] * mat_B[29][0] +
                mat_A[225][0] * mat_B[37][0] +
                mat_A[225][1] * mat_B[45][0] +
                mat_A[225][2] * mat_B[53][0] +
                mat_A[225][3] * mat_B[61][0] +
                mat_A[226][0] * mat_B[69][0] +
                mat_A[226][1] * mat_B[77][0] +
                mat_A[226][2] * mat_B[85][0] +
                mat_A[226][3] * mat_B[93][0] +
                mat_A[227][0] * mat_B[101][0] +
                mat_A[227][1] * mat_B[109][0] +
                mat_A[227][2] * mat_B[117][0] +
                mat_A[227][3] * mat_B[125][0] +
                mat_A[228][0] * mat_B[133][0] +
                mat_A[228][1] * mat_B[141][0] +
                mat_A[228][2] * mat_B[149][0] +
                mat_A[228][3] * mat_B[157][0] +
                mat_A[229][0] * mat_B[165][0] +
                mat_A[229][1] * mat_B[173][0] +
                mat_A[229][2] * mat_B[181][0] +
                mat_A[229][3] * mat_B[189][0] +
                mat_A[230][0] * mat_B[197][0] +
                mat_A[230][1] * mat_B[205][0] +
                mat_A[230][2] * mat_B[213][0] +
                mat_A[230][3] * mat_B[221][0] +
                mat_A[231][0] * mat_B[229][0] +
                mat_A[231][1] * mat_B[237][0] +
                mat_A[231][2] * mat_B[245][0] +
                mat_A[231][3] * mat_B[253][0];
    mat_C[229][1] <=
                mat_A[224][0] * mat_B[5][1] +
                mat_A[224][1] * mat_B[13][1] +
                mat_A[224][2] * mat_B[21][1] +
                mat_A[224][3] * mat_B[29][1] +
                mat_A[225][0] * mat_B[37][1] +
                mat_A[225][1] * mat_B[45][1] +
                mat_A[225][2] * mat_B[53][1] +
                mat_A[225][3] * mat_B[61][1] +
                mat_A[226][0] * mat_B[69][1] +
                mat_A[226][1] * mat_B[77][1] +
                mat_A[226][2] * mat_B[85][1] +
                mat_A[226][3] * mat_B[93][1] +
                mat_A[227][0] * mat_B[101][1] +
                mat_A[227][1] * mat_B[109][1] +
                mat_A[227][2] * mat_B[117][1] +
                mat_A[227][3] * mat_B[125][1] +
                mat_A[228][0] * mat_B[133][1] +
                mat_A[228][1] * mat_B[141][1] +
                mat_A[228][2] * mat_B[149][1] +
                mat_A[228][3] * mat_B[157][1] +
                mat_A[229][0] * mat_B[165][1] +
                mat_A[229][1] * mat_B[173][1] +
                mat_A[229][2] * mat_B[181][1] +
                mat_A[229][3] * mat_B[189][1] +
                mat_A[230][0] * mat_B[197][1] +
                mat_A[230][1] * mat_B[205][1] +
                mat_A[230][2] * mat_B[213][1] +
                mat_A[230][3] * mat_B[221][1] +
                mat_A[231][0] * mat_B[229][1] +
                mat_A[231][1] * mat_B[237][1] +
                mat_A[231][2] * mat_B[245][1] +
                mat_A[231][3] * mat_B[253][1];
    mat_C[229][2] <=
                mat_A[224][0] * mat_B[5][2] +
                mat_A[224][1] * mat_B[13][2] +
                mat_A[224][2] * mat_B[21][2] +
                mat_A[224][3] * mat_B[29][2] +
                mat_A[225][0] * mat_B[37][2] +
                mat_A[225][1] * mat_B[45][2] +
                mat_A[225][2] * mat_B[53][2] +
                mat_A[225][3] * mat_B[61][2] +
                mat_A[226][0] * mat_B[69][2] +
                mat_A[226][1] * mat_B[77][2] +
                mat_A[226][2] * mat_B[85][2] +
                mat_A[226][3] * mat_B[93][2] +
                mat_A[227][0] * mat_B[101][2] +
                mat_A[227][1] * mat_B[109][2] +
                mat_A[227][2] * mat_B[117][2] +
                mat_A[227][3] * mat_B[125][2] +
                mat_A[228][0] * mat_B[133][2] +
                mat_A[228][1] * mat_B[141][2] +
                mat_A[228][2] * mat_B[149][2] +
                mat_A[228][3] * mat_B[157][2] +
                mat_A[229][0] * mat_B[165][2] +
                mat_A[229][1] * mat_B[173][2] +
                mat_A[229][2] * mat_B[181][2] +
                mat_A[229][3] * mat_B[189][2] +
                mat_A[230][0] * mat_B[197][2] +
                mat_A[230][1] * mat_B[205][2] +
                mat_A[230][2] * mat_B[213][2] +
                mat_A[230][3] * mat_B[221][2] +
                mat_A[231][0] * mat_B[229][2] +
                mat_A[231][1] * mat_B[237][2] +
                mat_A[231][2] * mat_B[245][2] +
                mat_A[231][3] * mat_B[253][2];
    mat_C[229][3] <=
                mat_A[224][0] * mat_B[5][3] +
                mat_A[224][1] * mat_B[13][3] +
                mat_A[224][2] * mat_B[21][3] +
                mat_A[224][3] * mat_B[29][3] +
                mat_A[225][0] * mat_B[37][3] +
                mat_A[225][1] * mat_B[45][3] +
                mat_A[225][2] * mat_B[53][3] +
                mat_A[225][3] * mat_B[61][3] +
                mat_A[226][0] * mat_B[69][3] +
                mat_A[226][1] * mat_B[77][3] +
                mat_A[226][2] * mat_B[85][3] +
                mat_A[226][3] * mat_B[93][3] +
                mat_A[227][0] * mat_B[101][3] +
                mat_A[227][1] * mat_B[109][3] +
                mat_A[227][2] * mat_B[117][3] +
                mat_A[227][3] * mat_B[125][3] +
                mat_A[228][0] * mat_B[133][3] +
                mat_A[228][1] * mat_B[141][3] +
                mat_A[228][2] * mat_B[149][3] +
                mat_A[228][3] * mat_B[157][3] +
                mat_A[229][0] * mat_B[165][3] +
                mat_A[229][1] * mat_B[173][3] +
                mat_A[229][2] * mat_B[181][3] +
                mat_A[229][3] * mat_B[189][3] +
                mat_A[230][0] * mat_B[197][3] +
                mat_A[230][1] * mat_B[205][3] +
                mat_A[230][2] * mat_B[213][3] +
                mat_A[230][3] * mat_B[221][3] +
                mat_A[231][0] * mat_B[229][3] +
                mat_A[231][1] * mat_B[237][3] +
                mat_A[231][2] * mat_B[245][3] +
                mat_A[231][3] * mat_B[253][3];
    mat_C[230][0] <=
                mat_A[224][0] * mat_B[6][0] +
                mat_A[224][1] * mat_B[14][0] +
                mat_A[224][2] * mat_B[22][0] +
                mat_A[224][3] * mat_B[30][0] +
                mat_A[225][0] * mat_B[38][0] +
                mat_A[225][1] * mat_B[46][0] +
                mat_A[225][2] * mat_B[54][0] +
                mat_A[225][3] * mat_B[62][0] +
                mat_A[226][0] * mat_B[70][0] +
                mat_A[226][1] * mat_B[78][0] +
                mat_A[226][2] * mat_B[86][0] +
                mat_A[226][3] * mat_B[94][0] +
                mat_A[227][0] * mat_B[102][0] +
                mat_A[227][1] * mat_B[110][0] +
                mat_A[227][2] * mat_B[118][0] +
                mat_A[227][3] * mat_B[126][0] +
                mat_A[228][0] * mat_B[134][0] +
                mat_A[228][1] * mat_B[142][0] +
                mat_A[228][2] * mat_B[150][0] +
                mat_A[228][3] * mat_B[158][0] +
                mat_A[229][0] * mat_B[166][0] +
                mat_A[229][1] * mat_B[174][0] +
                mat_A[229][2] * mat_B[182][0] +
                mat_A[229][3] * mat_B[190][0] +
                mat_A[230][0] * mat_B[198][0] +
                mat_A[230][1] * mat_B[206][0] +
                mat_A[230][2] * mat_B[214][0] +
                mat_A[230][3] * mat_B[222][0] +
                mat_A[231][0] * mat_B[230][0] +
                mat_A[231][1] * mat_B[238][0] +
                mat_A[231][2] * mat_B[246][0] +
                mat_A[231][3] * mat_B[254][0];
    mat_C[230][1] <=
                mat_A[224][0] * mat_B[6][1] +
                mat_A[224][1] * mat_B[14][1] +
                mat_A[224][2] * mat_B[22][1] +
                mat_A[224][3] * mat_B[30][1] +
                mat_A[225][0] * mat_B[38][1] +
                mat_A[225][1] * mat_B[46][1] +
                mat_A[225][2] * mat_B[54][1] +
                mat_A[225][3] * mat_B[62][1] +
                mat_A[226][0] * mat_B[70][1] +
                mat_A[226][1] * mat_B[78][1] +
                mat_A[226][2] * mat_B[86][1] +
                mat_A[226][3] * mat_B[94][1] +
                mat_A[227][0] * mat_B[102][1] +
                mat_A[227][1] * mat_B[110][1] +
                mat_A[227][2] * mat_B[118][1] +
                mat_A[227][3] * mat_B[126][1] +
                mat_A[228][0] * mat_B[134][1] +
                mat_A[228][1] * mat_B[142][1] +
                mat_A[228][2] * mat_B[150][1] +
                mat_A[228][3] * mat_B[158][1] +
                mat_A[229][0] * mat_B[166][1] +
                mat_A[229][1] * mat_B[174][1] +
                mat_A[229][2] * mat_B[182][1] +
                mat_A[229][3] * mat_B[190][1] +
                mat_A[230][0] * mat_B[198][1] +
                mat_A[230][1] * mat_B[206][1] +
                mat_A[230][2] * mat_B[214][1] +
                mat_A[230][3] * mat_B[222][1] +
                mat_A[231][0] * mat_B[230][1] +
                mat_A[231][1] * mat_B[238][1] +
                mat_A[231][2] * mat_B[246][1] +
                mat_A[231][3] * mat_B[254][1];
    mat_C[230][2] <=
                mat_A[224][0] * mat_B[6][2] +
                mat_A[224][1] * mat_B[14][2] +
                mat_A[224][2] * mat_B[22][2] +
                mat_A[224][3] * mat_B[30][2] +
                mat_A[225][0] * mat_B[38][2] +
                mat_A[225][1] * mat_B[46][2] +
                mat_A[225][2] * mat_B[54][2] +
                mat_A[225][3] * mat_B[62][2] +
                mat_A[226][0] * mat_B[70][2] +
                mat_A[226][1] * mat_B[78][2] +
                mat_A[226][2] * mat_B[86][2] +
                mat_A[226][3] * mat_B[94][2] +
                mat_A[227][0] * mat_B[102][2] +
                mat_A[227][1] * mat_B[110][2] +
                mat_A[227][2] * mat_B[118][2] +
                mat_A[227][3] * mat_B[126][2] +
                mat_A[228][0] * mat_B[134][2] +
                mat_A[228][1] * mat_B[142][2] +
                mat_A[228][2] * mat_B[150][2] +
                mat_A[228][3] * mat_B[158][2] +
                mat_A[229][0] * mat_B[166][2] +
                mat_A[229][1] * mat_B[174][2] +
                mat_A[229][2] * mat_B[182][2] +
                mat_A[229][3] * mat_B[190][2] +
                mat_A[230][0] * mat_B[198][2] +
                mat_A[230][1] * mat_B[206][2] +
                mat_A[230][2] * mat_B[214][2] +
                mat_A[230][3] * mat_B[222][2] +
                mat_A[231][0] * mat_B[230][2] +
                mat_A[231][1] * mat_B[238][2] +
                mat_A[231][2] * mat_B[246][2] +
                mat_A[231][3] * mat_B[254][2];
    mat_C[230][3] <=
                mat_A[224][0] * mat_B[6][3] +
                mat_A[224][1] * mat_B[14][3] +
                mat_A[224][2] * mat_B[22][3] +
                mat_A[224][3] * mat_B[30][3] +
                mat_A[225][0] * mat_B[38][3] +
                mat_A[225][1] * mat_B[46][3] +
                mat_A[225][2] * mat_B[54][3] +
                mat_A[225][3] * mat_B[62][3] +
                mat_A[226][0] * mat_B[70][3] +
                mat_A[226][1] * mat_B[78][3] +
                mat_A[226][2] * mat_B[86][3] +
                mat_A[226][3] * mat_B[94][3] +
                mat_A[227][0] * mat_B[102][3] +
                mat_A[227][1] * mat_B[110][3] +
                mat_A[227][2] * mat_B[118][3] +
                mat_A[227][3] * mat_B[126][3] +
                mat_A[228][0] * mat_B[134][3] +
                mat_A[228][1] * mat_B[142][3] +
                mat_A[228][2] * mat_B[150][3] +
                mat_A[228][3] * mat_B[158][3] +
                mat_A[229][0] * mat_B[166][3] +
                mat_A[229][1] * mat_B[174][3] +
                mat_A[229][2] * mat_B[182][3] +
                mat_A[229][3] * mat_B[190][3] +
                mat_A[230][0] * mat_B[198][3] +
                mat_A[230][1] * mat_B[206][3] +
                mat_A[230][2] * mat_B[214][3] +
                mat_A[230][3] * mat_B[222][3] +
                mat_A[231][0] * mat_B[230][3] +
                mat_A[231][1] * mat_B[238][3] +
                mat_A[231][2] * mat_B[246][3] +
                mat_A[231][3] * mat_B[254][3];
    mat_C[231][0] <=
                mat_A[224][0] * mat_B[7][0] +
                mat_A[224][1] * mat_B[15][0] +
                mat_A[224][2] * mat_B[23][0] +
                mat_A[224][3] * mat_B[31][0] +
                mat_A[225][0] * mat_B[39][0] +
                mat_A[225][1] * mat_B[47][0] +
                mat_A[225][2] * mat_B[55][0] +
                mat_A[225][3] * mat_B[63][0] +
                mat_A[226][0] * mat_B[71][0] +
                mat_A[226][1] * mat_B[79][0] +
                mat_A[226][2] * mat_B[87][0] +
                mat_A[226][3] * mat_B[95][0] +
                mat_A[227][0] * mat_B[103][0] +
                mat_A[227][1] * mat_B[111][0] +
                mat_A[227][2] * mat_B[119][0] +
                mat_A[227][3] * mat_B[127][0] +
                mat_A[228][0] * mat_B[135][0] +
                mat_A[228][1] * mat_B[143][0] +
                mat_A[228][2] * mat_B[151][0] +
                mat_A[228][3] * mat_B[159][0] +
                mat_A[229][0] * mat_B[167][0] +
                mat_A[229][1] * mat_B[175][0] +
                mat_A[229][2] * mat_B[183][0] +
                mat_A[229][3] * mat_B[191][0] +
                mat_A[230][0] * mat_B[199][0] +
                mat_A[230][1] * mat_B[207][0] +
                mat_A[230][2] * mat_B[215][0] +
                mat_A[230][3] * mat_B[223][0] +
                mat_A[231][0] * mat_B[231][0] +
                mat_A[231][1] * mat_B[239][0] +
                mat_A[231][2] * mat_B[247][0] +
                mat_A[231][3] * mat_B[255][0];
    mat_C[231][1] <=
                mat_A[224][0] * mat_B[7][1] +
                mat_A[224][1] * mat_B[15][1] +
                mat_A[224][2] * mat_B[23][1] +
                mat_A[224][3] * mat_B[31][1] +
                mat_A[225][0] * mat_B[39][1] +
                mat_A[225][1] * mat_B[47][1] +
                mat_A[225][2] * mat_B[55][1] +
                mat_A[225][3] * mat_B[63][1] +
                mat_A[226][0] * mat_B[71][1] +
                mat_A[226][1] * mat_B[79][1] +
                mat_A[226][2] * mat_B[87][1] +
                mat_A[226][3] * mat_B[95][1] +
                mat_A[227][0] * mat_B[103][1] +
                mat_A[227][1] * mat_B[111][1] +
                mat_A[227][2] * mat_B[119][1] +
                mat_A[227][3] * mat_B[127][1] +
                mat_A[228][0] * mat_B[135][1] +
                mat_A[228][1] * mat_B[143][1] +
                mat_A[228][2] * mat_B[151][1] +
                mat_A[228][3] * mat_B[159][1] +
                mat_A[229][0] * mat_B[167][1] +
                mat_A[229][1] * mat_B[175][1] +
                mat_A[229][2] * mat_B[183][1] +
                mat_A[229][3] * mat_B[191][1] +
                mat_A[230][0] * mat_B[199][1] +
                mat_A[230][1] * mat_B[207][1] +
                mat_A[230][2] * mat_B[215][1] +
                mat_A[230][3] * mat_B[223][1] +
                mat_A[231][0] * mat_B[231][1] +
                mat_A[231][1] * mat_B[239][1] +
                mat_A[231][2] * mat_B[247][1] +
                mat_A[231][3] * mat_B[255][1];
    mat_C[231][2] <=
                mat_A[224][0] * mat_B[7][2] +
                mat_A[224][1] * mat_B[15][2] +
                mat_A[224][2] * mat_B[23][2] +
                mat_A[224][3] * mat_B[31][2] +
                mat_A[225][0] * mat_B[39][2] +
                mat_A[225][1] * mat_B[47][2] +
                mat_A[225][2] * mat_B[55][2] +
                mat_A[225][3] * mat_B[63][2] +
                mat_A[226][0] * mat_B[71][2] +
                mat_A[226][1] * mat_B[79][2] +
                mat_A[226][2] * mat_B[87][2] +
                mat_A[226][3] * mat_B[95][2] +
                mat_A[227][0] * mat_B[103][2] +
                mat_A[227][1] * mat_B[111][2] +
                mat_A[227][2] * mat_B[119][2] +
                mat_A[227][3] * mat_B[127][2] +
                mat_A[228][0] * mat_B[135][2] +
                mat_A[228][1] * mat_B[143][2] +
                mat_A[228][2] * mat_B[151][2] +
                mat_A[228][3] * mat_B[159][2] +
                mat_A[229][0] * mat_B[167][2] +
                mat_A[229][1] * mat_B[175][2] +
                mat_A[229][2] * mat_B[183][2] +
                mat_A[229][3] * mat_B[191][2] +
                mat_A[230][0] * mat_B[199][2] +
                mat_A[230][1] * mat_B[207][2] +
                mat_A[230][2] * mat_B[215][2] +
                mat_A[230][3] * mat_B[223][2] +
                mat_A[231][0] * mat_B[231][2] +
                mat_A[231][1] * mat_B[239][2] +
                mat_A[231][2] * mat_B[247][2] +
                mat_A[231][3] * mat_B[255][2];
    mat_C[231][3] <=
                mat_A[224][0] * mat_B[7][3] +
                mat_A[224][1] * mat_B[15][3] +
                mat_A[224][2] * mat_B[23][3] +
                mat_A[224][3] * mat_B[31][3] +
                mat_A[225][0] * mat_B[39][3] +
                mat_A[225][1] * mat_B[47][3] +
                mat_A[225][2] * mat_B[55][3] +
                mat_A[225][3] * mat_B[63][3] +
                mat_A[226][0] * mat_B[71][3] +
                mat_A[226][1] * mat_B[79][3] +
                mat_A[226][2] * mat_B[87][3] +
                mat_A[226][3] * mat_B[95][3] +
                mat_A[227][0] * mat_B[103][3] +
                mat_A[227][1] * mat_B[111][3] +
                mat_A[227][2] * mat_B[119][3] +
                mat_A[227][3] * mat_B[127][3] +
                mat_A[228][0] * mat_B[135][3] +
                mat_A[228][1] * mat_B[143][3] +
                mat_A[228][2] * mat_B[151][3] +
                mat_A[228][3] * mat_B[159][3] +
                mat_A[229][0] * mat_B[167][3] +
                mat_A[229][1] * mat_B[175][3] +
                mat_A[229][2] * mat_B[183][3] +
                mat_A[229][3] * mat_B[191][3] +
                mat_A[230][0] * mat_B[199][3] +
                mat_A[230][1] * mat_B[207][3] +
                mat_A[230][2] * mat_B[215][3] +
                mat_A[230][3] * mat_B[223][3] +
                mat_A[231][0] * mat_B[231][3] +
                mat_A[231][1] * mat_B[239][3] +
                mat_A[231][2] * mat_B[247][3] +
                mat_A[231][3] * mat_B[255][3];
    mat_C[232][0] <=
                mat_A[232][0] * mat_B[0][0] +
                mat_A[232][1] * mat_B[8][0] +
                mat_A[232][2] * mat_B[16][0] +
                mat_A[232][3] * mat_B[24][0] +
                mat_A[233][0] * mat_B[32][0] +
                mat_A[233][1] * mat_B[40][0] +
                mat_A[233][2] * mat_B[48][0] +
                mat_A[233][3] * mat_B[56][0] +
                mat_A[234][0] * mat_B[64][0] +
                mat_A[234][1] * mat_B[72][0] +
                mat_A[234][2] * mat_B[80][0] +
                mat_A[234][3] * mat_B[88][0] +
                mat_A[235][0] * mat_B[96][0] +
                mat_A[235][1] * mat_B[104][0] +
                mat_A[235][2] * mat_B[112][0] +
                mat_A[235][3] * mat_B[120][0] +
                mat_A[236][0] * mat_B[128][0] +
                mat_A[236][1] * mat_B[136][0] +
                mat_A[236][2] * mat_B[144][0] +
                mat_A[236][3] * mat_B[152][0] +
                mat_A[237][0] * mat_B[160][0] +
                mat_A[237][1] * mat_B[168][0] +
                mat_A[237][2] * mat_B[176][0] +
                mat_A[237][3] * mat_B[184][0] +
                mat_A[238][0] * mat_B[192][0] +
                mat_A[238][1] * mat_B[200][0] +
                mat_A[238][2] * mat_B[208][0] +
                mat_A[238][3] * mat_B[216][0] +
                mat_A[239][0] * mat_B[224][0] +
                mat_A[239][1] * mat_B[232][0] +
                mat_A[239][2] * mat_B[240][0] +
                mat_A[239][3] * mat_B[248][0];
    mat_C[232][1] <=
                mat_A[232][0] * mat_B[0][1] +
                mat_A[232][1] * mat_B[8][1] +
                mat_A[232][2] * mat_B[16][1] +
                mat_A[232][3] * mat_B[24][1] +
                mat_A[233][0] * mat_B[32][1] +
                mat_A[233][1] * mat_B[40][1] +
                mat_A[233][2] * mat_B[48][1] +
                mat_A[233][3] * mat_B[56][1] +
                mat_A[234][0] * mat_B[64][1] +
                mat_A[234][1] * mat_B[72][1] +
                mat_A[234][2] * mat_B[80][1] +
                mat_A[234][3] * mat_B[88][1] +
                mat_A[235][0] * mat_B[96][1] +
                mat_A[235][1] * mat_B[104][1] +
                mat_A[235][2] * mat_B[112][1] +
                mat_A[235][3] * mat_B[120][1] +
                mat_A[236][0] * mat_B[128][1] +
                mat_A[236][1] * mat_B[136][1] +
                mat_A[236][2] * mat_B[144][1] +
                mat_A[236][3] * mat_B[152][1] +
                mat_A[237][0] * mat_B[160][1] +
                mat_A[237][1] * mat_B[168][1] +
                mat_A[237][2] * mat_B[176][1] +
                mat_A[237][3] * mat_B[184][1] +
                mat_A[238][0] * mat_B[192][1] +
                mat_A[238][1] * mat_B[200][1] +
                mat_A[238][2] * mat_B[208][1] +
                mat_A[238][3] * mat_B[216][1] +
                mat_A[239][0] * mat_B[224][1] +
                mat_A[239][1] * mat_B[232][1] +
                mat_A[239][2] * mat_B[240][1] +
                mat_A[239][3] * mat_B[248][1];
    mat_C[232][2] <=
                mat_A[232][0] * mat_B[0][2] +
                mat_A[232][1] * mat_B[8][2] +
                mat_A[232][2] * mat_B[16][2] +
                mat_A[232][3] * mat_B[24][2] +
                mat_A[233][0] * mat_B[32][2] +
                mat_A[233][1] * mat_B[40][2] +
                mat_A[233][2] * mat_B[48][2] +
                mat_A[233][3] * mat_B[56][2] +
                mat_A[234][0] * mat_B[64][2] +
                mat_A[234][1] * mat_B[72][2] +
                mat_A[234][2] * mat_B[80][2] +
                mat_A[234][3] * mat_B[88][2] +
                mat_A[235][0] * mat_B[96][2] +
                mat_A[235][1] * mat_B[104][2] +
                mat_A[235][2] * mat_B[112][2] +
                mat_A[235][3] * mat_B[120][2] +
                mat_A[236][0] * mat_B[128][2] +
                mat_A[236][1] * mat_B[136][2] +
                mat_A[236][2] * mat_B[144][2] +
                mat_A[236][3] * mat_B[152][2] +
                mat_A[237][0] * mat_B[160][2] +
                mat_A[237][1] * mat_B[168][2] +
                mat_A[237][2] * mat_B[176][2] +
                mat_A[237][3] * mat_B[184][2] +
                mat_A[238][0] * mat_B[192][2] +
                mat_A[238][1] * mat_B[200][2] +
                mat_A[238][2] * mat_B[208][2] +
                mat_A[238][3] * mat_B[216][2] +
                mat_A[239][0] * mat_B[224][2] +
                mat_A[239][1] * mat_B[232][2] +
                mat_A[239][2] * mat_B[240][2] +
                mat_A[239][3] * mat_B[248][2];
    mat_C[232][3] <=
                mat_A[232][0] * mat_B[0][3] +
                mat_A[232][1] * mat_B[8][3] +
                mat_A[232][2] * mat_B[16][3] +
                mat_A[232][3] * mat_B[24][3] +
                mat_A[233][0] * mat_B[32][3] +
                mat_A[233][1] * mat_B[40][3] +
                mat_A[233][2] * mat_B[48][3] +
                mat_A[233][3] * mat_B[56][3] +
                mat_A[234][0] * mat_B[64][3] +
                mat_A[234][1] * mat_B[72][3] +
                mat_A[234][2] * mat_B[80][3] +
                mat_A[234][3] * mat_B[88][3] +
                mat_A[235][0] * mat_B[96][3] +
                mat_A[235][1] * mat_B[104][3] +
                mat_A[235][2] * mat_B[112][3] +
                mat_A[235][3] * mat_B[120][3] +
                mat_A[236][0] * mat_B[128][3] +
                mat_A[236][1] * mat_B[136][3] +
                mat_A[236][2] * mat_B[144][3] +
                mat_A[236][3] * mat_B[152][3] +
                mat_A[237][0] * mat_B[160][3] +
                mat_A[237][1] * mat_B[168][3] +
                mat_A[237][2] * mat_B[176][3] +
                mat_A[237][3] * mat_B[184][3] +
                mat_A[238][0] * mat_B[192][3] +
                mat_A[238][1] * mat_B[200][3] +
                mat_A[238][2] * mat_B[208][3] +
                mat_A[238][3] * mat_B[216][3] +
                mat_A[239][0] * mat_B[224][3] +
                mat_A[239][1] * mat_B[232][3] +
                mat_A[239][2] * mat_B[240][3] +
                mat_A[239][3] * mat_B[248][3];
    mat_C[233][0] <=
                mat_A[232][0] * mat_B[1][0] +
                mat_A[232][1] * mat_B[9][0] +
                mat_A[232][2] * mat_B[17][0] +
                mat_A[232][3] * mat_B[25][0] +
                mat_A[233][0] * mat_B[33][0] +
                mat_A[233][1] * mat_B[41][0] +
                mat_A[233][2] * mat_B[49][0] +
                mat_A[233][3] * mat_B[57][0] +
                mat_A[234][0] * mat_B[65][0] +
                mat_A[234][1] * mat_B[73][0] +
                mat_A[234][2] * mat_B[81][0] +
                mat_A[234][3] * mat_B[89][0] +
                mat_A[235][0] * mat_B[97][0] +
                mat_A[235][1] * mat_B[105][0] +
                mat_A[235][2] * mat_B[113][0] +
                mat_A[235][3] * mat_B[121][0] +
                mat_A[236][0] * mat_B[129][0] +
                mat_A[236][1] * mat_B[137][0] +
                mat_A[236][2] * mat_B[145][0] +
                mat_A[236][3] * mat_B[153][0] +
                mat_A[237][0] * mat_B[161][0] +
                mat_A[237][1] * mat_B[169][0] +
                mat_A[237][2] * mat_B[177][0] +
                mat_A[237][3] * mat_B[185][0] +
                mat_A[238][0] * mat_B[193][0] +
                mat_A[238][1] * mat_B[201][0] +
                mat_A[238][2] * mat_B[209][0] +
                mat_A[238][3] * mat_B[217][0] +
                mat_A[239][0] * mat_B[225][0] +
                mat_A[239][1] * mat_B[233][0] +
                mat_A[239][2] * mat_B[241][0] +
                mat_A[239][3] * mat_B[249][0];
    mat_C[233][1] <=
                mat_A[232][0] * mat_B[1][1] +
                mat_A[232][1] * mat_B[9][1] +
                mat_A[232][2] * mat_B[17][1] +
                mat_A[232][3] * mat_B[25][1] +
                mat_A[233][0] * mat_B[33][1] +
                mat_A[233][1] * mat_B[41][1] +
                mat_A[233][2] * mat_B[49][1] +
                mat_A[233][3] * mat_B[57][1] +
                mat_A[234][0] * mat_B[65][1] +
                mat_A[234][1] * mat_B[73][1] +
                mat_A[234][2] * mat_B[81][1] +
                mat_A[234][3] * mat_B[89][1] +
                mat_A[235][0] * mat_B[97][1] +
                mat_A[235][1] * mat_B[105][1] +
                mat_A[235][2] * mat_B[113][1] +
                mat_A[235][3] * mat_B[121][1] +
                mat_A[236][0] * mat_B[129][1] +
                mat_A[236][1] * mat_B[137][1] +
                mat_A[236][2] * mat_B[145][1] +
                mat_A[236][3] * mat_B[153][1] +
                mat_A[237][0] * mat_B[161][1] +
                mat_A[237][1] * mat_B[169][1] +
                mat_A[237][2] * mat_B[177][1] +
                mat_A[237][3] * mat_B[185][1] +
                mat_A[238][0] * mat_B[193][1] +
                mat_A[238][1] * mat_B[201][1] +
                mat_A[238][2] * mat_B[209][1] +
                mat_A[238][3] * mat_B[217][1] +
                mat_A[239][0] * mat_B[225][1] +
                mat_A[239][1] * mat_B[233][1] +
                mat_A[239][2] * mat_B[241][1] +
                mat_A[239][3] * mat_B[249][1];
    mat_C[233][2] <=
                mat_A[232][0] * mat_B[1][2] +
                mat_A[232][1] * mat_B[9][2] +
                mat_A[232][2] * mat_B[17][2] +
                mat_A[232][3] * mat_B[25][2] +
                mat_A[233][0] * mat_B[33][2] +
                mat_A[233][1] * mat_B[41][2] +
                mat_A[233][2] * mat_B[49][2] +
                mat_A[233][3] * mat_B[57][2] +
                mat_A[234][0] * mat_B[65][2] +
                mat_A[234][1] * mat_B[73][2] +
                mat_A[234][2] * mat_B[81][2] +
                mat_A[234][3] * mat_B[89][2] +
                mat_A[235][0] * mat_B[97][2] +
                mat_A[235][1] * mat_B[105][2] +
                mat_A[235][2] * mat_B[113][2] +
                mat_A[235][3] * mat_B[121][2] +
                mat_A[236][0] * mat_B[129][2] +
                mat_A[236][1] * mat_B[137][2] +
                mat_A[236][2] * mat_B[145][2] +
                mat_A[236][3] * mat_B[153][2] +
                mat_A[237][0] * mat_B[161][2] +
                mat_A[237][1] * mat_B[169][2] +
                mat_A[237][2] * mat_B[177][2] +
                mat_A[237][3] * mat_B[185][2] +
                mat_A[238][0] * mat_B[193][2] +
                mat_A[238][1] * mat_B[201][2] +
                mat_A[238][2] * mat_B[209][2] +
                mat_A[238][3] * mat_B[217][2] +
                mat_A[239][0] * mat_B[225][2] +
                mat_A[239][1] * mat_B[233][2] +
                mat_A[239][2] * mat_B[241][2] +
                mat_A[239][3] * mat_B[249][2];
    mat_C[233][3] <=
                mat_A[232][0] * mat_B[1][3] +
                mat_A[232][1] * mat_B[9][3] +
                mat_A[232][2] * mat_B[17][3] +
                mat_A[232][3] * mat_B[25][3] +
                mat_A[233][0] * mat_B[33][3] +
                mat_A[233][1] * mat_B[41][3] +
                mat_A[233][2] * mat_B[49][3] +
                mat_A[233][3] * mat_B[57][3] +
                mat_A[234][0] * mat_B[65][3] +
                mat_A[234][1] * mat_B[73][3] +
                mat_A[234][2] * mat_B[81][3] +
                mat_A[234][3] * mat_B[89][3] +
                mat_A[235][0] * mat_B[97][3] +
                mat_A[235][1] * mat_B[105][3] +
                mat_A[235][2] * mat_B[113][3] +
                mat_A[235][3] * mat_B[121][3] +
                mat_A[236][0] * mat_B[129][3] +
                mat_A[236][1] * mat_B[137][3] +
                mat_A[236][2] * mat_B[145][3] +
                mat_A[236][3] * mat_B[153][3] +
                mat_A[237][0] * mat_B[161][3] +
                mat_A[237][1] * mat_B[169][3] +
                mat_A[237][2] * mat_B[177][3] +
                mat_A[237][3] * mat_B[185][3] +
                mat_A[238][0] * mat_B[193][3] +
                mat_A[238][1] * mat_B[201][3] +
                mat_A[238][2] * mat_B[209][3] +
                mat_A[238][3] * mat_B[217][3] +
                mat_A[239][0] * mat_B[225][3] +
                mat_A[239][1] * mat_B[233][3] +
                mat_A[239][2] * mat_B[241][3] +
                mat_A[239][3] * mat_B[249][3];
    mat_C[234][0] <=
                mat_A[232][0] * mat_B[2][0] +
                mat_A[232][1] * mat_B[10][0] +
                mat_A[232][2] * mat_B[18][0] +
                mat_A[232][3] * mat_B[26][0] +
                mat_A[233][0] * mat_B[34][0] +
                mat_A[233][1] * mat_B[42][0] +
                mat_A[233][2] * mat_B[50][0] +
                mat_A[233][3] * mat_B[58][0] +
                mat_A[234][0] * mat_B[66][0] +
                mat_A[234][1] * mat_B[74][0] +
                mat_A[234][2] * mat_B[82][0] +
                mat_A[234][3] * mat_B[90][0] +
                mat_A[235][0] * mat_B[98][0] +
                mat_A[235][1] * mat_B[106][0] +
                mat_A[235][2] * mat_B[114][0] +
                mat_A[235][3] * mat_B[122][0] +
                mat_A[236][0] * mat_B[130][0] +
                mat_A[236][1] * mat_B[138][0] +
                mat_A[236][2] * mat_B[146][0] +
                mat_A[236][3] * mat_B[154][0] +
                mat_A[237][0] * mat_B[162][0] +
                mat_A[237][1] * mat_B[170][0] +
                mat_A[237][2] * mat_B[178][0] +
                mat_A[237][3] * mat_B[186][0] +
                mat_A[238][0] * mat_B[194][0] +
                mat_A[238][1] * mat_B[202][0] +
                mat_A[238][2] * mat_B[210][0] +
                mat_A[238][3] * mat_B[218][0] +
                mat_A[239][0] * mat_B[226][0] +
                mat_A[239][1] * mat_B[234][0] +
                mat_A[239][2] * mat_B[242][0] +
                mat_A[239][3] * mat_B[250][0];
    mat_C[234][1] <=
                mat_A[232][0] * mat_B[2][1] +
                mat_A[232][1] * mat_B[10][1] +
                mat_A[232][2] * mat_B[18][1] +
                mat_A[232][3] * mat_B[26][1] +
                mat_A[233][0] * mat_B[34][1] +
                mat_A[233][1] * mat_B[42][1] +
                mat_A[233][2] * mat_B[50][1] +
                mat_A[233][3] * mat_B[58][1] +
                mat_A[234][0] * mat_B[66][1] +
                mat_A[234][1] * mat_B[74][1] +
                mat_A[234][2] * mat_B[82][1] +
                mat_A[234][3] * mat_B[90][1] +
                mat_A[235][0] * mat_B[98][1] +
                mat_A[235][1] * mat_B[106][1] +
                mat_A[235][2] * mat_B[114][1] +
                mat_A[235][3] * mat_B[122][1] +
                mat_A[236][0] * mat_B[130][1] +
                mat_A[236][1] * mat_B[138][1] +
                mat_A[236][2] * mat_B[146][1] +
                mat_A[236][3] * mat_B[154][1] +
                mat_A[237][0] * mat_B[162][1] +
                mat_A[237][1] * mat_B[170][1] +
                mat_A[237][2] * mat_B[178][1] +
                mat_A[237][3] * mat_B[186][1] +
                mat_A[238][0] * mat_B[194][1] +
                mat_A[238][1] * mat_B[202][1] +
                mat_A[238][2] * mat_B[210][1] +
                mat_A[238][3] * mat_B[218][1] +
                mat_A[239][0] * mat_B[226][1] +
                mat_A[239][1] * mat_B[234][1] +
                mat_A[239][2] * mat_B[242][1] +
                mat_A[239][3] * mat_B[250][1];
    mat_C[234][2] <=
                mat_A[232][0] * mat_B[2][2] +
                mat_A[232][1] * mat_B[10][2] +
                mat_A[232][2] * mat_B[18][2] +
                mat_A[232][3] * mat_B[26][2] +
                mat_A[233][0] * mat_B[34][2] +
                mat_A[233][1] * mat_B[42][2] +
                mat_A[233][2] * mat_B[50][2] +
                mat_A[233][3] * mat_B[58][2] +
                mat_A[234][0] * mat_B[66][2] +
                mat_A[234][1] * mat_B[74][2] +
                mat_A[234][2] * mat_B[82][2] +
                mat_A[234][3] * mat_B[90][2] +
                mat_A[235][0] * mat_B[98][2] +
                mat_A[235][1] * mat_B[106][2] +
                mat_A[235][2] * mat_B[114][2] +
                mat_A[235][3] * mat_B[122][2] +
                mat_A[236][0] * mat_B[130][2] +
                mat_A[236][1] * mat_B[138][2] +
                mat_A[236][2] * mat_B[146][2] +
                mat_A[236][3] * mat_B[154][2] +
                mat_A[237][0] * mat_B[162][2] +
                mat_A[237][1] * mat_B[170][2] +
                mat_A[237][2] * mat_B[178][2] +
                mat_A[237][3] * mat_B[186][2] +
                mat_A[238][0] * mat_B[194][2] +
                mat_A[238][1] * mat_B[202][2] +
                mat_A[238][2] * mat_B[210][2] +
                mat_A[238][3] * mat_B[218][2] +
                mat_A[239][0] * mat_B[226][2] +
                mat_A[239][1] * mat_B[234][2] +
                mat_A[239][2] * mat_B[242][2] +
                mat_A[239][3] * mat_B[250][2];
    mat_C[234][3] <=
                mat_A[232][0] * mat_B[2][3] +
                mat_A[232][1] * mat_B[10][3] +
                mat_A[232][2] * mat_B[18][3] +
                mat_A[232][3] * mat_B[26][3] +
                mat_A[233][0] * mat_B[34][3] +
                mat_A[233][1] * mat_B[42][3] +
                mat_A[233][2] * mat_B[50][3] +
                mat_A[233][3] * mat_B[58][3] +
                mat_A[234][0] * mat_B[66][3] +
                mat_A[234][1] * mat_B[74][3] +
                mat_A[234][2] * mat_B[82][3] +
                mat_A[234][3] * mat_B[90][3] +
                mat_A[235][0] * mat_B[98][3] +
                mat_A[235][1] * mat_B[106][3] +
                mat_A[235][2] * mat_B[114][3] +
                mat_A[235][3] * mat_B[122][3] +
                mat_A[236][0] * mat_B[130][3] +
                mat_A[236][1] * mat_B[138][3] +
                mat_A[236][2] * mat_B[146][3] +
                mat_A[236][3] * mat_B[154][3] +
                mat_A[237][0] * mat_B[162][3] +
                mat_A[237][1] * mat_B[170][3] +
                mat_A[237][2] * mat_B[178][3] +
                mat_A[237][3] * mat_B[186][3] +
                mat_A[238][0] * mat_B[194][3] +
                mat_A[238][1] * mat_B[202][3] +
                mat_A[238][2] * mat_B[210][3] +
                mat_A[238][3] * mat_B[218][3] +
                mat_A[239][0] * mat_B[226][3] +
                mat_A[239][1] * mat_B[234][3] +
                mat_A[239][2] * mat_B[242][3] +
                mat_A[239][3] * mat_B[250][3];
    mat_C[235][0] <=
                mat_A[232][0] * mat_B[3][0] +
                mat_A[232][1] * mat_B[11][0] +
                mat_A[232][2] * mat_B[19][0] +
                mat_A[232][3] * mat_B[27][0] +
                mat_A[233][0] * mat_B[35][0] +
                mat_A[233][1] * mat_B[43][0] +
                mat_A[233][2] * mat_B[51][0] +
                mat_A[233][3] * mat_B[59][0] +
                mat_A[234][0] * mat_B[67][0] +
                mat_A[234][1] * mat_B[75][0] +
                mat_A[234][2] * mat_B[83][0] +
                mat_A[234][3] * mat_B[91][0] +
                mat_A[235][0] * mat_B[99][0] +
                mat_A[235][1] * mat_B[107][0] +
                mat_A[235][2] * mat_B[115][0] +
                mat_A[235][3] * mat_B[123][0] +
                mat_A[236][0] * mat_B[131][0] +
                mat_A[236][1] * mat_B[139][0] +
                mat_A[236][2] * mat_B[147][0] +
                mat_A[236][3] * mat_B[155][0] +
                mat_A[237][0] * mat_B[163][0] +
                mat_A[237][1] * mat_B[171][0] +
                mat_A[237][2] * mat_B[179][0] +
                mat_A[237][3] * mat_B[187][0] +
                mat_A[238][0] * mat_B[195][0] +
                mat_A[238][1] * mat_B[203][0] +
                mat_A[238][2] * mat_B[211][0] +
                mat_A[238][3] * mat_B[219][0] +
                mat_A[239][0] * mat_B[227][0] +
                mat_A[239][1] * mat_B[235][0] +
                mat_A[239][2] * mat_B[243][0] +
                mat_A[239][3] * mat_B[251][0];
    mat_C[235][1] <=
                mat_A[232][0] * mat_B[3][1] +
                mat_A[232][1] * mat_B[11][1] +
                mat_A[232][2] * mat_B[19][1] +
                mat_A[232][3] * mat_B[27][1] +
                mat_A[233][0] * mat_B[35][1] +
                mat_A[233][1] * mat_B[43][1] +
                mat_A[233][2] * mat_B[51][1] +
                mat_A[233][3] * mat_B[59][1] +
                mat_A[234][0] * mat_B[67][1] +
                mat_A[234][1] * mat_B[75][1] +
                mat_A[234][2] * mat_B[83][1] +
                mat_A[234][3] * mat_B[91][1] +
                mat_A[235][0] * mat_B[99][1] +
                mat_A[235][1] * mat_B[107][1] +
                mat_A[235][2] * mat_B[115][1] +
                mat_A[235][3] * mat_B[123][1] +
                mat_A[236][0] * mat_B[131][1] +
                mat_A[236][1] * mat_B[139][1] +
                mat_A[236][2] * mat_B[147][1] +
                mat_A[236][3] * mat_B[155][1] +
                mat_A[237][0] * mat_B[163][1] +
                mat_A[237][1] * mat_B[171][1] +
                mat_A[237][2] * mat_B[179][1] +
                mat_A[237][3] * mat_B[187][1] +
                mat_A[238][0] * mat_B[195][1] +
                mat_A[238][1] * mat_B[203][1] +
                mat_A[238][2] * mat_B[211][1] +
                mat_A[238][3] * mat_B[219][1] +
                mat_A[239][0] * mat_B[227][1] +
                mat_A[239][1] * mat_B[235][1] +
                mat_A[239][2] * mat_B[243][1] +
                mat_A[239][3] * mat_B[251][1];
    mat_C[235][2] <=
                mat_A[232][0] * mat_B[3][2] +
                mat_A[232][1] * mat_B[11][2] +
                mat_A[232][2] * mat_B[19][2] +
                mat_A[232][3] * mat_B[27][2] +
                mat_A[233][0] * mat_B[35][2] +
                mat_A[233][1] * mat_B[43][2] +
                mat_A[233][2] * mat_B[51][2] +
                mat_A[233][3] * mat_B[59][2] +
                mat_A[234][0] * mat_B[67][2] +
                mat_A[234][1] * mat_B[75][2] +
                mat_A[234][2] * mat_B[83][2] +
                mat_A[234][3] * mat_B[91][2] +
                mat_A[235][0] * mat_B[99][2] +
                mat_A[235][1] * mat_B[107][2] +
                mat_A[235][2] * mat_B[115][2] +
                mat_A[235][3] * mat_B[123][2] +
                mat_A[236][0] * mat_B[131][2] +
                mat_A[236][1] * mat_B[139][2] +
                mat_A[236][2] * mat_B[147][2] +
                mat_A[236][3] * mat_B[155][2] +
                mat_A[237][0] * mat_B[163][2] +
                mat_A[237][1] * mat_B[171][2] +
                mat_A[237][2] * mat_B[179][2] +
                mat_A[237][3] * mat_B[187][2] +
                mat_A[238][0] * mat_B[195][2] +
                mat_A[238][1] * mat_B[203][2] +
                mat_A[238][2] * mat_B[211][2] +
                mat_A[238][3] * mat_B[219][2] +
                mat_A[239][0] * mat_B[227][2] +
                mat_A[239][1] * mat_B[235][2] +
                mat_A[239][2] * mat_B[243][2] +
                mat_A[239][3] * mat_B[251][2];
    mat_C[235][3] <=
                mat_A[232][0] * mat_B[3][3] +
                mat_A[232][1] * mat_B[11][3] +
                mat_A[232][2] * mat_B[19][3] +
                mat_A[232][3] * mat_B[27][3] +
                mat_A[233][0] * mat_B[35][3] +
                mat_A[233][1] * mat_B[43][3] +
                mat_A[233][2] * mat_B[51][3] +
                mat_A[233][3] * mat_B[59][3] +
                mat_A[234][0] * mat_B[67][3] +
                mat_A[234][1] * mat_B[75][3] +
                mat_A[234][2] * mat_B[83][3] +
                mat_A[234][3] * mat_B[91][3] +
                mat_A[235][0] * mat_B[99][3] +
                mat_A[235][1] * mat_B[107][3] +
                mat_A[235][2] * mat_B[115][3] +
                mat_A[235][3] * mat_B[123][3] +
                mat_A[236][0] * mat_B[131][3] +
                mat_A[236][1] * mat_B[139][3] +
                mat_A[236][2] * mat_B[147][3] +
                mat_A[236][3] * mat_B[155][3] +
                mat_A[237][0] * mat_B[163][3] +
                mat_A[237][1] * mat_B[171][3] +
                mat_A[237][2] * mat_B[179][3] +
                mat_A[237][3] * mat_B[187][3] +
                mat_A[238][0] * mat_B[195][3] +
                mat_A[238][1] * mat_B[203][3] +
                mat_A[238][2] * mat_B[211][3] +
                mat_A[238][3] * mat_B[219][3] +
                mat_A[239][0] * mat_B[227][3] +
                mat_A[239][1] * mat_B[235][3] +
                mat_A[239][2] * mat_B[243][3] +
                mat_A[239][3] * mat_B[251][3];
    mat_C[236][0] <=
                mat_A[232][0] * mat_B[4][0] +
                mat_A[232][1] * mat_B[12][0] +
                mat_A[232][2] * mat_B[20][0] +
                mat_A[232][3] * mat_B[28][0] +
                mat_A[233][0] * mat_B[36][0] +
                mat_A[233][1] * mat_B[44][0] +
                mat_A[233][2] * mat_B[52][0] +
                mat_A[233][3] * mat_B[60][0] +
                mat_A[234][0] * mat_B[68][0] +
                mat_A[234][1] * mat_B[76][0] +
                mat_A[234][2] * mat_B[84][0] +
                mat_A[234][3] * mat_B[92][0] +
                mat_A[235][0] * mat_B[100][0] +
                mat_A[235][1] * mat_B[108][0] +
                mat_A[235][2] * mat_B[116][0] +
                mat_A[235][3] * mat_B[124][0] +
                mat_A[236][0] * mat_B[132][0] +
                mat_A[236][1] * mat_B[140][0] +
                mat_A[236][2] * mat_B[148][0] +
                mat_A[236][3] * mat_B[156][0] +
                mat_A[237][0] * mat_B[164][0] +
                mat_A[237][1] * mat_B[172][0] +
                mat_A[237][2] * mat_B[180][0] +
                mat_A[237][3] * mat_B[188][0] +
                mat_A[238][0] * mat_B[196][0] +
                mat_A[238][1] * mat_B[204][0] +
                mat_A[238][2] * mat_B[212][0] +
                mat_A[238][3] * mat_B[220][0] +
                mat_A[239][0] * mat_B[228][0] +
                mat_A[239][1] * mat_B[236][0] +
                mat_A[239][2] * mat_B[244][0] +
                mat_A[239][3] * mat_B[252][0];
    mat_C[236][1] <=
                mat_A[232][0] * mat_B[4][1] +
                mat_A[232][1] * mat_B[12][1] +
                mat_A[232][2] * mat_B[20][1] +
                mat_A[232][3] * mat_B[28][1] +
                mat_A[233][0] * mat_B[36][1] +
                mat_A[233][1] * mat_B[44][1] +
                mat_A[233][2] * mat_B[52][1] +
                mat_A[233][3] * mat_B[60][1] +
                mat_A[234][0] * mat_B[68][1] +
                mat_A[234][1] * mat_B[76][1] +
                mat_A[234][2] * mat_B[84][1] +
                mat_A[234][3] * mat_B[92][1] +
                mat_A[235][0] * mat_B[100][1] +
                mat_A[235][1] * mat_B[108][1] +
                mat_A[235][2] * mat_B[116][1] +
                mat_A[235][3] * mat_B[124][1] +
                mat_A[236][0] * mat_B[132][1] +
                mat_A[236][1] * mat_B[140][1] +
                mat_A[236][2] * mat_B[148][1] +
                mat_A[236][3] * mat_B[156][1] +
                mat_A[237][0] * mat_B[164][1] +
                mat_A[237][1] * mat_B[172][1] +
                mat_A[237][2] * mat_B[180][1] +
                mat_A[237][3] * mat_B[188][1] +
                mat_A[238][0] * mat_B[196][1] +
                mat_A[238][1] * mat_B[204][1] +
                mat_A[238][2] * mat_B[212][1] +
                mat_A[238][3] * mat_B[220][1] +
                mat_A[239][0] * mat_B[228][1] +
                mat_A[239][1] * mat_B[236][1] +
                mat_A[239][2] * mat_B[244][1] +
                mat_A[239][3] * mat_B[252][1];
    mat_C[236][2] <=
                mat_A[232][0] * mat_B[4][2] +
                mat_A[232][1] * mat_B[12][2] +
                mat_A[232][2] * mat_B[20][2] +
                mat_A[232][3] * mat_B[28][2] +
                mat_A[233][0] * mat_B[36][2] +
                mat_A[233][1] * mat_B[44][2] +
                mat_A[233][2] * mat_B[52][2] +
                mat_A[233][3] * mat_B[60][2] +
                mat_A[234][0] * mat_B[68][2] +
                mat_A[234][1] * mat_B[76][2] +
                mat_A[234][2] * mat_B[84][2] +
                mat_A[234][3] * mat_B[92][2] +
                mat_A[235][0] * mat_B[100][2] +
                mat_A[235][1] * mat_B[108][2] +
                mat_A[235][2] * mat_B[116][2] +
                mat_A[235][3] * mat_B[124][2] +
                mat_A[236][0] * mat_B[132][2] +
                mat_A[236][1] * mat_B[140][2] +
                mat_A[236][2] * mat_B[148][2] +
                mat_A[236][3] * mat_B[156][2] +
                mat_A[237][0] * mat_B[164][2] +
                mat_A[237][1] * mat_B[172][2] +
                mat_A[237][2] * mat_B[180][2] +
                mat_A[237][3] * mat_B[188][2] +
                mat_A[238][0] * mat_B[196][2] +
                mat_A[238][1] * mat_B[204][2] +
                mat_A[238][2] * mat_B[212][2] +
                mat_A[238][3] * mat_B[220][2] +
                mat_A[239][0] * mat_B[228][2] +
                mat_A[239][1] * mat_B[236][2] +
                mat_A[239][2] * mat_B[244][2] +
                mat_A[239][3] * mat_B[252][2];
    mat_C[236][3] <=
                mat_A[232][0] * mat_B[4][3] +
                mat_A[232][1] * mat_B[12][3] +
                mat_A[232][2] * mat_B[20][3] +
                mat_A[232][3] * mat_B[28][3] +
                mat_A[233][0] * mat_B[36][3] +
                mat_A[233][1] * mat_B[44][3] +
                mat_A[233][2] * mat_B[52][3] +
                mat_A[233][3] * mat_B[60][3] +
                mat_A[234][0] * mat_B[68][3] +
                mat_A[234][1] * mat_B[76][3] +
                mat_A[234][2] * mat_B[84][3] +
                mat_A[234][3] * mat_B[92][3] +
                mat_A[235][0] * mat_B[100][3] +
                mat_A[235][1] * mat_B[108][3] +
                mat_A[235][2] * mat_B[116][3] +
                mat_A[235][3] * mat_B[124][3] +
                mat_A[236][0] * mat_B[132][3] +
                mat_A[236][1] * mat_B[140][3] +
                mat_A[236][2] * mat_B[148][3] +
                mat_A[236][3] * mat_B[156][3] +
                mat_A[237][0] * mat_B[164][3] +
                mat_A[237][1] * mat_B[172][3] +
                mat_A[237][2] * mat_B[180][3] +
                mat_A[237][3] * mat_B[188][3] +
                mat_A[238][0] * mat_B[196][3] +
                mat_A[238][1] * mat_B[204][3] +
                mat_A[238][2] * mat_B[212][3] +
                mat_A[238][3] * mat_B[220][3] +
                mat_A[239][0] * mat_B[228][3] +
                mat_A[239][1] * mat_B[236][3] +
                mat_A[239][2] * mat_B[244][3] +
                mat_A[239][3] * mat_B[252][3];
    mat_C[237][0] <=
                mat_A[232][0] * mat_B[5][0] +
                mat_A[232][1] * mat_B[13][0] +
                mat_A[232][2] * mat_B[21][0] +
                mat_A[232][3] * mat_B[29][0] +
                mat_A[233][0] * mat_B[37][0] +
                mat_A[233][1] * mat_B[45][0] +
                mat_A[233][2] * mat_B[53][0] +
                mat_A[233][3] * mat_B[61][0] +
                mat_A[234][0] * mat_B[69][0] +
                mat_A[234][1] * mat_B[77][0] +
                mat_A[234][2] * mat_B[85][0] +
                mat_A[234][3] * mat_B[93][0] +
                mat_A[235][0] * mat_B[101][0] +
                mat_A[235][1] * mat_B[109][0] +
                mat_A[235][2] * mat_B[117][0] +
                mat_A[235][3] * mat_B[125][0] +
                mat_A[236][0] * mat_B[133][0] +
                mat_A[236][1] * mat_B[141][0] +
                mat_A[236][2] * mat_B[149][0] +
                mat_A[236][3] * mat_B[157][0] +
                mat_A[237][0] * mat_B[165][0] +
                mat_A[237][1] * mat_B[173][0] +
                mat_A[237][2] * mat_B[181][0] +
                mat_A[237][3] * mat_B[189][0] +
                mat_A[238][0] * mat_B[197][0] +
                mat_A[238][1] * mat_B[205][0] +
                mat_A[238][2] * mat_B[213][0] +
                mat_A[238][3] * mat_B[221][0] +
                mat_A[239][0] * mat_B[229][0] +
                mat_A[239][1] * mat_B[237][0] +
                mat_A[239][2] * mat_B[245][0] +
                mat_A[239][3] * mat_B[253][0];
    mat_C[237][1] <=
                mat_A[232][0] * mat_B[5][1] +
                mat_A[232][1] * mat_B[13][1] +
                mat_A[232][2] * mat_B[21][1] +
                mat_A[232][3] * mat_B[29][1] +
                mat_A[233][0] * mat_B[37][1] +
                mat_A[233][1] * mat_B[45][1] +
                mat_A[233][2] * mat_B[53][1] +
                mat_A[233][3] * mat_B[61][1] +
                mat_A[234][0] * mat_B[69][1] +
                mat_A[234][1] * mat_B[77][1] +
                mat_A[234][2] * mat_B[85][1] +
                mat_A[234][3] * mat_B[93][1] +
                mat_A[235][0] * mat_B[101][1] +
                mat_A[235][1] * mat_B[109][1] +
                mat_A[235][2] * mat_B[117][1] +
                mat_A[235][3] * mat_B[125][1] +
                mat_A[236][0] * mat_B[133][1] +
                mat_A[236][1] * mat_B[141][1] +
                mat_A[236][2] * mat_B[149][1] +
                mat_A[236][3] * mat_B[157][1] +
                mat_A[237][0] * mat_B[165][1] +
                mat_A[237][1] * mat_B[173][1] +
                mat_A[237][2] * mat_B[181][1] +
                mat_A[237][3] * mat_B[189][1] +
                mat_A[238][0] * mat_B[197][1] +
                mat_A[238][1] * mat_B[205][1] +
                mat_A[238][2] * mat_B[213][1] +
                mat_A[238][3] * mat_B[221][1] +
                mat_A[239][0] * mat_B[229][1] +
                mat_A[239][1] * mat_B[237][1] +
                mat_A[239][2] * mat_B[245][1] +
                mat_A[239][3] * mat_B[253][1];
    mat_C[237][2] <=
                mat_A[232][0] * mat_B[5][2] +
                mat_A[232][1] * mat_B[13][2] +
                mat_A[232][2] * mat_B[21][2] +
                mat_A[232][3] * mat_B[29][2] +
                mat_A[233][0] * mat_B[37][2] +
                mat_A[233][1] * mat_B[45][2] +
                mat_A[233][2] * mat_B[53][2] +
                mat_A[233][3] * mat_B[61][2] +
                mat_A[234][0] * mat_B[69][2] +
                mat_A[234][1] * mat_B[77][2] +
                mat_A[234][2] * mat_B[85][2] +
                mat_A[234][3] * mat_B[93][2] +
                mat_A[235][0] * mat_B[101][2] +
                mat_A[235][1] * mat_B[109][2] +
                mat_A[235][2] * mat_B[117][2] +
                mat_A[235][3] * mat_B[125][2] +
                mat_A[236][0] * mat_B[133][2] +
                mat_A[236][1] * mat_B[141][2] +
                mat_A[236][2] * mat_B[149][2] +
                mat_A[236][3] * mat_B[157][2] +
                mat_A[237][0] * mat_B[165][2] +
                mat_A[237][1] * mat_B[173][2] +
                mat_A[237][2] * mat_B[181][2] +
                mat_A[237][3] * mat_B[189][2] +
                mat_A[238][0] * mat_B[197][2] +
                mat_A[238][1] * mat_B[205][2] +
                mat_A[238][2] * mat_B[213][2] +
                mat_A[238][3] * mat_B[221][2] +
                mat_A[239][0] * mat_B[229][2] +
                mat_A[239][1] * mat_B[237][2] +
                mat_A[239][2] * mat_B[245][2] +
                mat_A[239][3] * mat_B[253][2];
    mat_C[237][3] <=
                mat_A[232][0] * mat_B[5][3] +
                mat_A[232][1] * mat_B[13][3] +
                mat_A[232][2] * mat_B[21][3] +
                mat_A[232][3] * mat_B[29][3] +
                mat_A[233][0] * mat_B[37][3] +
                mat_A[233][1] * mat_B[45][3] +
                mat_A[233][2] * mat_B[53][3] +
                mat_A[233][3] * mat_B[61][3] +
                mat_A[234][0] * mat_B[69][3] +
                mat_A[234][1] * mat_B[77][3] +
                mat_A[234][2] * mat_B[85][3] +
                mat_A[234][3] * mat_B[93][3] +
                mat_A[235][0] * mat_B[101][3] +
                mat_A[235][1] * mat_B[109][3] +
                mat_A[235][2] * mat_B[117][3] +
                mat_A[235][3] * mat_B[125][3] +
                mat_A[236][0] * mat_B[133][3] +
                mat_A[236][1] * mat_B[141][3] +
                mat_A[236][2] * mat_B[149][3] +
                mat_A[236][3] * mat_B[157][3] +
                mat_A[237][0] * mat_B[165][3] +
                mat_A[237][1] * mat_B[173][3] +
                mat_A[237][2] * mat_B[181][3] +
                mat_A[237][3] * mat_B[189][3] +
                mat_A[238][0] * mat_B[197][3] +
                mat_A[238][1] * mat_B[205][3] +
                mat_A[238][2] * mat_B[213][3] +
                mat_A[238][3] * mat_B[221][3] +
                mat_A[239][0] * mat_B[229][3] +
                mat_A[239][1] * mat_B[237][3] +
                mat_A[239][2] * mat_B[245][3] +
                mat_A[239][3] * mat_B[253][3];
    mat_C[238][0] <=
                mat_A[232][0] * mat_B[6][0] +
                mat_A[232][1] * mat_B[14][0] +
                mat_A[232][2] * mat_B[22][0] +
                mat_A[232][3] * mat_B[30][0] +
                mat_A[233][0] * mat_B[38][0] +
                mat_A[233][1] * mat_B[46][0] +
                mat_A[233][2] * mat_B[54][0] +
                mat_A[233][3] * mat_B[62][0] +
                mat_A[234][0] * mat_B[70][0] +
                mat_A[234][1] * mat_B[78][0] +
                mat_A[234][2] * mat_B[86][0] +
                mat_A[234][3] * mat_B[94][0] +
                mat_A[235][0] * mat_B[102][0] +
                mat_A[235][1] * mat_B[110][0] +
                mat_A[235][2] * mat_B[118][0] +
                mat_A[235][3] * mat_B[126][0] +
                mat_A[236][0] * mat_B[134][0] +
                mat_A[236][1] * mat_B[142][0] +
                mat_A[236][2] * mat_B[150][0] +
                mat_A[236][3] * mat_B[158][0] +
                mat_A[237][0] * mat_B[166][0] +
                mat_A[237][1] * mat_B[174][0] +
                mat_A[237][2] * mat_B[182][0] +
                mat_A[237][3] * mat_B[190][0] +
                mat_A[238][0] * mat_B[198][0] +
                mat_A[238][1] * mat_B[206][0] +
                mat_A[238][2] * mat_B[214][0] +
                mat_A[238][3] * mat_B[222][0] +
                mat_A[239][0] * mat_B[230][0] +
                mat_A[239][1] * mat_B[238][0] +
                mat_A[239][2] * mat_B[246][0] +
                mat_A[239][3] * mat_B[254][0];
    mat_C[238][1] <=
                mat_A[232][0] * mat_B[6][1] +
                mat_A[232][1] * mat_B[14][1] +
                mat_A[232][2] * mat_B[22][1] +
                mat_A[232][3] * mat_B[30][1] +
                mat_A[233][0] * mat_B[38][1] +
                mat_A[233][1] * mat_B[46][1] +
                mat_A[233][2] * mat_B[54][1] +
                mat_A[233][3] * mat_B[62][1] +
                mat_A[234][0] * mat_B[70][1] +
                mat_A[234][1] * mat_B[78][1] +
                mat_A[234][2] * mat_B[86][1] +
                mat_A[234][3] * mat_B[94][1] +
                mat_A[235][0] * mat_B[102][1] +
                mat_A[235][1] * mat_B[110][1] +
                mat_A[235][2] * mat_B[118][1] +
                mat_A[235][3] * mat_B[126][1] +
                mat_A[236][0] * mat_B[134][1] +
                mat_A[236][1] * mat_B[142][1] +
                mat_A[236][2] * mat_B[150][1] +
                mat_A[236][3] * mat_B[158][1] +
                mat_A[237][0] * mat_B[166][1] +
                mat_A[237][1] * mat_B[174][1] +
                mat_A[237][2] * mat_B[182][1] +
                mat_A[237][3] * mat_B[190][1] +
                mat_A[238][0] * mat_B[198][1] +
                mat_A[238][1] * mat_B[206][1] +
                mat_A[238][2] * mat_B[214][1] +
                mat_A[238][3] * mat_B[222][1] +
                mat_A[239][0] * mat_B[230][1] +
                mat_A[239][1] * mat_B[238][1] +
                mat_A[239][2] * mat_B[246][1] +
                mat_A[239][3] * mat_B[254][1];
    mat_C[238][2] <=
                mat_A[232][0] * mat_B[6][2] +
                mat_A[232][1] * mat_B[14][2] +
                mat_A[232][2] * mat_B[22][2] +
                mat_A[232][3] * mat_B[30][2] +
                mat_A[233][0] * mat_B[38][2] +
                mat_A[233][1] * mat_B[46][2] +
                mat_A[233][2] * mat_B[54][2] +
                mat_A[233][3] * mat_B[62][2] +
                mat_A[234][0] * mat_B[70][2] +
                mat_A[234][1] * mat_B[78][2] +
                mat_A[234][2] * mat_B[86][2] +
                mat_A[234][3] * mat_B[94][2] +
                mat_A[235][0] * mat_B[102][2] +
                mat_A[235][1] * mat_B[110][2] +
                mat_A[235][2] * mat_B[118][2] +
                mat_A[235][3] * mat_B[126][2] +
                mat_A[236][0] * mat_B[134][2] +
                mat_A[236][1] * mat_B[142][2] +
                mat_A[236][2] * mat_B[150][2] +
                mat_A[236][3] * mat_B[158][2] +
                mat_A[237][0] * mat_B[166][2] +
                mat_A[237][1] * mat_B[174][2] +
                mat_A[237][2] * mat_B[182][2] +
                mat_A[237][3] * mat_B[190][2] +
                mat_A[238][0] * mat_B[198][2] +
                mat_A[238][1] * mat_B[206][2] +
                mat_A[238][2] * mat_B[214][2] +
                mat_A[238][3] * mat_B[222][2] +
                mat_A[239][0] * mat_B[230][2] +
                mat_A[239][1] * mat_B[238][2] +
                mat_A[239][2] * mat_B[246][2] +
                mat_A[239][3] * mat_B[254][2];
    mat_C[238][3] <=
                mat_A[232][0] * mat_B[6][3] +
                mat_A[232][1] * mat_B[14][3] +
                mat_A[232][2] * mat_B[22][3] +
                mat_A[232][3] * mat_B[30][3] +
                mat_A[233][0] * mat_B[38][3] +
                mat_A[233][1] * mat_B[46][3] +
                mat_A[233][2] * mat_B[54][3] +
                mat_A[233][3] * mat_B[62][3] +
                mat_A[234][0] * mat_B[70][3] +
                mat_A[234][1] * mat_B[78][3] +
                mat_A[234][2] * mat_B[86][3] +
                mat_A[234][3] * mat_B[94][3] +
                mat_A[235][0] * mat_B[102][3] +
                mat_A[235][1] * mat_B[110][3] +
                mat_A[235][2] * mat_B[118][3] +
                mat_A[235][3] * mat_B[126][3] +
                mat_A[236][0] * mat_B[134][3] +
                mat_A[236][1] * mat_B[142][3] +
                mat_A[236][2] * mat_B[150][3] +
                mat_A[236][3] * mat_B[158][3] +
                mat_A[237][0] * mat_B[166][3] +
                mat_A[237][1] * mat_B[174][3] +
                mat_A[237][2] * mat_B[182][3] +
                mat_A[237][3] * mat_B[190][3] +
                mat_A[238][0] * mat_B[198][3] +
                mat_A[238][1] * mat_B[206][3] +
                mat_A[238][2] * mat_B[214][3] +
                mat_A[238][3] * mat_B[222][3] +
                mat_A[239][0] * mat_B[230][3] +
                mat_A[239][1] * mat_B[238][3] +
                mat_A[239][2] * mat_B[246][3] +
                mat_A[239][3] * mat_B[254][3];
    mat_C[239][0] <=
                mat_A[232][0] * mat_B[7][0] +
                mat_A[232][1] * mat_B[15][0] +
                mat_A[232][2] * mat_B[23][0] +
                mat_A[232][3] * mat_B[31][0] +
                mat_A[233][0] * mat_B[39][0] +
                mat_A[233][1] * mat_B[47][0] +
                mat_A[233][2] * mat_B[55][0] +
                mat_A[233][3] * mat_B[63][0] +
                mat_A[234][0] * mat_B[71][0] +
                mat_A[234][1] * mat_B[79][0] +
                mat_A[234][2] * mat_B[87][0] +
                mat_A[234][3] * mat_B[95][0] +
                mat_A[235][0] * mat_B[103][0] +
                mat_A[235][1] * mat_B[111][0] +
                mat_A[235][2] * mat_B[119][0] +
                mat_A[235][3] * mat_B[127][0] +
                mat_A[236][0] * mat_B[135][0] +
                mat_A[236][1] * mat_B[143][0] +
                mat_A[236][2] * mat_B[151][0] +
                mat_A[236][3] * mat_B[159][0] +
                mat_A[237][0] * mat_B[167][0] +
                mat_A[237][1] * mat_B[175][0] +
                mat_A[237][2] * mat_B[183][0] +
                mat_A[237][3] * mat_B[191][0] +
                mat_A[238][0] * mat_B[199][0] +
                mat_A[238][1] * mat_B[207][0] +
                mat_A[238][2] * mat_B[215][0] +
                mat_A[238][3] * mat_B[223][0] +
                mat_A[239][0] * mat_B[231][0] +
                mat_A[239][1] * mat_B[239][0] +
                mat_A[239][2] * mat_B[247][0] +
                mat_A[239][3] * mat_B[255][0];
    mat_C[239][1] <=
                mat_A[232][0] * mat_B[7][1] +
                mat_A[232][1] * mat_B[15][1] +
                mat_A[232][2] * mat_B[23][1] +
                mat_A[232][3] * mat_B[31][1] +
                mat_A[233][0] * mat_B[39][1] +
                mat_A[233][1] * mat_B[47][1] +
                mat_A[233][2] * mat_B[55][1] +
                mat_A[233][3] * mat_B[63][1] +
                mat_A[234][0] * mat_B[71][1] +
                mat_A[234][1] * mat_B[79][1] +
                mat_A[234][2] * mat_B[87][1] +
                mat_A[234][3] * mat_B[95][1] +
                mat_A[235][0] * mat_B[103][1] +
                mat_A[235][1] * mat_B[111][1] +
                mat_A[235][2] * mat_B[119][1] +
                mat_A[235][3] * mat_B[127][1] +
                mat_A[236][0] * mat_B[135][1] +
                mat_A[236][1] * mat_B[143][1] +
                mat_A[236][2] * mat_B[151][1] +
                mat_A[236][3] * mat_B[159][1] +
                mat_A[237][0] * mat_B[167][1] +
                mat_A[237][1] * mat_B[175][1] +
                mat_A[237][2] * mat_B[183][1] +
                mat_A[237][3] * mat_B[191][1] +
                mat_A[238][0] * mat_B[199][1] +
                mat_A[238][1] * mat_B[207][1] +
                mat_A[238][2] * mat_B[215][1] +
                mat_A[238][3] * mat_B[223][1] +
                mat_A[239][0] * mat_B[231][1] +
                mat_A[239][1] * mat_B[239][1] +
                mat_A[239][2] * mat_B[247][1] +
                mat_A[239][3] * mat_B[255][1];
    mat_C[239][2] <=
                mat_A[232][0] * mat_B[7][2] +
                mat_A[232][1] * mat_B[15][2] +
                mat_A[232][2] * mat_B[23][2] +
                mat_A[232][3] * mat_B[31][2] +
                mat_A[233][0] * mat_B[39][2] +
                mat_A[233][1] * mat_B[47][2] +
                mat_A[233][2] * mat_B[55][2] +
                mat_A[233][3] * mat_B[63][2] +
                mat_A[234][0] * mat_B[71][2] +
                mat_A[234][1] * mat_B[79][2] +
                mat_A[234][2] * mat_B[87][2] +
                mat_A[234][3] * mat_B[95][2] +
                mat_A[235][0] * mat_B[103][2] +
                mat_A[235][1] * mat_B[111][2] +
                mat_A[235][2] * mat_B[119][2] +
                mat_A[235][3] * mat_B[127][2] +
                mat_A[236][0] * mat_B[135][2] +
                mat_A[236][1] * mat_B[143][2] +
                mat_A[236][2] * mat_B[151][2] +
                mat_A[236][3] * mat_B[159][2] +
                mat_A[237][0] * mat_B[167][2] +
                mat_A[237][1] * mat_B[175][2] +
                mat_A[237][2] * mat_B[183][2] +
                mat_A[237][3] * mat_B[191][2] +
                mat_A[238][0] * mat_B[199][2] +
                mat_A[238][1] * mat_B[207][2] +
                mat_A[238][2] * mat_B[215][2] +
                mat_A[238][3] * mat_B[223][2] +
                mat_A[239][0] * mat_B[231][2] +
                mat_A[239][1] * mat_B[239][2] +
                mat_A[239][2] * mat_B[247][2] +
                mat_A[239][3] * mat_B[255][2];
    mat_C[239][3] <=
                mat_A[232][0] * mat_B[7][3] +
                mat_A[232][1] * mat_B[15][3] +
                mat_A[232][2] * mat_B[23][3] +
                mat_A[232][3] * mat_B[31][3] +
                mat_A[233][0] * mat_B[39][3] +
                mat_A[233][1] * mat_B[47][3] +
                mat_A[233][2] * mat_B[55][3] +
                mat_A[233][3] * mat_B[63][3] +
                mat_A[234][0] * mat_B[71][3] +
                mat_A[234][1] * mat_B[79][3] +
                mat_A[234][2] * mat_B[87][3] +
                mat_A[234][3] * mat_B[95][3] +
                mat_A[235][0] * mat_B[103][3] +
                mat_A[235][1] * mat_B[111][3] +
                mat_A[235][2] * mat_B[119][3] +
                mat_A[235][3] * mat_B[127][3] +
                mat_A[236][0] * mat_B[135][3] +
                mat_A[236][1] * mat_B[143][3] +
                mat_A[236][2] * mat_B[151][3] +
                mat_A[236][3] * mat_B[159][3] +
                mat_A[237][0] * mat_B[167][3] +
                mat_A[237][1] * mat_B[175][3] +
                mat_A[237][2] * mat_B[183][3] +
                mat_A[237][3] * mat_B[191][3] +
                mat_A[238][0] * mat_B[199][3] +
                mat_A[238][1] * mat_B[207][3] +
                mat_A[238][2] * mat_B[215][3] +
                mat_A[238][3] * mat_B[223][3] +
                mat_A[239][0] * mat_B[231][3] +
                mat_A[239][1] * mat_B[239][3] +
                mat_A[239][2] * mat_B[247][3] +
                mat_A[239][3] * mat_B[255][3];
    mat_C[240][0] <=
                mat_A[240][0] * mat_B[0][0] +
                mat_A[240][1] * mat_B[8][0] +
                mat_A[240][2] * mat_B[16][0] +
                mat_A[240][3] * mat_B[24][0] +
                mat_A[241][0] * mat_B[32][0] +
                mat_A[241][1] * mat_B[40][0] +
                mat_A[241][2] * mat_B[48][0] +
                mat_A[241][3] * mat_B[56][0] +
                mat_A[242][0] * mat_B[64][0] +
                mat_A[242][1] * mat_B[72][0] +
                mat_A[242][2] * mat_B[80][0] +
                mat_A[242][3] * mat_B[88][0] +
                mat_A[243][0] * mat_B[96][0] +
                mat_A[243][1] * mat_B[104][0] +
                mat_A[243][2] * mat_B[112][0] +
                mat_A[243][3] * mat_B[120][0] +
                mat_A[244][0] * mat_B[128][0] +
                mat_A[244][1] * mat_B[136][0] +
                mat_A[244][2] * mat_B[144][0] +
                mat_A[244][3] * mat_B[152][0] +
                mat_A[245][0] * mat_B[160][0] +
                mat_A[245][1] * mat_B[168][0] +
                mat_A[245][2] * mat_B[176][0] +
                mat_A[245][3] * mat_B[184][0] +
                mat_A[246][0] * mat_B[192][0] +
                mat_A[246][1] * mat_B[200][0] +
                mat_A[246][2] * mat_B[208][0] +
                mat_A[246][3] * mat_B[216][0] +
                mat_A[247][0] * mat_B[224][0] +
                mat_A[247][1] * mat_B[232][0] +
                mat_A[247][2] * mat_B[240][0] +
                mat_A[247][3] * mat_B[248][0];
    mat_C[240][1] <=
                mat_A[240][0] * mat_B[0][1] +
                mat_A[240][1] * mat_B[8][1] +
                mat_A[240][2] * mat_B[16][1] +
                mat_A[240][3] * mat_B[24][1] +
                mat_A[241][0] * mat_B[32][1] +
                mat_A[241][1] * mat_B[40][1] +
                mat_A[241][2] * mat_B[48][1] +
                mat_A[241][3] * mat_B[56][1] +
                mat_A[242][0] * mat_B[64][1] +
                mat_A[242][1] * mat_B[72][1] +
                mat_A[242][2] * mat_B[80][1] +
                mat_A[242][3] * mat_B[88][1] +
                mat_A[243][0] * mat_B[96][1] +
                mat_A[243][1] * mat_B[104][1] +
                mat_A[243][2] * mat_B[112][1] +
                mat_A[243][3] * mat_B[120][1] +
                mat_A[244][0] * mat_B[128][1] +
                mat_A[244][1] * mat_B[136][1] +
                mat_A[244][2] * mat_B[144][1] +
                mat_A[244][3] * mat_B[152][1] +
                mat_A[245][0] * mat_B[160][1] +
                mat_A[245][1] * mat_B[168][1] +
                mat_A[245][2] * mat_B[176][1] +
                mat_A[245][3] * mat_B[184][1] +
                mat_A[246][0] * mat_B[192][1] +
                mat_A[246][1] * mat_B[200][1] +
                mat_A[246][2] * mat_B[208][1] +
                mat_A[246][3] * mat_B[216][1] +
                mat_A[247][0] * mat_B[224][1] +
                mat_A[247][1] * mat_B[232][1] +
                mat_A[247][2] * mat_B[240][1] +
                mat_A[247][3] * mat_B[248][1];
    mat_C[240][2] <=
                mat_A[240][0] * mat_B[0][2] +
                mat_A[240][1] * mat_B[8][2] +
                mat_A[240][2] * mat_B[16][2] +
                mat_A[240][3] * mat_B[24][2] +
                mat_A[241][0] * mat_B[32][2] +
                mat_A[241][1] * mat_B[40][2] +
                mat_A[241][2] * mat_B[48][2] +
                mat_A[241][3] * mat_B[56][2] +
                mat_A[242][0] * mat_B[64][2] +
                mat_A[242][1] * mat_B[72][2] +
                mat_A[242][2] * mat_B[80][2] +
                mat_A[242][3] * mat_B[88][2] +
                mat_A[243][0] * mat_B[96][2] +
                mat_A[243][1] * mat_B[104][2] +
                mat_A[243][2] * mat_B[112][2] +
                mat_A[243][3] * mat_B[120][2] +
                mat_A[244][0] * mat_B[128][2] +
                mat_A[244][1] * mat_B[136][2] +
                mat_A[244][2] * mat_B[144][2] +
                mat_A[244][3] * mat_B[152][2] +
                mat_A[245][0] * mat_B[160][2] +
                mat_A[245][1] * mat_B[168][2] +
                mat_A[245][2] * mat_B[176][2] +
                mat_A[245][3] * mat_B[184][2] +
                mat_A[246][0] * mat_B[192][2] +
                mat_A[246][1] * mat_B[200][2] +
                mat_A[246][2] * mat_B[208][2] +
                mat_A[246][3] * mat_B[216][2] +
                mat_A[247][0] * mat_B[224][2] +
                mat_A[247][1] * mat_B[232][2] +
                mat_A[247][2] * mat_B[240][2] +
                mat_A[247][3] * mat_B[248][2];
    mat_C[240][3] <=
                mat_A[240][0] * mat_B[0][3] +
                mat_A[240][1] * mat_B[8][3] +
                mat_A[240][2] * mat_B[16][3] +
                mat_A[240][3] * mat_B[24][3] +
                mat_A[241][0] * mat_B[32][3] +
                mat_A[241][1] * mat_B[40][3] +
                mat_A[241][2] * mat_B[48][3] +
                mat_A[241][3] * mat_B[56][3] +
                mat_A[242][0] * mat_B[64][3] +
                mat_A[242][1] * mat_B[72][3] +
                mat_A[242][2] * mat_B[80][3] +
                mat_A[242][3] * mat_B[88][3] +
                mat_A[243][0] * mat_B[96][3] +
                mat_A[243][1] * mat_B[104][3] +
                mat_A[243][2] * mat_B[112][3] +
                mat_A[243][3] * mat_B[120][3] +
                mat_A[244][0] * mat_B[128][3] +
                mat_A[244][1] * mat_B[136][3] +
                mat_A[244][2] * mat_B[144][3] +
                mat_A[244][3] * mat_B[152][3] +
                mat_A[245][0] * mat_B[160][3] +
                mat_A[245][1] * mat_B[168][3] +
                mat_A[245][2] * mat_B[176][3] +
                mat_A[245][3] * mat_B[184][3] +
                mat_A[246][0] * mat_B[192][3] +
                mat_A[246][1] * mat_B[200][3] +
                mat_A[246][2] * mat_B[208][3] +
                mat_A[246][3] * mat_B[216][3] +
                mat_A[247][0] * mat_B[224][3] +
                mat_A[247][1] * mat_B[232][3] +
                mat_A[247][2] * mat_B[240][3] +
                mat_A[247][3] * mat_B[248][3];
    mat_C[241][0] <=
                mat_A[240][0] * mat_B[1][0] +
                mat_A[240][1] * mat_B[9][0] +
                mat_A[240][2] * mat_B[17][0] +
                mat_A[240][3] * mat_B[25][0] +
                mat_A[241][0] * mat_B[33][0] +
                mat_A[241][1] * mat_B[41][0] +
                mat_A[241][2] * mat_B[49][0] +
                mat_A[241][3] * mat_B[57][0] +
                mat_A[242][0] * mat_B[65][0] +
                mat_A[242][1] * mat_B[73][0] +
                mat_A[242][2] * mat_B[81][0] +
                mat_A[242][3] * mat_B[89][0] +
                mat_A[243][0] * mat_B[97][0] +
                mat_A[243][1] * mat_B[105][0] +
                mat_A[243][2] * mat_B[113][0] +
                mat_A[243][3] * mat_B[121][0] +
                mat_A[244][0] * mat_B[129][0] +
                mat_A[244][1] * mat_B[137][0] +
                mat_A[244][2] * mat_B[145][0] +
                mat_A[244][3] * mat_B[153][0] +
                mat_A[245][0] * mat_B[161][0] +
                mat_A[245][1] * mat_B[169][0] +
                mat_A[245][2] * mat_B[177][0] +
                mat_A[245][3] * mat_B[185][0] +
                mat_A[246][0] * mat_B[193][0] +
                mat_A[246][1] * mat_B[201][0] +
                mat_A[246][2] * mat_B[209][0] +
                mat_A[246][3] * mat_B[217][0] +
                mat_A[247][0] * mat_B[225][0] +
                mat_A[247][1] * mat_B[233][0] +
                mat_A[247][2] * mat_B[241][0] +
                mat_A[247][3] * mat_B[249][0];
    mat_C[241][1] <=
                mat_A[240][0] * mat_B[1][1] +
                mat_A[240][1] * mat_B[9][1] +
                mat_A[240][2] * mat_B[17][1] +
                mat_A[240][3] * mat_B[25][1] +
                mat_A[241][0] * mat_B[33][1] +
                mat_A[241][1] * mat_B[41][1] +
                mat_A[241][2] * mat_B[49][1] +
                mat_A[241][3] * mat_B[57][1] +
                mat_A[242][0] * mat_B[65][1] +
                mat_A[242][1] * mat_B[73][1] +
                mat_A[242][2] * mat_B[81][1] +
                mat_A[242][3] * mat_B[89][1] +
                mat_A[243][0] * mat_B[97][1] +
                mat_A[243][1] * mat_B[105][1] +
                mat_A[243][2] * mat_B[113][1] +
                mat_A[243][3] * mat_B[121][1] +
                mat_A[244][0] * mat_B[129][1] +
                mat_A[244][1] * mat_B[137][1] +
                mat_A[244][2] * mat_B[145][1] +
                mat_A[244][3] * mat_B[153][1] +
                mat_A[245][0] * mat_B[161][1] +
                mat_A[245][1] * mat_B[169][1] +
                mat_A[245][2] * mat_B[177][1] +
                mat_A[245][3] * mat_B[185][1] +
                mat_A[246][0] * mat_B[193][1] +
                mat_A[246][1] * mat_B[201][1] +
                mat_A[246][2] * mat_B[209][1] +
                mat_A[246][3] * mat_B[217][1] +
                mat_A[247][0] * mat_B[225][1] +
                mat_A[247][1] * mat_B[233][1] +
                mat_A[247][2] * mat_B[241][1] +
                mat_A[247][3] * mat_B[249][1];
    mat_C[241][2] <=
                mat_A[240][0] * mat_B[1][2] +
                mat_A[240][1] * mat_B[9][2] +
                mat_A[240][2] * mat_B[17][2] +
                mat_A[240][3] * mat_B[25][2] +
                mat_A[241][0] * mat_B[33][2] +
                mat_A[241][1] * mat_B[41][2] +
                mat_A[241][2] * mat_B[49][2] +
                mat_A[241][3] * mat_B[57][2] +
                mat_A[242][0] * mat_B[65][2] +
                mat_A[242][1] * mat_B[73][2] +
                mat_A[242][2] * mat_B[81][2] +
                mat_A[242][3] * mat_B[89][2] +
                mat_A[243][0] * mat_B[97][2] +
                mat_A[243][1] * mat_B[105][2] +
                mat_A[243][2] * mat_B[113][2] +
                mat_A[243][3] * mat_B[121][2] +
                mat_A[244][0] * mat_B[129][2] +
                mat_A[244][1] * mat_B[137][2] +
                mat_A[244][2] * mat_B[145][2] +
                mat_A[244][3] * mat_B[153][2] +
                mat_A[245][0] * mat_B[161][2] +
                mat_A[245][1] * mat_B[169][2] +
                mat_A[245][2] * mat_B[177][2] +
                mat_A[245][3] * mat_B[185][2] +
                mat_A[246][0] * mat_B[193][2] +
                mat_A[246][1] * mat_B[201][2] +
                mat_A[246][2] * mat_B[209][2] +
                mat_A[246][3] * mat_B[217][2] +
                mat_A[247][0] * mat_B[225][2] +
                mat_A[247][1] * mat_B[233][2] +
                mat_A[247][2] * mat_B[241][2] +
                mat_A[247][3] * mat_B[249][2];
    mat_C[241][3] <=
                mat_A[240][0] * mat_B[1][3] +
                mat_A[240][1] * mat_B[9][3] +
                mat_A[240][2] * mat_B[17][3] +
                mat_A[240][3] * mat_B[25][3] +
                mat_A[241][0] * mat_B[33][3] +
                mat_A[241][1] * mat_B[41][3] +
                mat_A[241][2] * mat_B[49][3] +
                mat_A[241][3] * mat_B[57][3] +
                mat_A[242][0] * mat_B[65][3] +
                mat_A[242][1] * mat_B[73][3] +
                mat_A[242][2] * mat_B[81][3] +
                mat_A[242][3] * mat_B[89][3] +
                mat_A[243][0] * mat_B[97][3] +
                mat_A[243][1] * mat_B[105][3] +
                mat_A[243][2] * mat_B[113][3] +
                mat_A[243][3] * mat_B[121][3] +
                mat_A[244][0] * mat_B[129][3] +
                mat_A[244][1] * mat_B[137][3] +
                mat_A[244][2] * mat_B[145][3] +
                mat_A[244][3] * mat_B[153][3] +
                mat_A[245][0] * mat_B[161][3] +
                mat_A[245][1] * mat_B[169][3] +
                mat_A[245][2] * mat_B[177][3] +
                mat_A[245][3] * mat_B[185][3] +
                mat_A[246][0] * mat_B[193][3] +
                mat_A[246][1] * mat_B[201][3] +
                mat_A[246][2] * mat_B[209][3] +
                mat_A[246][3] * mat_B[217][3] +
                mat_A[247][0] * mat_B[225][3] +
                mat_A[247][1] * mat_B[233][3] +
                mat_A[247][2] * mat_B[241][3] +
                mat_A[247][3] * mat_B[249][3];
    mat_C[242][0] <=
                mat_A[240][0] * mat_B[2][0] +
                mat_A[240][1] * mat_B[10][0] +
                mat_A[240][2] * mat_B[18][0] +
                mat_A[240][3] * mat_B[26][0] +
                mat_A[241][0] * mat_B[34][0] +
                mat_A[241][1] * mat_B[42][0] +
                mat_A[241][2] * mat_B[50][0] +
                mat_A[241][3] * mat_B[58][0] +
                mat_A[242][0] * mat_B[66][0] +
                mat_A[242][1] * mat_B[74][0] +
                mat_A[242][2] * mat_B[82][0] +
                mat_A[242][3] * mat_B[90][0] +
                mat_A[243][0] * mat_B[98][0] +
                mat_A[243][1] * mat_B[106][0] +
                mat_A[243][2] * mat_B[114][0] +
                mat_A[243][3] * mat_B[122][0] +
                mat_A[244][0] * mat_B[130][0] +
                mat_A[244][1] * mat_B[138][0] +
                mat_A[244][2] * mat_B[146][0] +
                mat_A[244][3] * mat_B[154][0] +
                mat_A[245][0] * mat_B[162][0] +
                mat_A[245][1] * mat_B[170][0] +
                mat_A[245][2] * mat_B[178][0] +
                mat_A[245][3] * mat_B[186][0] +
                mat_A[246][0] * mat_B[194][0] +
                mat_A[246][1] * mat_B[202][0] +
                mat_A[246][2] * mat_B[210][0] +
                mat_A[246][3] * mat_B[218][0] +
                mat_A[247][0] * mat_B[226][0] +
                mat_A[247][1] * mat_B[234][0] +
                mat_A[247][2] * mat_B[242][0] +
                mat_A[247][3] * mat_B[250][0];
    mat_C[242][1] <=
                mat_A[240][0] * mat_B[2][1] +
                mat_A[240][1] * mat_B[10][1] +
                mat_A[240][2] * mat_B[18][1] +
                mat_A[240][3] * mat_B[26][1] +
                mat_A[241][0] * mat_B[34][1] +
                mat_A[241][1] * mat_B[42][1] +
                mat_A[241][2] * mat_B[50][1] +
                mat_A[241][3] * mat_B[58][1] +
                mat_A[242][0] * mat_B[66][1] +
                mat_A[242][1] * mat_B[74][1] +
                mat_A[242][2] * mat_B[82][1] +
                mat_A[242][3] * mat_B[90][1] +
                mat_A[243][0] * mat_B[98][1] +
                mat_A[243][1] * mat_B[106][1] +
                mat_A[243][2] * mat_B[114][1] +
                mat_A[243][3] * mat_B[122][1] +
                mat_A[244][0] * mat_B[130][1] +
                mat_A[244][1] * mat_B[138][1] +
                mat_A[244][2] * mat_B[146][1] +
                mat_A[244][3] * mat_B[154][1] +
                mat_A[245][0] * mat_B[162][1] +
                mat_A[245][1] * mat_B[170][1] +
                mat_A[245][2] * mat_B[178][1] +
                mat_A[245][3] * mat_B[186][1] +
                mat_A[246][0] * mat_B[194][1] +
                mat_A[246][1] * mat_B[202][1] +
                mat_A[246][2] * mat_B[210][1] +
                mat_A[246][3] * mat_B[218][1] +
                mat_A[247][0] * mat_B[226][1] +
                mat_A[247][1] * mat_B[234][1] +
                mat_A[247][2] * mat_B[242][1] +
                mat_A[247][3] * mat_B[250][1];
    mat_C[242][2] <=
                mat_A[240][0] * mat_B[2][2] +
                mat_A[240][1] * mat_B[10][2] +
                mat_A[240][2] * mat_B[18][2] +
                mat_A[240][3] * mat_B[26][2] +
                mat_A[241][0] * mat_B[34][2] +
                mat_A[241][1] * mat_B[42][2] +
                mat_A[241][2] * mat_B[50][2] +
                mat_A[241][3] * mat_B[58][2] +
                mat_A[242][0] * mat_B[66][2] +
                mat_A[242][1] * mat_B[74][2] +
                mat_A[242][2] * mat_B[82][2] +
                mat_A[242][3] * mat_B[90][2] +
                mat_A[243][0] * mat_B[98][2] +
                mat_A[243][1] * mat_B[106][2] +
                mat_A[243][2] * mat_B[114][2] +
                mat_A[243][3] * mat_B[122][2] +
                mat_A[244][0] * mat_B[130][2] +
                mat_A[244][1] * mat_B[138][2] +
                mat_A[244][2] * mat_B[146][2] +
                mat_A[244][3] * mat_B[154][2] +
                mat_A[245][0] * mat_B[162][2] +
                mat_A[245][1] * mat_B[170][2] +
                mat_A[245][2] * mat_B[178][2] +
                mat_A[245][3] * mat_B[186][2] +
                mat_A[246][0] * mat_B[194][2] +
                mat_A[246][1] * mat_B[202][2] +
                mat_A[246][2] * mat_B[210][2] +
                mat_A[246][3] * mat_B[218][2] +
                mat_A[247][0] * mat_B[226][2] +
                mat_A[247][1] * mat_B[234][2] +
                mat_A[247][2] * mat_B[242][2] +
                mat_A[247][3] * mat_B[250][2];
    mat_C[242][3] <=
                mat_A[240][0] * mat_B[2][3] +
                mat_A[240][1] * mat_B[10][3] +
                mat_A[240][2] * mat_B[18][3] +
                mat_A[240][3] * mat_B[26][3] +
                mat_A[241][0] * mat_B[34][3] +
                mat_A[241][1] * mat_B[42][3] +
                mat_A[241][2] * mat_B[50][3] +
                mat_A[241][3] * mat_B[58][3] +
                mat_A[242][0] * mat_B[66][3] +
                mat_A[242][1] * mat_B[74][3] +
                mat_A[242][2] * mat_B[82][3] +
                mat_A[242][3] * mat_B[90][3] +
                mat_A[243][0] * mat_B[98][3] +
                mat_A[243][1] * mat_B[106][3] +
                mat_A[243][2] * mat_B[114][3] +
                mat_A[243][3] * mat_B[122][3] +
                mat_A[244][0] * mat_B[130][3] +
                mat_A[244][1] * mat_B[138][3] +
                mat_A[244][2] * mat_B[146][3] +
                mat_A[244][3] * mat_B[154][3] +
                mat_A[245][0] * mat_B[162][3] +
                mat_A[245][1] * mat_B[170][3] +
                mat_A[245][2] * mat_B[178][3] +
                mat_A[245][3] * mat_B[186][3] +
                mat_A[246][0] * mat_B[194][3] +
                mat_A[246][1] * mat_B[202][3] +
                mat_A[246][2] * mat_B[210][3] +
                mat_A[246][3] * mat_B[218][3] +
                mat_A[247][0] * mat_B[226][3] +
                mat_A[247][1] * mat_B[234][3] +
                mat_A[247][2] * mat_B[242][3] +
                mat_A[247][3] * mat_B[250][3];
    mat_C[243][0] <=
                mat_A[240][0] * mat_B[3][0] +
                mat_A[240][1] * mat_B[11][0] +
                mat_A[240][2] * mat_B[19][0] +
                mat_A[240][3] * mat_B[27][0] +
                mat_A[241][0] * mat_B[35][0] +
                mat_A[241][1] * mat_B[43][0] +
                mat_A[241][2] * mat_B[51][0] +
                mat_A[241][3] * mat_B[59][0] +
                mat_A[242][0] * mat_B[67][0] +
                mat_A[242][1] * mat_B[75][0] +
                mat_A[242][2] * mat_B[83][0] +
                mat_A[242][3] * mat_B[91][0] +
                mat_A[243][0] * mat_B[99][0] +
                mat_A[243][1] * mat_B[107][0] +
                mat_A[243][2] * mat_B[115][0] +
                mat_A[243][3] * mat_B[123][0] +
                mat_A[244][0] * mat_B[131][0] +
                mat_A[244][1] * mat_B[139][0] +
                mat_A[244][2] * mat_B[147][0] +
                mat_A[244][3] * mat_B[155][0] +
                mat_A[245][0] * mat_B[163][0] +
                mat_A[245][1] * mat_B[171][0] +
                mat_A[245][2] * mat_B[179][0] +
                mat_A[245][3] * mat_B[187][0] +
                mat_A[246][0] * mat_B[195][0] +
                mat_A[246][1] * mat_B[203][0] +
                mat_A[246][2] * mat_B[211][0] +
                mat_A[246][3] * mat_B[219][0] +
                mat_A[247][0] * mat_B[227][0] +
                mat_A[247][1] * mat_B[235][0] +
                mat_A[247][2] * mat_B[243][0] +
                mat_A[247][3] * mat_B[251][0];
    mat_C[243][1] <=
                mat_A[240][0] * mat_B[3][1] +
                mat_A[240][1] * mat_B[11][1] +
                mat_A[240][2] * mat_B[19][1] +
                mat_A[240][3] * mat_B[27][1] +
                mat_A[241][0] * mat_B[35][1] +
                mat_A[241][1] * mat_B[43][1] +
                mat_A[241][2] * mat_B[51][1] +
                mat_A[241][3] * mat_B[59][1] +
                mat_A[242][0] * mat_B[67][1] +
                mat_A[242][1] * mat_B[75][1] +
                mat_A[242][2] * mat_B[83][1] +
                mat_A[242][3] * mat_B[91][1] +
                mat_A[243][0] * mat_B[99][1] +
                mat_A[243][1] * mat_B[107][1] +
                mat_A[243][2] * mat_B[115][1] +
                mat_A[243][3] * mat_B[123][1] +
                mat_A[244][0] * mat_B[131][1] +
                mat_A[244][1] * mat_B[139][1] +
                mat_A[244][2] * mat_B[147][1] +
                mat_A[244][3] * mat_B[155][1] +
                mat_A[245][0] * mat_B[163][1] +
                mat_A[245][1] * mat_B[171][1] +
                mat_A[245][2] * mat_B[179][1] +
                mat_A[245][3] * mat_B[187][1] +
                mat_A[246][0] * mat_B[195][1] +
                mat_A[246][1] * mat_B[203][1] +
                mat_A[246][2] * mat_B[211][1] +
                mat_A[246][3] * mat_B[219][1] +
                mat_A[247][0] * mat_B[227][1] +
                mat_A[247][1] * mat_B[235][1] +
                mat_A[247][2] * mat_B[243][1] +
                mat_A[247][3] * mat_B[251][1];
    mat_C[243][2] <=
                mat_A[240][0] * mat_B[3][2] +
                mat_A[240][1] * mat_B[11][2] +
                mat_A[240][2] * mat_B[19][2] +
                mat_A[240][3] * mat_B[27][2] +
                mat_A[241][0] * mat_B[35][2] +
                mat_A[241][1] * mat_B[43][2] +
                mat_A[241][2] * mat_B[51][2] +
                mat_A[241][3] * mat_B[59][2] +
                mat_A[242][0] * mat_B[67][2] +
                mat_A[242][1] * mat_B[75][2] +
                mat_A[242][2] * mat_B[83][2] +
                mat_A[242][3] * mat_B[91][2] +
                mat_A[243][0] * mat_B[99][2] +
                mat_A[243][1] * mat_B[107][2] +
                mat_A[243][2] * mat_B[115][2] +
                mat_A[243][3] * mat_B[123][2] +
                mat_A[244][0] * mat_B[131][2] +
                mat_A[244][1] * mat_B[139][2] +
                mat_A[244][2] * mat_B[147][2] +
                mat_A[244][3] * mat_B[155][2] +
                mat_A[245][0] * mat_B[163][2] +
                mat_A[245][1] * mat_B[171][2] +
                mat_A[245][2] * mat_B[179][2] +
                mat_A[245][3] * mat_B[187][2] +
                mat_A[246][0] * mat_B[195][2] +
                mat_A[246][1] * mat_B[203][2] +
                mat_A[246][2] * mat_B[211][2] +
                mat_A[246][3] * mat_B[219][2] +
                mat_A[247][0] * mat_B[227][2] +
                mat_A[247][1] * mat_B[235][2] +
                mat_A[247][2] * mat_B[243][2] +
                mat_A[247][3] * mat_B[251][2];
    mat_C[243][3] <=
                mat_A[240][0] * mat_B[3][3] +
                mat_A[240][1] * mat_B[11][3] +
                mat_A[240][2] * mat_B[19][3] +
                mat_A[240][3] * mat_B[27][3] +
                mat_A[241][0] * mat_B[35][3] +
                mat_A[241][1] * mat_B[43][3] +
                mat_A[241][2] * mat_B[51][3] +
                mat_A[241][3] * mat_B[59][3] +
                mat_A[242][0] * mat_B[67][3] +
                mat_A[242][1] * mat_B[75][3] +
                mat_A[242][2] * mat_B[83][3] +
                mat_A[242][3] * mat_B[91][3] +
                mat_A[243][0] * mat_B[99][3] +
                mat_A[243][1] * mat_B[107][3] +
                mat_A[243][2] * mat_B[115][3] +
                mat_A[243][3] * mat_B[123][3] +
                mat_A[244][0] * mat_B[131][3] +
                mat_A[244][1] * mat_B[139][3] +
                mat_A[244][2] * mat_B[147][3] +
                mat_A[244][3] * mat_B[155][3] +
                mat_A[245][0] * mat_B[163][3] +
                mat_A[245][1] * mat_B[171][3] +
                mat_A[245][2] * mat_B[179][3] +
                mat_A[245][3] * mat_B[187][3] +
                mat_A[246][0] * mat_B[195][3] +
                mat_A[246][1] * mat_B[203][3] +
                mat_A[246][2] * mat_B[211][3] +
                mat_A[246][3] * mat_B[219][3] +
                mat_A[247][0] * mat_B[227][3] +
                mat_A[247][1] * mat_B[235][3] +
                mat_A[247][2] * mat_B[243][3] +
                mat_A[247][3] * mat_B[251][3];
    mat_C[244][0] <=
                mat_A[240][0] * mat_B[4][0] +
                mat_A[240][1] * mat_B[12][0] +
                mat_A[240][2] * mat_B[20][0] +
                mat_A[240][3] * mat_B[28][0] +
                mat_A[241][0] * mat_B[36][0] +
                mat_A[241][1] * mat_B[44][0] +
                mat_A[241][2] * mat_B[52][0] +
                mat_A[241][3] * mat_B[60][0] +
                mat_A[242][0] * mat_B[68][0] +
                mat_A[242][1] * mat_B[76][0] +
                mat_A[242][2] * mat_B[84][0] +
                mat_A[242][3] * mat_B[92][0] +
                mat_A[243][0] * mat_B[100][0] +
                mat_A[243][1] * mat_B[108][0] +
                mat_A[243][2] * mat_B[116][0] +
                mat_A[243][3] * mat_B[124][0] +
                mat_A[244][0] * mat_B[132][0] +
                mat_A[244][1] * mat_B[140][0] +
                mat_A[244][2] * mat_B[148][0] +
                mat_A[244][3] * mat_B[156][0] +
                mat_A[245][0] * mat_B[164][0] +
                mat_A[245][1] * mat_B[172][0] +
                mat_A[245][2] * mat_B[180][0] +
                mat_A[245][3] * mat_B[188][0] +
                mat_A[246][0] * mat_B[196][0] +
                mat_A[246][1] * mat_B[204][0] +
                mat_A[246][2] * mat_B[212][0] +
                mat_A[246][3] * mat_B[220][0] +
                mat_A[247][0] * mat_B[228][0] +
                mat_A[247][1] * mat_B[236][0] +
                mat_A[247][2] * mat_B[244][0] +
                mat_A[247][3] * mat_B[252][0];
    mat_C[244][1] <=
                mat_A[240][0] * mat_B[4][1] +
                mat_A[240][1] * mat_B[12][1] +
                mat_A[240][2] * mat_B[20][1] +
                mat_A[240][3] * mat_B[28][1] +
                mat_A[241][0] * mat_B[36][1] +
                mat_A[241][1] * mat_B[44][1] +
                mat_A[241][2] * mat_B[52][1] +
                mat_A[241][3] * mat_B[60][1] +
                mat_A[242][0] * mat_B[68][1] +
                mat_A[242][1] * mat_B[76][1] +
                mat_A[242][2] * mat_B[84][1] +
                mat_A[242][3] * mat_B[92][1] +
                mat_A[243][0] * mat_B[100][1] +
                mat_A[243][1] * mat_B[108][1] +
                mat_A[243][2] * mat_B[116][1] +
                mat_A[243][3] * mat_B[124][1] +
                mat_A[244][0] * mat_B[132][1] +
                mat_A[244][1] * mat_B[140][1] +
                mat_A[244][2] * mat_B[148][1] +
                mat_A[244][3] * mat_B[156][1] +
                mat_A[245][0] * mat_B[164][1] +
                mat_A[245][1] * mat_B[172][1] +
                mat_A[245][2] * mat_B[180][1] +
                mat_A[245][3] * mat_B[188][1] +
                mat_A[246][0] * mat_B[196][1] +
                mat_A[246][1] * mat_B[204][1] +
                mat_A[246][2] * mat_B[212][1] +
                mat_A[246][3] * mat_B[220][1] +
                mat_A[247][0] * mat_B[228][1] +
                mat_A[247][1] * mat_B[236][1] +
                mat_A[247][2] * mat_B[244][1] +
                mat_A[247][3] * mat_B[252][1];
    mat_C[244][2] <=
                mat_A[240][0] * mat_B[4][2] +
                mat_A[240][1] * mat_B[12][2] +
                mat_A[240][2] * mat_B[20][2] +
                mat_A[240][3] * mat_B[28][2] +
                mat_A[241][0] * mat_B[36][2] +
                mat_A[241][1] * mat_B[44][2] +
                mat_A[241][2] * mat_B[52][2] +
                mat_A[241][3] * mat_B[60][2] +
                mat_A[242][0] * mat_B[68][2] +
                mat_A[242][1] * mat_B[76][2] +
                mat_A[242][2] * mat_B[84][2] +
                mat_A[242][3] * mat_B[92][2] +
                mat_A[243][0] * mat_B[100][2] +
                mat_A[243][1] * mat_B[108][2] +
                mat_A[243][2] * mat_B[116][2] +
                mat_A[243][3] * mat_B[124][2] +
                mat_A[244][0] * mat_B[132][2] +
                mat_A[244][1] * mat_B[140][2] +
                mat_A[244][2] * mat_B[148][2] +
                mat_A[244][3] * mat_B[156][2] +
                mat_A[245][0] * mat_B[164][2] +
                mat_A[245][1] * mat_B[172][2] +
                mat_A[245][2] * mat_B[180][2] +
                mat_A[245][3] * mat_B[188][2] +
                mat_A[246][0] * mat_B[196][2] +
                mat_A[246][1] * mat_B[204][2] +
                mat_A[246][2] * mat_B[212][2] +
                mat_A[246][3] * mat_B[220][2] +
                mat_A[247][0] * mat_B[228][2] +
                mat_A[247][1] * mat_B[236][2] +
                mat_A[247][2] * mat_B[244][2] +
                mat_A[247][3] * mat_B[252][2];
    mat_C[244][3] <=
                mat_A[240][0] * mat_B[4][3] +
                mat_A[240][1] * mat_B[12][3] +
                mat_A[240][2] * mat_B[20][3] +
                mat_A[240][3] * mat_B[28][3] +
                mat_A[241][0] * mat_B[36][3] +
                mat_A[241][1] * mat_B[44][3] +
                mat_A[241][2] * mat_B[52][3] +
                mat_A[241][3] * mat_B[60][3] +
                mat_A[242][0] * mat_B[68][3] +
                mat_A[242][1] * mat_B[76][3] +
                mat_A[242][2] * mat_B[84][3] +
                mat_A[242][3] * mat_B[92][3] +
                mat_A[243][0] * mat_B[100][3] +
                mat_A[243][1] * mat_B[108][3] +
                mat_A[243][2] * mat_B[116][3] +
                mat_A[243][3] * mat_B[124][3] +
                mat_A[244][0] * mat_B[132][3] +
                mat_A[244][1] * mat_B[140][3] +
                mat_A[244][2] * mat_B[148][3] +
                mat_A[244][3] * mat_B[156][3] +
                mat_A[245][0] * mat_B[164][3] +
                mat_A[245][1] * mat_B[172][3] +
                mat_A[245][2] * mat_B[180][3] +
                mat_A[245][3] * mat_B[188][3] +
                mat_A[246][0] * mat_B[196][3] +
                mat_A[246][1] * mat_B[204][3] +
                mat_A[246][2] * mat_B[212][3] +
                mat_A[246][3] * mat_B[220][3] +
                mat_A[247][0] * mat_B[228][3] +
                mat_A[247][1] * mat_B[236][3] +
                mat_A[247][2] * mat_B[244][3] +
                mat_A[247][3] * mat_B[252][3];
    mat_C[245][0] <=
                mat_A[240][0] * mat_B[5][0] +
                mat_A[240][1] * mat_B[13][0] +
                mat_A[240][2] * mat_B[21][0] +
                mat_A[240][3] * mat_B[29][0] +
                mat_A[241][0] * mat_B[37][0] +
                mat_A[241][1] * mat_B[45][0] +
                mat_A[241][2] * mat_B[53][0] +
                mat_A[241][3] * mat_B[61][0] +
                mat_A[242][0] * mat_B[69][0] +
                mat_A[242][1] * mat_B[77][0] +
                mat_A[242][2] * mat_B[85][0] +
                mat_A[242][3] * mat_B[93][0] +
                mat_A[243][0] * mat_B[101][0] +
                mat_A[243][1] * mat_B[109][0] +
                mat_A[243][2] * mat_B[117][0] +
                mat_A[243][3] * mat_B[125][0] +
                mat_A[244][0] * mat_B[133][0] +
                mat_A[244][1] * mat_B[141][0] +
                mat_A[244][2] * mat_B[149][0] +
                mat_A[244][3] * mat_B[157][0] +
                mat_A[245][0] * mat_B[165][0] +
                mat_A[245][1] * mat_B[173][0] +
                mat_A[245][2] * mat_B[181][0] +
                mat_A[245][3] * mat_B[189][0] +
                mat_A[246][0] * mat_B[197][0] +
                mat_A[246][1] * mat_B[205][0] +
                mat_A[246][2] * mat_B[213][0] +
                mat_A[246][3] * mat_B[221][0] +
                mat_A[247][0] * mat_B[229][0] +
                mat_A[247][1] * mat_B[237][0] +
                mat_A[247][2] * mat_B[245][0] +
                mat_A[247][3] * mat_B[253][0];
    mat_C[245][1] <=
                mat_A[240][0] * mat_B[5][1] +
                mat_A[240][1] * mat_B[13][1] +
                mat_A[240][2] * mat_B[21][1] +
                mat_A[240][3] * mat_B[29][1] +
                mat_A[241][0] * mat_B[37][1] +
                mat_A[241][1] * mat_B[45][1] +
                mat_A[241][2] * mat_B[53][1] +
                mat_A[241][3] * mat_B[61][1] +
                mat_A[242][0] * mat_B[69][1] +
                mat_A[242][1] * mat_B[77][1] +
                mat_A[242][2] * mat_B[85][1] +
                mat_A[242][3] * mat_B[93][1] +
                mat_A[243][0] * mat_B[101][1] +
                mat_A[243][1] * mat_B[109][1] +
                mat_A[243][2] * mat_B[117][1] +
                mat_A[243][3] * mat_B[125][1] +
                mat_A[244][0] * mat_B[133][1] +
                mat_A[244][1] * mat_B[141][1] +
                mat_A[244][2] * mat_B[149][1] +
                mat_A[244][3] * mat_B[157][1] +
                mat_A[245][0] * mat_B[165][1] +
                mat_A[245][1] * mat_B[173][1] +
                mat_A[245][2] * mat_B[181][1] +
                mat_A[245][3] * mat_B[189][1] +
                mat_A[246][0] * mat_B[197][1] +
                mat_A[246][1] * mat_B[205][1] +
                mat_A[246][2] * mat_B[213][1] +
                mat_A[246][3] * mat_B[221][1] +
                mat_A[247][0] * mat_B[229][1] +
                mat_A[247][1] * mat_B[237][1] +
                mat_A[247][2] * mat_B[245][1] +
                mat_A[247][3] * mat_B[253][1];
    mat_C[245][2] <=
                mat_A[240][0] * mat_B[5][2] +
                mat_A[240][1] * mat_B[13][2] +
                mat_A[240][2] * mat_B[21][2] +
                mat_A[240][3] * mat_B[29][2] +
                mat_A[241][0] * mat_B[37][2] +
                mat_A[241][1] * mat_B[45][2] +
                mat_A[241][2] * mat_B[53][2] +
                mat_A[241][3] * mat_B[61][2] +
                mat_A[242][0] * mat_B[69][2] +
                mat_A[242][1] * mat_B[77][2] +
                mat_A[242][2] * mat_B[85][2] +
                mat_A[242][3] * mat_B[93][2] +
                mat_A[243][0] * mat_B[101][2] +
                mat_A[243][1] * mat_B[109][2] +
                mat_A[243][2] * mat_B[117][2] +
                mat_A[243][3] * mat_B[125][2] +
                mat_A[244][0] * mat_B[133][2] +
                mat_A[244][1] * mat_B[141][2] +
                mat_A[244][2] * mat_B[149][2] +
                mat_A[244][3] * mat_B[157][2] +
                mat_A[245][0] * mat_B[165][2] +
                mat_A[245][1] * mat_B[173][2] +
                mat_A[245][2] * mat_B[181][2] +
                mat_A[245][3] * mat_B[189][2] +
                mat_A[246][0] * mat_B[197][2] +
                mat_A[246][1] * mat_B[205][2] +
                mat_A[246][2] * mat_B[213][2] +
                mat_A[246][3] * mat_B[221][2] +
                mat_A[247][0] * mat_B[229][2] +
                mat_A[247][1] * mat_B[237][2] +
                mat_A[247][2] * mat_B[245][2] +
                mat_A[247][3] * mat_B[253][2];
    mat_C[245][3] <=
                mat_A[240][0] * mat_B[5][3] +
                mat_A[240][1] * mat_B[13][3] +
                mat_A[240][2] * mat_B[21][3] +
                mat_A[240][3] * mat_B[29][3] +
                mat_A[241][0] * mat_B[37][3] +
                mat_A[241][1] * mat_B[45][3] +
                mat_A[241][2] * mat_B[53][3] +
                mat_A[241][3] * mat_B[61][3] +
                mat_A[242][0] * mat_B[69][3] +
                mat_A[242][1] * mat_B[77][3] +
                mat_A[242][2] * mat_B[85][3] +
                mat_A[242][3] * mat_B[93][3] +
                mat_A[243][0] * mat_B[101][3] +
                mat_A[243][1] * mat_B[109][3] +
                mat_A[243][2] * mat_B[117][3] +
                mat_A[243][3] * mat_B[125][3] +
                mat_A[244][0] * mat_B[133][3] +
                mat_A[244][1] * mat_B[141][3] +
                mat_A[244][2] * mat_B[149][3] +
                mat_A[244][3] * mat_B[157][3] +
                mat_A[245][0] * mat_B[165][3] +
                mat_A[245][1] * mat_B[173][3] +
                mat_A[245][2] * mat_B[181][3] +
                mat_A[245][3] * mat_B[189][3] +
                mat_A[246][0] * mat_B[197][3] +
                mat_A[246][1] * mat_B[205][3] +
                mat_A[246][2] * mat_B[213][3] +
                mat_A[246][3] * mat_B[221][3] +
                mat_A[247][0] * mat_B[229][3] +
                mat_A[247][1] * mat_B[237][3] +
                mat_A[247][2] * mat_B[245][3] +
                mat_A[247][3] * mat_B[253][3];
    mat_C[246][0] <=
                mat_A[240][0] * mat_B[6][0] +
                mat_A[240][1] * mat_B[14][0] +
                mat_A[240][2] * mat_B[22][0] +
                mat_A[240][3] * mat_B[30][0] +
                mat_A[241][0] * mat_B[38][0] +
                mat_A[241][1] * mat_B[46][0] +
                mat_A[241][2] * mat_B[54][0] +
                mat_A[241][3] * mat_B[62][0] +
                mat_A[242][0] * mat_B[70][0] +
                mat_A[242][1] * mat_B[78][0] +
                mat_A[242][2] * mat_B[86][0] +
                mat_A[242][3] * mat_B[94][0] +
                mat_A[243][0] * mat_B[102][0] +
                mat_A[243][1] * mat_B[110][0] +
                mat_A[243][2] * mat_B[118][0] +
                mat_A[243][3] * mat_B[126][0] +
                mat_A[244][0] * mat_B[134][0] +
                mat_A[244][1] * mat_B[142][0] +
                mat_A[244][2] * mat_B[150][0] +
                mat_A[244][3] * mat_B[158][0] +
                mat_A[245][0] * mat_B[166][0] +
                mat_A[245][1] * mat_B[174][0] +
                mat_A[245][2] * mat_B[182][0] +
                mat_A[245][3] * mat_B[190][0] +
                mat_A[246][0] * mat_B[198][0] +
                mat_A[246][1] * mat_B[206][0] +
                mat_A[246][2] * mat_B[214][0] +
                mat_A[246][3] * mat_B[222][0] +
                mat_A[247][0] * mat_B[230][0] +
                mat_A[247][1] * mat_B[238][0] +
                mat_A[247][2] * mat_B[246][0] +
                mat_A[247][3] * mat_B[254][0];
    mat_C[246][1] <=
                mat_A[240][0] * mat_B[6][1] +
                mat_A[240][1] * mat_B[14][1] +
                mat_A[240][2] * mat_B[22][1] +
                mat_A[240][3] * mat_B[30][1] +
                mat_A[241][0] * mat_B[38][1] +
                mat_A[241][1] * mat_B[46][1] +
                mat_A[241][2] * mat_B[54][1] +
                mat_A[241][3] * mat_B[62][1] +
                mat_A[242][0] * mat_B[70][1] +
                mat_A[242][1] * mat_B[78][1] +
                mat_A[242][2] * mat_B[86][1] +
                mat_A[242][3] * mat_B[94][1] +
                mat_A[243][0] * mat_B[102][1] +
                mat_A[243][1] * mat_B[110][1] +
                mat_A[243][2] * mat_B[118][1] +
                mat_A[243][3] * mat_B[126][1] +
                mat_A[244][0] * mat_B[134][1] +
                mat_A[244][1] * mat_B[142][1] +
                mat_A[244][2] * mat_B[150][1] +
                mat_A[244][3] * mat_B[158][1] +
                mat_A[245][0] * mat_B[166][1] +
                mat_A[245][1] * mat_B[174][1] +
                mat_A[245][2] * mat_B[182][1] +
                mat_A[245][3] * mat_B[190][1] +
                mat_A[246][0] * mat_B[198][1] +
                mat_A[246][1] * mat_B[206][1] +
                mat_A[246][2] * mat_B[214][1] +
                mat_A[246][3] * mat_B[222][1] +
                mat_A[247][0] * mat_B[230][1] +
                mat_A[247][1] * mat_B[238][1] +
                mat_A[247][2] * mat_B[246][1] +
                mat_A[247][3] * mat_B[254][1];
    mat_C[246][2] <=
                mat_A[240][0] * mat_B[6][2] +
                mat_A[240][1] * mat_B[14][2] +
                mat_A[240][2] * mat_B[22][2] +
                mat_A[240][3] * mat_B[30][2] +
                mat_A[241][0] * mat_B[38][2] +
                mat_A[241][1] * mat_B[46][2] +
                mat_A[241][2] * mat_B[54][2] +
                mat_A[241][3] * mat_B[62][2] +
                mat_A[242][0] * mat_B[70][2] +
                mat_A[242][1] * mat_B[78][2] +
                mat_A[242][2] * mat_B[86][2] +
                mat_A[242][3] * mat_B[94][2] +
                mat_A[243][0] * mat_B[102][2] +
                mat_A[243][1] * mat_B[110][2] +
                mat_A[243][2] * mat_B[118][2] +
                mat_A[243][3] * mat_B[126][2] +
                mat_A[244][0] * mat_B[134][2] +
                mat_A[244][1] * mat_B[142][2] +
                mat_A[244][2] * mat_B[150][2] +
                mat_A[244][3] * mat_B[158][2] +
                mat_A[245][0] * mat_B[166][2] +
                mat_A[245][1] * mat_B[174][2] +
                mat_A[245][2] * mat_B[182][2] +
                mat_A[245][3] * mat_B[190][2] +
                mat_A[246][0] * mat_B[198][2] +
                mat_A[246][1] * mat_B[206][2] +
                mat_A[246][2] * mat_B[214][2] +
                mat_A[246][3] * mat_B[222][2] +
                mat_A[247][0] * mat_B[230][2] +
                mat_A[247][1] * mat_B[238][2] +
                mat_A[247][2] * mat_B[246][2] +
                mat_A[247][3] * mat_B[254][2];
    mat_C[246][3] <=
                mat_A[240][0] * mat_B[6][3] +
                mat_A[240][1] * mat_B[14][3] +
                mat_A[240][2] * mat_B[22][3] +
                mat_A[240][3] * mat_B[30][3] +
                mat_A[241][0] * mat_B[38][3] +
                mat_A[241][1] * mat_B[46][3] +
                mat_A[241][2] * mat_B[54][3] +
                mat_A[241][3] * mat_B[62][3] +
                mat_A[242][0] * mat_B[70][3] +
                mat_A[242][1] * mat_B[78][3] +
                mat_A[242][2] * mat_B[86][3] +
                mat_A[242][3] * mat_B[94][3] +
                mat_A[243][0] * mat_B[102][3] +
                mat_A[243][1] * mat_B[110][3] +
                mat_A[243][2] * mat_B[118][3] +
                mat_A[243][3] * mat_B[126][3] +
                mat_A[244][0] * mat_B[134][3] +
                mat_A[244][1] * mat_B[142][3] +
                mat_A[244][2] * mat_B[150][3] +
                mat_A[244][3] * mat_B[158][3] +
                mat_A[245][0] * mat_B[166][3] +
                mat_A[245][1] * mat_B[174][3] +
                mat_A[245][2] * mat_B[182][3] +
                mat_A[245][3] * mat_B[190][3] +
                mat_A[246][0] * mat_B[198][3] +
                mat_A[246][1] * mat_B[206][3] +
                mat_A[246][2] * mat_B[214][3] +
                mat_A[246][3] * mat_B[222][3] +
                mat_A[247][0] * mat_B[230][3] +
                mat_A[247][1] * mat_B[238][3] +
                mat_A[247][2] * mat_B[246][3] +
                mat_A[247][3] * mat_B[254][3];
    mat_C[247][0] <=
                mat_A[240][0] * mat_B[7][0] +
                mat_A[240][1] * mat_B[15][0] +
                mat_A[240][2] * mat_B[23][0] +
                mat_A[240][3] * mat_B[31][0] +
                mat_A[241][0] * mat_B[39][0] +
                mat_A[241][1] * mat_B[47][0] +
                mat_A[241][2] * mat_B[55][0] +
                mat_A[241][3] * mat_B[63][0] +
                mat_A[242][0] * mat_B[71][0] +
                mat_A[242][1] * mat_B[79][0] +
                mat_A[242][2] * mat_B[87][0] +
                mat_A[242][3] * mat_B[95][0] +
                mat_A[243][0] * mat_B[103][0] +
                mat_A[243][1] * mat_B[111][0] +
                mat_A[243][2] * mat_B[119][0] +
                mat_A[243][3] * mat_B[127][0] +
                mat_A[244][0] * mat_B[135][0] +
                mat_A[244][1] * mat_B[143][0] +
                mat_A[244][2] * mat_B[151][0] +
                mat_A[244][3] * mat_B[159][0] +
                mat_A[245][0] * mat_B[167][0] +
                mat_A[245][1] * mat_B[175][0] +
                mat_A[245][2] * mat_B[183][0] +
                mat_A[245][3] * mat_B[191][0] +
                mat_A[246][0] * mat_B[199][0] +
                mat_A[246][1] * mat_B[207][0] +
                mat_A[246][2] * mat_B[215][0] +
                mat_A[246][3] * mat_B[223][0] +
                mat_A[247][0] * mat_B[231][0] +
                mat_A[247][1] * mat_B[239][0] +
                mat_A[247][2] * mat_B[247][0] +
                mat_A[247][3] * mat_B[255][0];
    mat_C[247][1] <=
                mat_A[240][0] * mat_B[7][1] +
                mat_A[240][1] * mat_B[15][1] +
                mat_A[240][2] * mat_B[23][1] +
                mat_A[240][3] * mat_B[31][1] +
                mat_A[241][0] * mat_B[39][1] +
                mat_A[241][1] * mat_B[47][1] +
                mat_A[241][2] * mat_B[55][1] +
                mat_A[241][3] * mat_B[63][1] +
                mat_A[242][0] * mat_B[71][1] +
                mat_A[242][1] * mat_B[79][1] +
                mat_A[242][2] * mat_B[87][1] +
                mat_A[242][3] * mat_B[95][1] +
                mat_A[243][0] * mat_B[103][1] +
                mat_A[243][1] * mat_B[111][1] +
                mat_A[243][2] * mat_B[119][1] +
                mat_A[243][3] * mat_B[127][1] +
                mat_A[244][0] * mat_B[135][1] +
                mat_A[244][1] * mat_B[143][1] +
                mat_A[244][2] * mat_B[151][1] +
                mat_A[244][3] * mat_B[159][1] +
                mat_A[245][0] * mat_B[167][1] +
                mat_A[245][1] * mat_B[175][1] +
                mat_A[245][2] * mat_B[183][1] +
                mat_A[245][3] * mat_B[191][1] +
                mat_A[246][0] * mat_B[199][1] +
                mat_A[246][1] * mat_B[207][1] +
                mat_A[246][2] * mat_B[215][1] +
                mat_A[246][3] * mat_B[223][1] +
                mat_A[247][0] * mat_B[231][1] +
                mat_A[247][1] * mat_B[239][1] +
                mat_A[247][2] * mat_B[247][1] +
                mat_A[247][3] * mat_B[255][1];
    mat_C[247][2] <=
                mat_A[240][0] * mat_B[7][2] +
                mat_A[240][1] * mat_B[15][2] +
                mat_A[240][2] * mat_B[23][2] +
                mat_A[240][3] * mat_B[31][2] +
                mat_A[241][0] * mat_B[39][2] +
                mat_A[241][1] * mat_B[47][2] +
                mat_A[241][2] * mat_B[55][2] +
                mat_A[241][3] * mat_B[63][2] +
                mat_A[242][0] * mat_B[71][2] +
                mat_A[242][1] * mat_B[79][2] +
                mat_A[242][2] * mat_B[87][2] +
                mat_A[242][3] * mat_B[95][2] +
                mat_A[243][0] * mat_B[103][2] +
                mat_A[243][1] * mat_B[111][2] +
                mat_A[243][2] * mat_B[119][2] +
                mat_A[243][3] * mat_B[127][2] +
                mat_A[244][0] * mat_B[135][2] +
                mat_A[244][1] * mat_B[143][2] +
                mat_A[244][2] * mat_B[151][2] +
                mat_A[244][3] * mat_B[159][2] +
                mat_A[245][0] * mat_B[167][2] +
                mat_A[245][1] * mat_B[175][2] +
                mat_A[245][2] * mat_B[183][2] +
                mat_A[245][3] * mat_B[191][2] +
                mat_A[246][0] * mat_B[199][2] +
                mat_A[246][1] * mat_B[207][2] +
                mat_A[246][2] * mat_B[215][2] +
                mat_A[246][3] * mat_B[223][2] +
                mat_A[247][0] * mat_B[231][2] +
                mat_A[247][1] * mat_B[239][2] +
                mat_A[247][2] * mat_B[247][2] +
                mat_A[247][3] * mat_B[255][2];
    mat_C[247][3] <=
                mat_A[240][0] * mat_B[7][3] +
                mat_A[240][1] * mat_B[15][3] +
                mat_A[240][2] * mat_B[23][3] +
                mat_A[240][3] * mat_B[31][3] +
                mat_A[241][0] * mat_B[39][3] +
                mat_A[241][1] * mat_B[47][3] +
                mat_A[241][2] * mat_B[55][3] +
                mat_A[241][3] * mat_B[63][3] +
                mat_A[242][0] * mat_B[71][3] +
                mat_A[242][1] * mat_B[79][3] +
                mat_A[242][2] * mat_B[87][3] +
                mat_A[242][3] * mat_B[95][3] +
                mat_A[243][0] * mat_B[103][3] +
                mat_A[243][1] * mat_B[111][3] +
                mat_A[243][2] * mat_B[119][3] +
                mat_A[243][3] * mat_B[127][3] +
                mat_A[244][0] * mat_B[135][3] +
                mat_A[244][1] * mat_B[143][3] +
                mat_A[244][2] * mat_B[151][3] +
                mat_A[244][3] * mat_B[159][3] +
                mat_A[245][0] * mat_B[167][3] +
                mat_A[245][1] * mat_B[175][3] +
                mat_A[245][2] * mat_B[183][3] +
                mat_A[245][3] * mat_B[191][3] +
                mat_A[246][0] * mat_B[199][3] +
                mat_A[246][1] * mat_B[207][3] +
                mat_A[246][2] * mat_B[215][3] +
                mat_A[246][3] * mat_B[223][3] +
                mat_A[247][0] * mat_B[231][3] +
                mat_A[247][1] * mat_B[239][3] +
                mat_A[247][2] * mat_B[247][3] +
                mat_A[247][3] * mat_B[255][3];
    mat_C[248][0] <=
                mat_A[248][0] * mat_B[0][0] +
                mat_A[248][1] * mat_B[8][0] +
                mat_A[248][2] * mat_B[16][0] +
                mat_A[248][3] * mat_B[24][0] +
                mat_A[249][0] * mat_B[32][0] +
                mat_A[249][1] * mat_B[40][0] +
                mat_A[249][2] * mat_B[48][0] +
                mat_A[249][3] * mat_B[56][0] +
                mat_A[250][0] * mat_B[64][0] +
                mat_A[250][1] * mat_B[72][0] +
                mat_A[250][2] * mat_B[80][0] +
                mat_A[250][3] * mat_B[88][0] +
                mat_A[251][0] * mat_B[96][0] +
                mat_A[251][1] * mat_B[104][0] +
                mat_A[251][2] * mat_B[112][0] +
                mat_A[251][3] * mat_B[120][0] +
                mat_A[252][0] * mat_B[128][0] +
                mat_A[252][1] * mat_B[136][0] +
                mat_A[252][2] * mat_B[144][0] +
                mat_A[252][3] * mat_B[152][0] +
                mat_A[253][0] * mat_B[160][0] +
                mat_A[253][1] * mat_B[168][0] +
                mat_A[253][2] * mat_B[176][0] +
                mat_A[253][3] * mat_B[184][0] +
                mat_A[254][0] * mat_B[192][0] +
                mat_A[254][1] * mat_B[200][0] +
                mat_A[254][2] * mat_B[208][0] +
                mat_A[254][3] * mat_B[216][0] +
                mat_A[255][0] * mat_B[224][0] +
                mat_A[255][1] * mat_B[232][0] +
                mat_A[255][2] * mat_B[240][0] +
                mat_A[255][3] * mat_B[248][0];
    mat_C[248][1] <=
                mat_A[248][0] * mat_B[0][1] +
                mat_A[248][1] * mat_B[8][1] +
                mat_A[248][2] * mat_B[16][1] +
                mat_A[248][3] * mat_B[24][1] +
                mat_A[249][0] * mat_B[32][1] +
                mat_A[249][1] * mat_B[40][1] +
                mat_A[249][2] * mat_B[48][1] +
                mat_A[249][3] * mat_B[56][1] +
                mat_A[250][0] * mat_B[64][1] +
                mat_A[250][1] * mat_B[72][1] +
                mat_A[250][2] * mat_B[80][1] +
                mat_A[250][3] * mat_B[88][1] +
                mat_A[251][0] * mat_B[96][1] +
                mat_A[251][1] * mat_B[104][1] +
                mat_A[251][2] * mat_B[112][1] +
                mat_A[251][3] * mat_B[120][1] +
                mat_A[252][0] * mat_B[128][1] +
                mat_A[252][1] * mat_B[136][1] +
                mat_A[252][2] * mat_B[144][1] +
                mat_A[252][3] * mat_B[152][1] +
                mat_A[253][0] * mat_B[160][1] +
                mat_A[253][1] * mat_B[168][1] +
                mat_A[253][2] * mat_B[176][1] +
                mat_A[253][3] * mat_B[184][1] +
                mat_A[254][0] * mat_B[192][1] +
                mat_A[254][1] * mat_B[200][1] +
                mat_A[254][2] * mat_B[208][1] +
                mat_A[254][3] * mat_B[216][1] +
                mat_A[255][0] * mat_B[224][1] +
                mat_A[255][1] * mat_B[232][1] +
                mat_A[255][2] * mat_B[240][1] +
                mat_A[255][3] * mat_B[248][1];
    mat_C[248][2] <=
                mat_A[248][0] * mat_B[0][2] +
                mat_A[248][1] * mat_B[8][2] +
                mat_A[248][2] * mat_B[16][2] +
                mat_A[248][3] * mat_B[24][2] +
                mat_A[249][0] * mat_B[32][2] +
                mat_A[249][1] * mat_B[40][2] +
                mat_A[249][2] * mat_B[48][2] +
                mat_A[249][3] * mat_B[56][2] +
                mat_A[250][0] * mat_B[64][2] +
                mat_A[250][1] * mat_B[72][2] +
                mat_A[250][2] * mat_B[80][2] +
                mat_A[250][3] * mat_B[88][2] +
                mat_A[251][0] * mat_B[96][2] +
                mat_A[251][1] * mat_B[104][2] +
                mat_A[251][2] * mat_B[112][2] +
                mat_A[251][3] * mat_B[120][2] +
                mat_A[252][0] * mat_B[128][2] +
                mat_A[252][1] * mat_B[136][2] +
                mat_A[252][2] * mat_B[144][2] +
                mat_A[252][3] * mat_B[152][2] +
                mat_A[253][0] * mat_B[160][2] +
                mat_A[253][1] * mat_B[168][2] +
                mat_A[253][2] * mat_B[176][2] +
                mat_A[253][3] * mat_B[184][2] +
                mat_A[254][0] * mat_B[192][2] +
                mat_A[254][1] * mat_B[200][2] +
                mat_A[254][2] * mat_B[208][2] +
                mat_A[254][3] * mat_B[216][2] +
                mat_A[255][0] * mat_B[224][2] +
                mat_A[255][1] * mat_B[232][2] +
                mat_A[255][2] * mat_B[240][2] +
                mat_A[255][3] * mat_B[248][2];
    mat_C[248][3] <=
                mat_A[248][0] * mat_B[0][3] +
                mat_A[248][1] * mat_B[8][3] +
                mat_A[248][2] * mat_B[16][3] +
                mat_A[248][3] * mat_B[24][3] +
                mat_A[249][0] * mat_B[32][3] +
                mat_A[249][1] * mat_B[40][3] +
                mat_A[249][2] * mat_B[48][3] +
                mat_A[249][3] * mat_B[56][3] +
                mat_A[250][0] * mat_B[64][3] +
                mat_A[250][1] * mat_B[72][3] +
                mat_A[250][2] * mat_B[80][3] +
                mat_A[250][3] * mat_B[88][3] +
                mat_A[251][0] * mat_B[96][3] +
                mat_A[251][1] * mat_B[104][3] +
                mat_A[251][2] * mat_B[112][3] +
                mat_A[251][3] * mat_B[120][3] +
                mat_A[252][0] * mat_B[128][3] +
                mat_A[252][1] * mat_B[136][3] +
                mat_A[252][2] * mat_B[144][3] +
                mat_A[252][3] * mat_B[152][3] +
                mat_A[253][0] * mat_B[160][3] +
                mat_A[253][1] * mat_B[168][3] +
                mat_A[253][2] * mat_B[176][3] +
                mat_A[253][3] * mat_B[184][3] +
                mat_A[254][0] * mat_B[192][3] +
                mat_A[254][1] * mat_B[200][3] +
                mat_A[254][2] * mat_B[208][3] +
                mat_A[254][3] * mat_B[216][3] +
                mat_A[255][0] * mat_B[224][3] +
                mat_A[255][1] * mat_B[232][3] +
                mat_A[255][2] * mat_B[240][3] +
                mat_A[255][3] * mat_B[248][3];
    mat_C[249][0] <=
                mat_A[248][0] * mat_B[1][0] +
                mat_A[248][1] * mat_B[9][0] +
                mat_A[248][2] * mat_B[17][0] +
                mat_A[248][3] * mat_B[25][0] +
                mat_A[249][0] * mat_B[33][0] +
                mat_A[249][1] * mat_B[41][0] +
                mat_A[249][2] * mat_B[49][0] +
                mat_A[249][3] * mat_B[57][0] +
                mat_A[250][0] * mat_B[65][0] +
                mat_A[250][1] * mat_B[73][0] +
                mat_A[250][2] * mat_B[81][0] +
                mat_A[250][3] * mat_B[89][0] +
                mat_A[251][0] * mat_B[97][0] +
                mat_A[251][1] * mat_B[105][0] +
                mat_A[251][2] * mat_B[113][0] +
                mat_A[251][3] * mat_B[121][0] +
                mat_A[252][0] * mat_B[129][0] +
                mat_A[252][1] * mat_B[137][0] +
                mat_A[252][2] * mat_B[145][0] +
                mat_A[252][3] * mat_B[153][0] +
                mat_A[253][0] * mat_B[161][0] +
                mat_A[253][1] * mat_B[169][0] +
                mat_A[253][2] * mat_B[177][0] +
                mat_A[253][3] * mat_B[185][0] +
                mat_A[254][0] * mat_B[193][0] +
                mat_A[254][1] * mat_B[201][0] +
                mat_A[254][2] * mat_B[209][0] +
                mat_A[254][3] * mat_B[217][0] +
                mat_A[255][0] * mat_B[225][0] +
                mat_A[255][1] * mat_B[233][0] +
                mat_A[255][2] * mat_B[241][0] +
                mat_A[255][3] * mat_B[249][0];
    mat_C[249][1] <=
                mat_A[248][0] * mat_B[1][1] +
                mat_A[248][1] * mat_B[9][1] +
                mat_A[248][2] * mat_B[17][1] +
                mat_A[248][3] * mat_B[25][1] +
                mat_A[249][0] * mat_B[33][1] +
                mat_A[249][1] * mat_B[41][1] +
                mat_A[249][2] * mat_B[49][1] +
                mat_A[249][3] * mat_B[57][1] +
                mat_A[250][0] * mat_B[65][1] +
                mat_A[250][1] * mat_B[73][1] +
                mat_A[250][2] * mat_B[81][1] +
                mat_A[250][3] * mat_B[89][1] +
                mat_A[251][0] * mat_B[97][1] +
                mat_A[251][1] * mat_B[105][1] +
                mat_A[251][2] * mat_B[113][1] +
                mat_A[251][3] * mat_B[121][1] +
                mat_A[252][0] * mat_B[129][1] +
                mat_A[252][1] * mat_B[137][1] +
                mat_A[252][2] * mat_B[145][1] +
                mat_A[252][3] * mat_B[153][1] +
                mat_A[253][0] * mat_B[161][1] +
                mat_A[253][1] * mat_B[169][1] +
                mat_A[253][2] * mat_B[177][1] +
                mat_A[253][3] * mat_B[185][1] +
                mat_A[254][0] * mat_B[193][1] +
                mat_A[254][1] * mat_B[201][1] +
                mat_A[254][2] * mat_B[209][1] +
                mat_A[254][3] * mat_B[217][1] +
                mat_A[255][0] * mat_B[225][1] +
                mat_A[255][1] * mat_B[233][1] +
                mat_A[255][2] * mat_B[241][1] +
                mat_A[255][3] * mat_B[249][1];
    mat_C[249][2] <=
                mat_A[248][0] * mat_B[1][2] +
                mat_A[248][1] * mat_B[9][2] +
                mat_A[248][2] * mat_B[17][2] +
                mat_A[248][3] * mat_B[25][2] +
                mat_A[249][0] * mat_B[33][2] +
                mat_A[249][1] * mat_B[41][2] +
                mat_A[249][2] * mat_B[49][2] +
                mat_A[249][3] * mat_B[57][2] +
                mat_A[250][0] * mat_B[65][2] +
                mat_A[250][1] * mat_B[73][2] +
                mat_A[250][2] * mat_B[81][2] +
                mat_A[250][3] * mat_B[89][2] +
                mat_A[251][0] * mat_B[97][2] +
                mat_A[251][1] * mat_B[105][2] +
                mat_A[251][2] * mat_B[113][2] +
                mat_A[251][3] * mat_B[121][2] +
                mat_A[252][0] * mat_B[129][2] +
                mat_A[252][1] * mat_B[137][2] +
                mat_A[252][2] * mat_B[145][2] +
                mat_A[252][3] * mat_B[153][2] +
                mat_A[253][0] * mat_B[161][2] +
                mat_A[253][1] * mat_B[169][2] +
                mat_A[253][2] * mat_B[177][2] +
                mat_A[253][3] * mat_B[185][2] +
                mat_A[254][0] * mat_B[193][2] +
                mat_A[254][1] * mat_B[201][2] +
                mat_A[254][2] * mat_B[209][2] +
                mat_A[254][3] * mat_B[217][2] +
                mat_A[255][0] * mat_B[225][2] +
                mat_A[255][1] * mat_B[233][2] +
                mat_A[255][2] * mat_B[241][2] +
                mat_A[255][3] * mat_B[249][2];
    mat_C[249][3] <=
                mat_A[248][0] * mat_B[1][3] +
                mat_A[248][1] * mat_B[9][3] +
                mat_A[248][2] * mat_B[17][3] +
                mat_A[248][3] * mat_B[25][3] +
                mat_A[249][0] * mat_B[33][3] +
                mat_A[249][1] * mat_B[41][3] +
                mat_A[249][2] * mat_B[49][3] +
                mat_A[249][3] * mat_B[57][3] +
                mat_A[250][0] * mat_B[65][3] +
                mat_A[250][1] * mat_B[73][3] +
                mat_A[250][2] * mat_B[81][3] +
                mat_A[250][3] * mat_B[89][3] +
                mat_A[251][0] * mat_B[97][3] +
                mat_A[251][1] * mat_B[105][3] +
                mat_A[251][2] * mat_B[113][3] +
                mat_A[251][3] * mat_B[121][3] +
                mat_A[252][0] * mat_B[129][3] +
                mat_A[252][1] * mat_B[137][3] +
                mat_A[252][2] * mat_B[145][3] +
                mat_A[252][3] * mat_B[153][3] +
                mat_A[253][0] * mat_B[161][3] +
                mat_A[253][1] * mat_B[169][3] +
                mat_A[253][2] * mat_B[177][3] +
                mat_A[253][3] * mat_B[185][3] +
                mat_A[254][0] * mat_B[193][3] +
                mat_A[254][1] * mat_B[201][3] +
                mat_A[254][2] * mat_B[209][3] +
                mat_A[254][3] * mat_B[217][3] +
                mat_A[255][0] * mat_B[225][3] +
                mat_A[255][1] * mat_B[233][3] +
                mat_A[255][2] * mat_B[241][3] +
                mat_A[255][3] * mat_B[249][3];
    mat_C[250][0] <=
                mat_A[248][0] * mat_B[2][0] +
                mat_A[248][1] * mat_B[10][0] +
                mat_A[248][2] * mat_B[18][0] +
                mat_A[248][3] * mat_B[26][0] +
                mat_A[249][0] * mat_B[34][0] +
                mat_A[249][1] * mat_B[42][0] +
                mat_A[249][2] * mat_B[50][0] +
                mat_A[249][3] * mat_B[58][0] +
                mat_A[250][0] * mat_B[66][0] +
                mat_A[250][1] * mat_B[74][0] +
                mat_A[250][2] * mat_B[82][0] +
                mat_A[250][3] * mat_B[90][0] +
                mat_A[251][0] * mat_B[98][0] +
                mat_A[251][1] * mat_B[106][0] +
                mat_A[251][2] * mat_B[114][0] +
                mat_A[251][3] * mat_B[122][0] +
                mat_A[252][0] * mat_B[130][0] +
                mat_A[252][1] * mat_B[138][0] +
                mat_A[252][2] * mat_B[146][0] +
                mat_A[252][3] * mat_B[154][0] +
                mat_A[253][0] * mat_B[162][0] +
                mat_A[253][1] * mat_B[170][0] +
                mat_A[253][2] * mat_B[178][0] +
                mat_A[253][3] * mat_B[186][0] +
                mat_A[254][0] * mat_B[194][0] +
                mat_A[254][1] * mat_B[202][0] +
                mat_A[254][2] * mat_B[210][0] +
                mat_A[254][3] * mat_B[218][0] +
                mat_A[255][0] * mat_B[226][0] +
                mat_A[255][1] * mat_B[234][0] +
                mat_A[255][2] * mat_B[242][0] +
                mat_A[255][3] * mat_B[250][0];
    mat_C[250][1] <=
                mat_A[248][0] * mat_B[2][1] +
                mat_A[248][1] * mat_B[10][1] +
                mat_A[248][2] * mat_B[18][1] +
                mat_A[248][3] * mat_B[26][1] +
                mat_A[249][0] * mat_B[34][1] +
                mat_A[249][1] * mat_B[42][1] +
                mat_A[249][2] * mat_B[50][1] +
                mat_A[249][3] * mat_B[58][1] +
                mat_A[250][0] * mat_B[66][1] +
                mat_A[250][1] * mat_B[74][1] +
                mat_A[250][2] * mat_B[82][1] +
                mat_A[250][3] * mat_B[90][1] +
                mat_A[251][0] * mat_B[98][1] +
                mat_A[251][1] * mat_B[106][1] +
                mat_A[251][2] * mat_B[114][1] +
                mat_A[251][3] * mat_B[122][1] +
                mat_A[252][0] * mat_B[130][1] +
                mat_A[252][1] * mat_B[138][1] +
                mat_A[252][2] * mat_B[146][1] +
                mat_A[252][3] * mat_B[154][1] +
                mat_A[253][0] * mat_B[162][1] +
                mat_A[253][1] * mat_B[170][1] +
                mat_A[253][2] * mat_B[178][1] +
                mat_A[253][3] * mat_B[186][1] +
                mat_A[254][0] * mat_B[194][1] +
                mat_A[254][1] * mat_B[202][1] +
                mat_A[254][2] * mat_B[210][1] +
                mat_A[254][3] * mat_B[218][1] +
                mat_A[255][0] * mat_B[226][1] +
                mat_A[255][1] * mat_B[234][1] +
                mat_A[255][2] * mat_B[242][1] +
                mat_A[255][3] * mat_B[250][1];
    mat_C[250][2] <=
                mat_A[248][0] * mat_B[2][2] +
                mat_A[248][1] * mat_B[10][2] +
                mat_A[248][2] * mat_B[18][2] +
                mat_A[248][3] * mat_B[26][2] +
                mat_A[249][0] * mat_B[34][2] +
                mat_A[249][1] * mat_B[42][2] +
                mat_A[249][2] * mat_B[50][2] +
                mat_A[249][3] * mat_B[58][2] +
                mat_A[250][0] * mat_B[66][2] +
                mat_A[250][1] * mat_B[74][2] +
                mat_A[250][2] * mat_B[82][2] +
                mat_A[250][3] * mat_B[90][2] +
                mat_A[251][0] * mat_B[98][2] +
                mat_A[251][1] * mat_B[106][2] +
                mat_A[251][2] * mat_B[114][2] +
                mat_A[251][3] * mat_B[122][2] +
                mat_A[252][0] * mat_B[130][2] +
                mat_A[252][1] * mat_B[138][2] +
                mat_A[252][2] * mat_B[146][2] +
                mat_A[252][3] * mat_B[154][2] +
                mat_A[253][0] * mat_B[162][2] +
                mat_A[253][1] * mat_B[170][2] +
                mat_A[253][2] * mat_B[178][2] +
                mat_A[253][3] * mat_B[186][2] +
                mat_A[254][0] * mat_B[194][2] +
                mat_A[254][1] * mat_B[202][2] +
                mat_A[254][2] * mat_B[210][2] +
                mat_A[254][3] * mat_B[218][2] +
                mat_A[255][0] * mat_B[226][2] +
                mat_A[255][1] * mat_B[234][2] +
                mat_A[255][2] * mat_B[242][2] +
                mat_A[255][3] * mat_B[250][2];
    mat_C[250][3] <=
                mat_A[248][0] * mat_B[2][3] +
                mat_A[248][1] * mat_B[10][3] +
                mat_A[248][2] * mat_B[18][3] +
                mat_A[248][3] * mat_B[26][3] +
                mat_A[249][0] * mat_B[34][3] +
                mat_A[249][1] * mat_B[42][3] +
                mat_A[249][2] * mat_B[50][3] +
                mat_A[249][3] * mat_B[58][3] +
                mat_A[250][0] * mat_B[66][3] +
                mat_A[250][1] * mat_B[74][3] +
                mat_A[250][2] * mat_B[82][3] +
                mat_A[250][3] * mat_B[90][3] +
                mat_A[251][0] * mat_B[98][3] +
                mat_A[251][1] * mat_B[106][3] +
                mat_A[251][2] * mat_B[114][3] +
                mat_A[251][3] * mat_B[122][3] +
                mat_A[252][0] * mat_B[130][3] +
                mat_A[252][1] * mat_B[138][3] +
                mat_A[252][2] * mat_B[146][3] +
                mat_A[252][3] * mat_B[154][3] +
                mat_A[253][0] * mat_B[162][3] +
                mat_A[253][1] * mat_B[170][3] +
                mat_A[253][2] * mat_B[178][3] +
                mat_A[253][3] * mat_B[186][3] +
                mat_A[254][0] * mat_B[194][3] +
                mat_A[254][1] * mat_B[202][3] +
                mat_A[254][2] * mat_B[210][3] +
                mat_A[254][3] * mat_B[218][3] +
                mat_A[255][0] * mat_B[226][3] +
                mat_A[255][1] * mat_B[234][3] +
                mat_A[255][2] * mat_B[242][3] +
                mat_A[255][3] * mat_B[250][3];
    mat_C[251][0] <=
                mat_A[248][0] * mat_B[3][0] +
                mat_A[248][1] * mat_B[11][0] +
                mat_A[248][2] * mat_B[19][0] +
                mat_A[248][3] * mat_B[27][0] +
                mat_A[249][0] * mat_B[35][0] +
                mat_A[249][1] * mat_B[43][0] +
                mat_A[249][2] * mat_B[51][0] +
                mat_A[249][3] * mat_B[59][0] +
                mat_A[250][0] * mat_B[67][0] +
                mat_A[250][1] * mat_B[75][0] +
                mat_A[250][2] * mat_B[83][0] +
                mat_A[250][3] * mat_B[91][0] +
                mat_A[251][0] * mat_B[99][0] +
                mat_A[251][1] * mat_B[107][0] +
                mat_A[251][2] * mat_B[115][0] +
                mat_A[251][3] * mat_B[123][0] +
                mat_A[252][0] * mat_B[131][0] +
                mat_A[252][1] * mat_B[139][0] +
                mat_A[252][2] * mat_B[147][0] +
                mat_A[252][3] * mat_B[155][0] +
                mat_A[253][0] * mat_B[163][0] +
                mat_A[253][1] * mat_B[171][0] +
                mat_A[253][2] * mat_B[179][0] +
                mat_A[253][3] * mat_B[187][0] +
                mat_A[254][0] * mat_B[195][0] +
                mat_A[254][1] * mat_B[203][0] +
                mat_A[254][2] * mat_B[211][0] +
                mat_A[254][3] * mat_B[219][0] +
                mat_A[255][0] * mat_B[227][0] +
                mat_A[255][1] * mat_B[235][0] +
                mat_A[255][2] * mat_B[243][0] +
                mat_A[255][3] * mat_B[251][0];
    mat_C[251][1] <=
                mat_A[248][0] * mat_B[3][1] +
                mat_A[248][1] * mat_B[11][1] +
                mat_A[248][2] * mat_B[19][1] +
                mat_A[248][3] * mat_B[27][1] +
                mat_A[249][0] * mat_B[35][1] +
                mat_A[249][1] * mat_B[43][1] +
                mat_A[249][2] * mat_B[51][1] +
                mat_A[249][3] * mat_B[59][1] +
                mat_A[250][0] * mat_B[67][1] +
                mat_A[250][1] * mat_B[75][1] +
                mat_A[250][2] * mat_B[83][1] +
                mat_A[250][3] * mat_B[91][1] +
                mat_A[251][0] * mat_B[99][1] +
                mat_A[251][1] * mat_B[107][1] +
                mat_A[251][2] * mat_B[115][1] +
                mat_A[251][3] * mat_B[123][1] +
                mat_A[252][0] * mat_B[131][1] +
                mat_A[252][1] * mat_B[139][1] +
                mat_A[252][2] * mat_B[147][1] +
                mat_A[252][3] * mat_B[155][1] +
                mat_A[253][0] * mat_B[163][1] +
                mat_A[253][1] * mat_B[171][1] +
                mat_A[253][2] * mat_B[179][1] +
                mat_A[253][3] * mat_B[187][1] +
                mat_A[254][0] * mat_B[195][1] +
                mat_A[254][1] * mat_B[203][1] +
                mat_A[254][2] * mat_B[211][1] +
                mat_A[254][3] * mat_B[219][1] +
                mat_A[255][0] * mat_B[227][1] +
                mat_A[255][1] * mat_B[235][1] +
                mat_A[255][2] * mat_B[243][1] +
                mat_A[255][3] * mat_B[251][1];
    mat_C[251][2] <=
                mat_A[248][0] * mat_B[3][2] +
                mat_A[248][1] * mat_B[11][2] +
                mat_A[248][2] * mat_B[19][2] +
                mat_A[248][3] * mat_B[27][2] +
                mat_A[249][0] * mat_B[35][2] +
                mat_A[249][1] * mat_B[43][2] +
                mat_A[249][2] * mat_B[51][2] +
                mat_A[249][3] * mat_B[59][2] +
                mat_A[250][0] * mat_B[67][2] +
                mat_A[250][1] * mat_B[75][2] +
                mat_A[250][2] * mat_B[83][2] +
                mat_A[250][3] * mat_B[91][2] +
                mat_A[251][0] * mat_B[99][2] +
                mat_A[251][1] * mat_B[107][2] +
                mat_A[251][2] * mat_B[115][2] +
                mat_A[251][3] * mat_B[123][2] +
                mat_A[252][0] * mat_B[131][2] +
                mat_A[252][1] * mat_B[139][2] +
                mat_A[252][2] * mat_B[147][2] +
                mat_A[252][3] * mat_B[155][2] +
                mat_A[253][0] * mat_B[163][2] +
                mat_A[253][1] * mat_B[171][2] +
                mat_A[253][2] * mat_B[179][2] +
                mat_A[253][3] * mat_B[187][2] +
                mat_A[254][0] * mat_B[195][2] +
                mat_A[254][1] * mat_B[203][2] +
                mat_A[254][2] * mat_B[211][2] +
                mat_A[254][3] * mat_B[219][2] +
                mat_A[255][0] * mat_B[227][2] +
                mat_A[255][1] * mat_B[235][2] +
                mat_A[255][2] * mat_B[243][2] +
                mat_A[255][3] * mat_B[251][2];
    mat_C[251][3] <=
                mat_A[248][0] * mat_B[3][3] +
                mat_A[248][1] * mat_B[11][3] +
                mat_A[248][2] * mat_B[19][3] +
                mat_A[248][3] * mat_B[27][3] +
                mat_A[249][0] * mat_B[35][3] +
                mat_A[249][1] * mat_B[43][3] +
                mat_A[249][2] * mat_B[51][3] +
                mat_A[249][3] * mat_B[59][3] +
                mat_A[250][0] * mat_B[67][3] +
                mat_A[250][1] * mat_B[75][3] +
                mat_A[250][2] * mat_B[83][3] +
                mat_A[250][3] * mat_B[91][3] +
                mat_A[251][0] * mat_B[99][3] +
                mat_A[251][1] * mat_B[107][3] +
                mat_A[251][2] * mat_B[115][3] +
                mat_A[251][3] * mat_B[123][3] +
                mat_A[252][0] * mat_B[131][3] +
                mat_A[252][1] * mat_B[139][3] +
                mat_A[252][2] * mat_B[147][3] +
                mat_A[252][3] * mat_B[155][3] +
                mat_A[253][0] * mat_B[163][3] +
                mat_A[253][1] * mat_B[171][3] +
                mat_A[253][2] * mat_B[179][3] +
                mat_A[253][3] * mat_B[187][3] +
                mat_A[254][0] * mat_B[195][3] +
                mat_A[254][1] * mat_B[203][3] +
                mat_A[254][2] * mat_B[211][3] +
                mat_A[254][3] * mat_B[219][3] +
                mat_A[255][0] * mat_B[227][3] +
                mat_A[255][1] * mat_B[235][3] +
                mat_A[255][2] * mat_B[243][3] +
                mat_A[255][3] * mat_B[251][3];
    mat_C[252][0] <=
                mat_A[248][0] * mat_B[4][0] +
                mat_A[248][1] * mat_B[12][0] +
                mat_A[248][2] * mat_B[20][0] +
                mat_A[248][3] * mat_B[28][0] +
                mat_A[249][0] * mat_B[36][0] +
                mat_A[249][1] * mat_B[44][0] +
                mat_A[249][2] * mat_B[52][0] +
                mat_A[249][3] * mat_B[60][0] +
                mat_A[250][0] * mat_B[68][0] +
                mat_A[250][1] * mat_B[76][0] +
                mat_A[250][2] * mat_B[84][0] +
                mat_A[250][3] * mat_B[92][0] +
                mat_A[251][0] * mat_B[100][0] +
                mat_A[251][1] * mat_B[108][0] +
                mat_A[251][2] * mat_B[116][0] +
                mat_A[251][3] * mat_B[124][0] +
                mat_A[252][0] * mat_B[132][0] +
                mat_A[252][1] * mat_B[140][0] +
                mat_A[252][2] * mat_B[148][0] +
                mat_A[252][3] * mat_B[156][0] +
                mat_A[253][0] * mat_B[164][0] +
                mat_A[253][1] * mat_B[172][0] +
                mat_A[253][2] * mat_B[180][0] +
                mat_A[253][3] * mat_B[188][0] +
                mat_A[254][0] * mat_B[196][0] +
                mat_A[254][1] * mat_B[204][0] +
                mat_A[254][2] * mat_B[212][0] +
                mat_A[254][3] * mat_B[220][0] +
                mat_A[255][0] * mat_B[228][0] +
                mat_A[255][1] * mat_B[236][0] +
                mat_A[255][2] * mat_B[244][0] +
                mat_A[255][3] * mat_B[252][0];
    mat_C[252][1] <=
                mat_A[248][0] * mat_B[4][1] +
                mat_A[248][1] * mat_B[12][1] +
                mat_A[248][2] * mat_B[20][1] +
                mat_A[248][3] * mat_B[28][1] +
                mat_A[249][0] * mat_B[36][1] +
                mat_A[249][1] * mat_B[44][1] +
                mat_A[249][2] * mat_B[52][1] +
                mat_A[249][3] * mat_B[60][1] +
                mat_A[250][0] * mat_B[68][1] +
                mat_A[250][1] * mat_B[76][1] +
                mat_A[250][2] * mat_B[84][1] +
                mat_A[250][3] * mat_B[92][1] +
                mat_A[251][0] * mat_B[100][1] +
                mat_A[251][1] * mat_B[108][1] +
                mat_A[251][2] * mat_B[116][1] +
                mat_A[251][3] * mat_B[124][1] +
                mat_A[252][0] * mat_B[132][1] +
                mat_A[252][1] * mat_B[140][1] +
                mat_A[252][2] * mat_B[148][1] +
                mat_A[252][3] * mat_B[156][1] +
                mat_A[253][0] * mat_B[164][1] +
                mat_A[253][1] * mat_B[172][1] +
                mat_A[253][2] * mat_B[180][1] +
                mat_A[253][3] * mat_B[188][1] +
                mat_A[254][0] * mat_B[196][1] +
                mat_A[254][1] * mat_B[204][1] +
                mat_A[254][2] * mat_B[212][1] +
                mat_A[254][3] * mat_B[220][1] +
                mat_A[255][0] * mat_B[228][1] +
                mat_A[255][1] * mat_B[236][1] +
                mat_A[255][2] * mat_B[244][1] +
                mat_A[255][3] * mat_B[252][1];
    mat_C[252][2] <=
                mat_A[248][0] * mat_B[4][2] +
                mat_A[248][1] * mat_B[12][2] +
                mat_A[248][2] * mat_B[20][2] +
                mat_A[248][3] * mat_B[28][2] +
                mat_A[249][0] * mat_B[36][2] +
                mat_A[249][1] * mat_B[44][2] +
                mat_A[249][2] * mat_B[52][2] +
                mat_A[249][3] * mat_B[60][2] +
                mat_A[250][0] * mat_B[68][2] +
                mat_A[250][1] * mat_B[76][2] +
                mat_A[250][2] * mat_B[84][2] +
                mat_A[250][3] * mat_B[92][2] +
                mat_A[251][0] * mat_B[100][2] +
                mat_A[251][1] * mat_B[108][2] +
                mat_A[251][2] * mat_B[116][2] +
                mat_A[251][3] * mat_B[124][2] +
                mat_A[252][0] * mat_B[132][2] +
                mat_A[252][1] * mat_B[140][2] +
                mat_A[252][2] * mat_B[148][2] +
                mat_A[252][3] * mat_B[156][2] +
                mat_A[253][0] * mat_B[164][2] +
                mat_A[253][1] * mat_B[172][2] +
                mat_A[253][2] * mat_B[180][2] +
                mat_A[253][3] * mat_B[188][2] +
                mat_A[254][0] * mat_B[196][2] +
                mat_A[254][1] * mat_B[204][2] +
                mat_A[254][2] * mat_B[212][2] +
                mat_A[254][3] * mat_B[220][2] +
                mat_A[255][0] * mat_B[228][2] +
                mat_A[255][1] * mat_B[236][2] +
                mat_A[255][2] * mat_B[244][2] +
                mat_A[255][3] * mat_B[252][2];
    mat_C[252][3] <=
                mat_A[248][0] * mat_B[4][3] +
                mat_A[248][1] * mat_B[12][3] +
                mat_A[248][2] * mat_B[20][3] +
                mat_A[248][3] * mat_B[28][3] +
                mat_A[249][0] * mat_B[36][3] +
                mat_A[249][1] * mat_B[44][3] +
                mat_A[249][2] * mat_B[52][3] +
                mat_A[249][3] * mat_B[60][3] +
                mat_A[250][0] * mat_B[68][3] +
                mat_A[250][1] * mat_B[76][3] +
                mat_A[250][2] * mat_B[84][3] +
                mat_A[250][3] * mat_B[92][3] +
                mat_A[251][0] * mat_B[100][3] +
                mat_A[251][1] * mat_B[108][3] +
                mat_A[251][2] * mat_B[116][3] +
                mat_A[251][3] * mat_B[124][3] +
                mat_A[252][0] * mat_B[132][3] +
                mat_A[252][1] * mat_B[140][3] +
                mat_A[252][2] * mat_B[148][3] +
                mat_A[252][3] * mat_B[156][3] +
                mat_A[253][0] * mat_B[164][3] +
                mat_A[253][1] * mat_B[172][3] +
                mat_A[253][2] * mat_B[180][3] +
                mat_A[253][3] * mat_B[188][3] +
                mat_A[254][0] * mat_B[196][3] +
                mat_A[254][1] * mat_B[204][3] +
                mat_A[254][2] * mat_B[212][3] +
                mat_A[254][3] * mat_B[220][3] +
                mat_A[255][0] * mat_B[228][3] +
                mat_A[255][1] * mat_B[236][3] +
                mat_A[255][2] * mat_B[244][3] +
                mat_A[255][3] * mat_B[252][3];
    mat_C[253][0] <=
                mat_A[248][0] * mat_B[5][0] +
                mat_A[248][1] * mat_B[13][0] +
                mat_A[248][2] * mat_B[21][0] +
                mat_A[248][3] * mat_B[29][0] +
                mat_A[249][0] * mat_B[37][0] +
                mat_A[249][1] * mat_B[45][0] +
                mat_A[249][2] * mat_B[53][0] +
                mat_A[249][3] * mat_B[61][0] +
                mat_A[250][0] * mat_B[69][0] +
                mat_A[250][1] * mat_B[77][0] +
                mat_A[250][2] * mat_B[85][0] +
                mat_A[250][3] * mat_B[93][0] +
                mat_A[251][0] * mat_B[101][0] +
                mat_A[251][1] * mat_B[109][0] +
                mat_A[251][2] * mat_B[117][0] +
                mat_A[251][3] * mat_B[125][0] +
                mat_A[252][0] * mat_B[133][0] +
                mat_A[252][1] * mat_B[141][0] +
                mat_A[252][2] * mat_B[149][0] +
                mat_A[252][3] * mat_B[157][0] +
                mat_A[253][0] * mat_B[165][0] +
                mat_A[253][1] * mat_B[173][0] +
                mat_A[253][2] * mat_B[181][0] +
                mat_A[253][3] * mat_B[189][0] +
                mat_A[254][0] * mat_B[197][0] +
                mat_A[254][1] * mat_B[205][0] +
                mat_A[254][2] * mat_B[213][0] +
                mat_A[254][3] * mat_B[221][0] +
                mat_A[255][0] * mat_B[229][0] +
                mat_A[255][1] * mat_B[237][0] +
                mat_A[255][2] * mat_B[245][0] +
                mat_A[255][3] * mat_B[253][0];
    mat_C[253][1] <=
                mat_A[248][0] * mat_B[5][1] +
                mat_A[248][1] * mat_B[13][1] +
                mat_A[248][2] * mat_B[21][1] +
                mat_A[248][3] * mat_B[29][1] +
                mat_A[249][0] * mat_B[37][1] +
                mat_A[249][1] * mat_B[45][1] +
                mat_A[249][2] * mat_B[53][1] +
                mat_A[249][3] * mat_B[61][1] +
                mat_A[250][0] * mat_B[69][1] +
                mat_A[250][1] * mat_B[77][1] +
                mat_A[250][2] * mat_B[85][1] +
                mat_A[250][3] * mat_B[93][1] +
                mat_A[251][0] * mat_B[101][1] +
                mat_A[251][1] * mat_B[109][1] +
                mat_A[251][2] * mat_B[117][1] +
                mat_A[251][3] * mat_B[125][1] +
                mat_A[252][0] * mat_B[133][1] +
                mat_A[252][1] * mat_B[141][1] +
                mat_A[252][2] * mat_B[149][1] +
                mat_A[252][3] * mat_B[157][1] +
                mat_A[253][0] * mat_B[165][1] +
                mat_A[253][1] * mat_B[173][1] +
                mat_A[253][2] * mat_B[181][1] +
                mat_A[253][3] * mat_B[189][1] +
                mat_A[254][0] * mat_B[197][1] +
                mat_A[254][1] * mat_B[205][1] +
                mat_A[254][2] * mat_B[213][1] +
                mat_A[254][3] * mat_B[221][1] +
                mat_A[255][0] * mat_B[229][1] +
                mat_A[255][1] * mat_B[237][1] +
                mat_A[255][2] * mat_B[245][1] +
                mat_A[255][3] * mat_B[253][1];
    mat_C[253][2] <=
                mat_A[248][0] * mat_B[5][2] +
                mat_A[248][1] * mat_B[13][2] +
                mat_A[248][2] * mat_B[21][2] +
                mat_A[248][3] * mat_B[29][2] +
                mat_A[249][0] * mat_B[37][2] +
                mat_A[249][1] * mat_B[45][2] +
                mat_A[249][2] * mat_B[53][2] +
                mat_A[249][3] * mat_B[61][2] +
                mat_A[250][0] * mat_B[69][2] +
                mat_A[250][1] * mat_B[77][2] +
                mat_A[250][2] * mat_B[85][2] +
                mat_A[250][3] * mat_B[93][2] +
                mat_A[251][0] * mat_B[101][2] +
                mat_A[251][1] * mat_B[109][2] +
                mat_A[251][2] * mat_B[117][2] +
                mat_A[251][3] * mat_B[125][2] +
                mat_A[252][0] * mat_B[133][2] +
                mat_A[252][1] * mat_B[141][2] +
                mat_A[252][2] * mat_B[149][2] +
                mat_A[252][3] * mat_B[157][2] +
                mat_A[253][0] * mat_B[165][2] +
                mat_A[253][1] * mat_B[173][2] +
                mat_A[253][2] * mat_B[181][2] +
                mat_A[253][3] * mat_B[189][2] +
                mat_A[254][0] * mat_B[197][2] +
                mat_A[254][1] * mat_B[205][2] +
                mat_A[254][2] * mat_B[213][2] +
                mat_A[254][3] * mat_B[221][2] +
                mat_A[255][0] * mat_B[229][2] +
                mat_A[255][1] * mat_B[237][2] +
                mat_A[255][2] * mat_B[245][2] +
                mat_A[255][3] * mat_B[253][2];
    mat_C[253][3] <=
                mat_A[248][0] * mat_B[5][3] +
                mat_A[248][1] * mat_B[13][3] +
                mat_A[248][2] * mat_B[21][3] +
                mat_A[248][3] * mat_B[29][3] +
                mat_A[249][0] * mat_B[37][3] +
                mat_A[249][1] * mat_B[45][3] +
                mat_A[249][2] * mat_B[53][3] +
                mat_A[249][3] * mat_B[61][3] +
                mat_A[250][0] * mat_B[69][3] +
                mat_A[250][1] * mat_B[77][3] +
                mat_A[250][2] * mat_B[85][3] +
                mat_A[250][3] * mat_B[93][3] +
                mat_A[251][0] * mat_B[101][3] +
                mat_A[251][1] * mat_B[109][3] +
                mat_A[251][2] * mat_B[117][3] +
                mat_A[251][3] * mat_B[125][3] +
                mat_A[252][0] * mat_B[133][3] +
                mat_A[252][1] * mat_B[141][3] +
                mat_A[252][2] * mat_B[149][3] +
                mat_A[252][3] * mat_B[157][3] +
                mat_A[253][0] * mat_B[165][3] +
                mat_A[253][1] * mat_B[173][3] +
                mat_A[253][2] * mat_B[181][3] +
                mat_A[253][3] * mat_B[189][3] +
                mat_A[254][0] * mat_B[197][3] +
                mat_A[254][1] * mat_B[205][3] +
                mat_A[254][2] * mat_B[213][3] +
                mat_A[254][3] * mat_B[221][3] +
                mat_A[255][0] * mat_B[229][3] +
                mat_A[255][1] * mat_B[237][3] +
                mat_A[255][2] * mat_B[245][3] +
                mat_A[255][3] * mat_B[253][3];
    mat_C[254][0] <=
                mat_A[248][0] * mat_B[6][0] +
                mat_A[248][1] * mat_B[14][0] +
                mat_A[248][2] * mat_B[22][0] +
                mat_A[248][3] * mat_B[30][0] +
                mat_A[249][0] * mat_B[38][0] +
                mat_A[249][1] * mat_B[46][0] +
                mat_A[249][2] * mat_B[54][0] +
                mat_A[249][3] * mat_B[62][0] +
                mat_A[250][0] * mat_B[70][0] +
                mat_A[250][1] * mat_B[78][0] +
                mat_A[250][2] * mat_B[86][0] +
                mat_A[250][3] * mat_B[94][0] +
                mat_A[251][0] * mat_B[102][0] +
                mat_A[251][1] * mat_B[110][0] +
                mat_A[251][2] * mat_B[118][0] +
                mat_A[251][3] * mat_B[126][0] +
                mat_A[252][0] * mat_B[134][0] +
                mat_A[252][1] * mat_B[142][0] +
                mat_A[252][2] * mat_B[150][0] +
                mat_A[252][3] * mat_B[158][0] +
                mat_A[253][0] * mat_B[166][0] +
                mat_A[253][1] * mat_B[174][0] +
                mat_A[253][2] * mat_B[182][0] +
                mat_A[253][3] * mat_B[190][0] +
                mat_A[254][0] * mat_B[198][0] +
                mat_A[254][1] * mat_B[206][0] +
                mat_A[254][2] * mat_B[214][0] +
                mat_A[254][3] * mat_B[222][0] +
                mat_A[255][0] * mat_B[230][0] +
                mat_A[255][1] * mat_B[238][0] +
                mat_A[255][2] * mat_B[246][0] +
                mat_A[255][3] * mat_B[254][0];
    mat_C[254][1] <=
                mat_A[248][0] * mat_B[6][1] +
                mat_A[248][1] * mat_B[14][1] +
                mat_A[248][2] * mat_B[22][1] +
                mat_A[248][3] * mat_B[30][1] +
                mat_A[249][0] * mat_B[38][1] +
                mat_A[249][1] * mat_B[46][1] +
                mat_A[249][2] * mat_B[54][1] +
                mat_A[249][3] * mat_B[62][1] +
                mat_A[250][0] * mat_B[70][1] +
                mat_A[250][1] * mat_B[78][1] +
                mat_A[250][2] * mat_B[86][1] +
                mat_A[250][3] * mat_B[94][1] +
                mat_A[251][0] * mat_B[102][1] +
                mat_A[251][1] * mat_B[110][1] +
                mat_A[251][2] * mat_B[118][1] +
                mat_A[251][3] * mat_B[126][1] +
                mat_A[252][0] * mat_B[134][1] +
                mat_A[252][1] * mat_B[142][1] +
                mat_A[252][2] * mat_B[150][1] +
                mat_A[252][3] * mat_B[158][1] +
                mat_A[253][0] * mat_B[166][1] +
                mat_A[253][1] * mat_B[174][1] +
                mat_A[253][2] * mat_B[182][1] +
                mat_A[253][3] * mat_B[190][1] +
                mat_A[254][0] * mat_B[198][1] +
                mat_A[254][1] * mat_B[206][1] +
                mat_A[254][2] * mat_B[214][1] +
                mat_A[254][3] * mat_B[222][1] +
                mat_A[255][0] * mat_B[230][1] +
                mat_A[255][1] * mat_B[238][1] +
                mat_A[255][2] * mat_B[246][1] +
                mat_A[255][3] * mat_B[254][1];
    mat_C[254][2] <=
                mat_A[248][0] * mat_B[6][2] +
                mat_A[248][1] * mat_B[14][2] +
                mat_A[248][2] * mat_B[22][2] +
                mat_A[248][3] * mat_B[30][2] +
                mat_A[249][0] * mat_B[38][2] +
                mat_A[249][1] * mat_B[46][2] +
                mat_A[249][2] * mat_B[54][2] +
                mat_A[249][3] * mat_B[62][2] +
                mat_A[250][0] * mat_B[70][2] +
                mat_A[250][1] * mat_B[78][2] +
                mat_A[250][2] * mat_B[86][2] +
                mat_A[250][3] * mat_B[94][2] +
                mat_A[251][0] * mat_B[102][2] +
                mat_A[251][1] * mat_B[110][2] +
                mat_A[251][2] * mat_B[118][2] +
                mat_A[251][3] * mat_B[126][2] +
                mat_A[252][0] * mat_B[134][2] +
                mat_A[252][1] * mat_B[142][2] +
                mat_A[252][2] * mat_B[150][2] +
                mat_A[252][3] * mat_B[158][2] +
                mat_A[253][0] * mat_B[166][2] +
                mat_A[253][1] * mat_B[174][2] +
                mat_A[253][2] * mat_B[182][2] +
                mat_A[253][3] * mat_B[190][2] +
                mat_A[254][0] * mat_B[198][2] +
                mat_A[254][1] * mat_B[206][2] +
                mat_A[254][2] * mat_B[214][2] +
                mat_A[254][3] * mat_B[222][2] +
                mat_A[255][0] * mat_B[230][2] +
                mat_A[255][1] * mat_B[238][2] +
                mat_A[255][2] * mat_B[246][2] +
                mat_A[255][3] * mat_B[254][2];
    mat_C[254][3] <=
                mat_A[248][0] * mat_B[6][3] +
                mat_A[248][1] * mat_B[14][3] +
                mat_A[248][2] * mat_B[22][3] +
                mat_A[248][3] * mat_B[30][3] +
                mat_A[249][0] * mat_B[38][3] +
                mat_A[249][1] * mat_B[46][3] +
                mat_A[249][2] * mat_B[54][3] +
                mat_A[249][3] * mat_B[62][3] +
                mat_A[250][0] * mat_B[70][3] +
                mat_A[250][1] * mat_B[78][3] +
                mat_A[250][2] * mat_B[86][3] +
                mat_A[250][3] * mat_B[94][3] +
                mat_A[251][0] * mat_B[102][3] +
                mat_A[251][1] * mat_B[110][3] +
                mat_A[251][2] * mat_B[118][3] +
                mat_A[251][3] * mat_B[126][3] +
                mat_A[252][0] * mat_B[134][3] +
                mat_A[252][1] * mat_B[142][3] +
                mat_A[252][2] * mat_B[150][3] +
                mat_A[252][3] * mat_B[158][3] +
                mat_A[253][0] * mat_B[166][3] +
                mat_A[253][1] * mat_B[174][3] +
                mat_A[253][2] * mat_B[182][3] +
                mat_A[253][3] * mat_B[190][3] +
                mat_A[254][0] * mat_B[198][3] +
                mat_A[254][1] * mat_B[206][3] +
                mat_A[254][2] * mat_B[214][3] +
                mat_A[254][3] * mat_B[222][3] +
                mat_A[255][0] * mat_B[230][3] +
                mat_A[255][1] * mat_B[238][3] +
                mat_A[255][2] * mat_B[246][3] +
                mat_A[255][3] * mat_B[254][3];
    mat_C[255][0] <=
                mat_A[248][0] * mat_B[7][0] +
                mat_A[248][1] * mat_B[15][0] +
                mat_A[248][2] * mat_B[23][0] +
                mat_A[248][3] * mat_B[31][0] +
                mat_A[249][0] * mat_B[39][0] +
                mat_A[249][1] * mat_B[47][0] +
                mat_A[249][2] * mat_B[55][0] +
                mat_A[249][3] * mat_B[63][0] +
                mat_A[250][0] * mat_B[71][0] +
                mat_A[250][1] * mat_B[79][0] +
                mat_A[250][2] * mat_B[87][0] +
                mat_A[250][3] * mat_B[95][0] +
                mat_A[251][0] * mat_B[103][0] +
                mat_A[251][1] * mat_B[111][0] +
                mat_A[251][2] * mat_B[119][0] +
                mat_A[251][3] * mat_B[127][0] +
                mat_A[252][0] * mat_B[135][0] +
                mat_A[252][1] * mat_B[143][0] +
                mat_A[252][2] * mat_B[151][0] +
                mat_A[252][3] * mat_B[159][0] +
                mat_A[253][0] * mat_B[167][0] +
                mat_A[253][1] * mat_B[175][0] +
                mat_A[253][2] * mat_B[183][0] +
                mat_A[253][3] * mat_B[191][0] +
                mat_A[254][0] * mat_B[199][0] +
                mat_A[254][1] * mat_B[207][0] +
                mat_A[254][2] * mat_B[215][0] +
                mat_A[254][3] * mat_B[223][0] +
                mat_A[255][0] * mat_B[231][0] +
                mat_A[255][1] * mat_B[239][0] +
                mat_A[255][2] * mat_B[247][0] +
                mat_A[255][3] * mat_B[255][0];
    mat_C[255][1] <=
                mat_A[248][0] * mat_B[7][1] +
                mat_A[248][1] * mat_B[15][1] +
                mat_A[248][2] * mat_B[23][1] +
                mat_A[248][3] * mat_B[31][1] +
                mat_A[249][0] * mat_B[39][1] +
                mat_A[249][1] * mat_B[47][1] +
                mat_A[249][2] * mat_B[55][1] +
                mat_A[249][3] * mat_B[63][1] +
                mat_A[250][0] * mat_B[71][1] +
                mat_A[250][1] * mat_B[79][1] +
                mat_A[250][2] * mat_B[87][1] +
                mat_A[250][3] * mat_B[95][1] +
                mat_A[251][0] * mat_B[103][1] +
                mat_A[251][1] * mat_B[111][1] +
                mat_A[251][2] * mat_B[119][1] +
                mat_A[251][3] * mat_B[127][1] +
                mat_A[252][0] * mat_B[135][1] +
                mat_A[252][1] * mat_B[143][1] +
                mat_A[252][2] * mat_B[151][1] +
                mat_A[252][3] * mat_B[159][1] +
                mat_A[253][0] * mat_B[167][1] +
                mat_A[253][1] * mat_B[175][1] +
                mat_A[253][2] * mat_B[183][1] +
                mat_A[253][3] * mat_B[191][1] +
                mat_A[254][0] * mat_B[199][1] +
                mat_A[254][1] * mat_B[207][1] +
                mat_A[254][2] * mat_B[215][1] +
                mat_A[254][3] * mat_B[223][1] +
                mat_A[255][0] * mat_B[231][1] +
                mat_A[255][1] * mat_B[239][1] +
                mat_A[255][2] * mat_B[247][1] +
                mat_A[255][3] * mat_B[255][1];
    mat_C[255][2] <=
                mat_A[248][0] * mat_B[7][2] +
                mat_A[248][1] * mat_B[15][2] +
                mat_A[248][2] * mat_B[23][2] +
                mat_A[248][3] * mat_B[31][2] +
                mat_A[249][0] * mat_B[39][2] +
                mat_A[249][1] * mat_B[47][2] +
                mat_A[249][2] * mat_B[55][2] +
                mat_A[249][3] * mat_B[63][2] +
                mat_A[250][0] * mat_B[71][2] +
                mat_A[250][1] * mat_B[79][2] +
                mat_A[250][2] * mat_B[87][2] +
                mat_A[250][3] * mat_B[95][2] +
                mat_A[251][0] * mat_B[103][2] +
                mat_A[251][1] * mat_B[111][2] +
                mat_A[251][2] * mat_B[119][2] +
                mat_A[251][3] * mat_B[127][2] +
                mat_A[252][0] * mat_B[135][2] +
                mat_A[252][1] * mat_B[143][2] +
                mat_A[252][2] * mat_B[151][2] +
                mat_A[252][3] * mat_B[159][2] +
                mat_A[253][0] * mat_B[167][2] +
                mat_A[253][1] * mat_B[175][2] +
                mat_A[253][2] * mat_B[183][2] +
                mat_A[253][3] * mat_B[191][2] +
                mat_A[254][0] * mat_B[199][2] +
                mat_A[254][1] * mat_B[207][2] +
                mat_A[254][2] * mat_B[215][2] +
                mat_A[254][3] * mat_B[223][2] +
                mat_A[255][0] * mat_B[231][2] +
                mat_A[255][1] * mat_B[239][2] +
                mat_A[255][2] * mat_B[247][2] +
                mat_A[255][3] * mat_B[255][2];
    mat_C[255][3] <=
                mat_A[248][0] * mat_B[7][3] +
                mat_A[248][1] * mat_B[15][3] +
                mat_A[248][2] * mat_B[23][3] +
                mat_A[248][3] * mat_B[31][3] +
                mat_A[249][0] * mat_B[39][3] +
                mat_A[249][1] * mat_B[47][3] +
                mat_A[249][2] * mat_B[55][3] +
                mat_A[249][3] * mat_B[63][3] +
                mat_A[250][0] * mat_B[71][3] +
                mat_A[250][1] * mat_B[79][3] +
                mat_A[250][2] * mat_B[87][3] +
                mat_A[250][3] * mat_B[95][3] +
                mat_A[251][0] * mat_B[103][3] +
                mat_A[251][1] * mat_B[111][3] +
                mat_A[251][2] * mat_B[119][3] +
                mat_A[251][3] * mat_B[127][3] +
                mat_A[252][0] * mat_B[135][3] +
                mat_A[252][1] * mat_B[143][3] +
                mat_A[252][2] * mat_B[151][3] +
                mat_A[252][3] * mat_B[159][3] +
                mat_A[253][0] * mat_B[167][3] +
                mat_A[253][1] * mat_B[175][3] +
                mat_A[253][2] * mat_B[183][3] +
                mat_A[253][3] * mat_B[191][3] +
                mat_A[254][0] * mat_B[199][3] +
                mat_A[254][1] * mat_B[207][3] +
                mat_A[254][2] * mat_B[215][3] +
                mat_A[254][3] * mat_B[223][3] +
                mat_A[255][0] * mat_B[231][3] +
                mat_A[255][1] * mat_B[239][3] +
                mat_A[255][2] * mat_B[247][3] +
                mat_A[255][3] * mat_B[255][3];
                  end
endmodule
